module configurable_param_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_addr[0] ;
 wire \rd_addr[1] ;
 wire \rd_addr[2] ;
 wire \rd_addr[3] ;
 wire \rd_data_reg[0] ;
 wire \rd_data_reg[1] ;
 wire \rd_data_reg[2] ;
 wire \rd_data_reg[3] ;
 wire \rd_data_reg[4] ;
 wire \rd_data_reg[5] ;
 wire \rd_data_reg[6] ;
 wire \rd_data_reg[7] ;
 wire \rd_ptr[4] ;
 wire rd_valid;
 wire \wr_addr[0] ;
 wire \wr_addr[1] ;
 wire \wr_addr[2] ;
 wire \wr_addr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net25;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _340_ (.A1(\wr_ptr[4] ),
    .A2(\rd_ptr[4] ),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _341_ (.A1(_330_),
    .A2(_325_),
    .A3(_328_),
    .A4(_322_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _342_ (.A1(_152_),
    .A2(_153_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _343_ (.I(_154_),
    .ZN(net15));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _344_ (.A1(\wr_ptr[4] ),
    .A2(\rd_ptr[4] ),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _345_ (.A1(_155_),
    .A2(_153_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _346_ (.I(_156_),
    .ZN(net16));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _347_ (.A1(net2),
    .A2(_154_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _348_ (.I(_157_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _349_ (.I(\rd_addr[1] ),
    .Z(_158_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _350_ (.I(_158_),
    .Z(_159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _351_ (.I(_159_),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _352_ (.I(\rd_addr[3] ),
    .Z(_160_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _353_ (.I(_160_),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _354_ (.I(\rd_addr[2] ),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _355_ (.I(_161_),
    .Z(_326_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _356_ (.I(_329_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _357_ (.I(\wr_addr[0] ),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _358_ (.I(\wr_addr[1] ),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _359_ (.I(_322_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _360_ (.I(_321_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _361_ (.A1(_329_),
    .A2(_162_),
    .B(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _362_ (.A1(_328_),
    .A2(_164_),
    .B(_327_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _363_ (.A1(_325_),
    .A2(_165_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _364_ (.I(_330_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _365_ (.A1(_167_),
    .A2(_320_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _366_ (.A1(_325_),
    .A2(_328_),
    .A3(_319_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _367_ (.A1(_325_),
    .A2(_327_),
    .B(_169_),
    .C(_324_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _368_ (.A1(_155_),
    .A2(_170_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _369_ (.A1(_328_),
    .A2(_319_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _370_ (.A1(net13),
    .A2(_168_),
    .B(_171_),
    .C(_172_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _371_ (.A1(_166_),
    .A2(_173_),
    .B(_154_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _372_ (.A1(_325_),
    .A2(_165_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _373_ (.A1(_167_),
    .A2(net14),
    .B(_320_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _374_ (.A1(_172_),
    .A2(_175_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _375_ (.A1(_174_),
    .A2(_176_),
    .B(_171_),
    .C(_156_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _376_ (.I(net4),
    .Z(_177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _377_ (.I(\wr_addr[3] ),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _378_ (.I(\wr_addr[2] ),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _379_ (.A1(net12),
    .A2(_178_),
    .A3(_179_),
    .A4(_156_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _380_ (.A1(_333_),
    .A2(_180_),
    .Z(_181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _381_ (.I0(\mem[0][0] ),
    .I1(_177_),
    .S(_181_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _382_ (.I(net5),
    .Z(_182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _383_ (.I0(\mem[0][1] ),
    .I1(_182_),
    .S(_181_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _384_ (.I(net6),
    .Z(_183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _385_ (.I0(\mem[0][2] ),
    .I1(_183_),
    .S(_181_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _386_ (.I(net7),
    .Z(_184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _387_ (.I0(\mem[0][3] ),
    .I1(_184_),
    .S(_181_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _388_ (.I(net8),
    .Z(_185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _389_ (.I0(\mem[0][4] ),
    .I1(_185_),
    .S(_181_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _390_ (.I(net9),
    .Z(_186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _391_ (.I0(\mem[0][5] ),
    .I1(_186_),
    .S(_181_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _392_ (.I(net10),
    .Z(_187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _393_ (.I0(\mem[0][6] ),
    .I1(_187_),
    .S(_181_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _394_ (.I(net11),
    .Z(_188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _395_ (.I0(\mem[0][7] ),
    .I1(_188_),
    .S(_181_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _396_ (.A1(net12),
    .A2(\wr_addr[3] ),
    .A3(_179_),
    .A4(_156_),
    .Z(_189_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _397_ (.A1(_334_),
    .A2(_189_),
    .Z(_190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _398_ (.I0(\mem[10][0] ),
    .I1(_177_),
    .S(_190_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _399_ (.I0(\mem[10][1] ),
    .I1(_182_),
    .S(_190_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _400_ (.I0(\mem[10][2] ),
    .I1(_183_),
    .S(_190_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _401_ (.I0(\mem[10][3] ),
    .I1(_184_),
    .S(_190_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _402_ (.I0(\mem[10][4] ),
    .I1(_185_),
    .S(_190_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _403_ (.I0(\mem[10][5] ),
    .I1(_186_),
    .S(_190_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _404_ (.I0(\mem[10][6] ),
    .I1(_187_),
    .S(_190_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _405_ (.I0(\mem[10][7] ),
    .I1(_188_),
    .S(_190_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _406_ (.A1(_338_),
    .A2(_189_),
    .Z(_191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _407_ (.I0(\mem[11][0] ),
    .I1(_177_),
    .S(_191_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _408_ (.I0(\mem[11][1] ),
    .I1(_182_),
    .S(_191_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _409_ (.I0(\mem[11][2] ),
    .I1(_183_),
    .S(_191_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _410_ (.I0(\mem[11][3] ),
    .I1(_184_),
    .S(_191_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _411_ (.I0(\mem[11][4] ),
    .I1(_185_),
    .S(_191_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _412_ (.I0(\mem[11][5] ),
    .I1(_186_),
    .S(_191_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _413_ (.I0(\mem[11][6] ),
    .I1(_187_),
    .S(_191_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _414_ (.I0(\mem[11][7] ),
    .I1(_188_),
    .S(_191_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _415_ (.A1(net12),
    .A2(\wr_addr[3] ),
    .A3(\wr_addr[2] ),
    .A4(_156_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _416_ (.A1(_333_),
    .A2(_192_),
    .Z(_193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _417_ (.I0(\mem[12][0] ),
    .I1(_177_),
    .S(_193_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _418_ (.I0(\mem[12][1] ),
    .I1(_182_),
    .S(_193_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _419_ (.I0(\mem[12][2] ),
    .I1(_183_),
    .S(_193_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _420_ (.I0(\mem[12][3] ),
    .I1(_184_),
    .S(_193_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _421_ (.I0(\mem[12][4] ),
    .I1(_185_),
    .S(_193_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _422_ (.I0(\mem[12][5] ),
    .I1(_186_),
    .S(_193_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _423_ (.I0(\mem[12][6] ),
    .I1(_187_),
    .S(_193_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _424_ (.I0(\mem[12][7] ),
    .I1(_188_),
    .S(_193_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _425_ (.A1(_336_),
    .A2(_192_),
    .Z(_194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _426_ (.I0(\mem[13][0] ),
    .I1(_177_),
    .S(_194_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _427_ (.I0(\mem[13][1] ),
    .I1(_182_),
    .S(_194_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _428_ (.I0(\mem[13][2] ),
    .I1(_183_),
    .S(_194_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _429_ (.I0(\mem[13][3] ),
    .I1(_184_),
    .S(_194_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _430_ (.I0(\mem[13][4] ),
    .I1(_185_),
    .S(_194_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _431_ (.I0(\mem[13][5] ),
    .I1(_186_),
    .S(_194_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _432_ (.I0(\mem[13][6] ),
    .I1(_187_),
    .S(_194_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _433_ (.I0(\mem[13][7] ),
    .I1(_188_),
    .S(_194_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _434_ (.A1(_334_),
    .A2(_192_),
    .Z(_195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _435_ (.I0(\mem[14][0] ),
    .I1(_177_),
    .S(_195_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _436_ (.I0(\mem[14][1] ),
    .I1(_182_),
    .S(_195_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _437_ (.I0(\mem[14][2] ),
    .I1(_183_),
    .S(_195_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _438_ (.I0(\mem[14][3] ),
    .I1(_184_),
    .S(_195_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _439_ (.I0(\mem[14][4] ),
    .I1(_185_),
    .S(_195_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _440_ (.I0(\mem[14][5] ),
    .I1(_186_),
    .S(_195_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _441_ (.I0(\mem[14][6] ),
    .I1(_187_),
    .S(_195_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _442_ (.I0(\mem[14][7] ),
    .I1(_188_),
    .S(_195_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _443_ (.A1(_338_),
    .A2(_192_),
    .Z(_196_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _444_ (.I(_196_),
    .Z(_197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _445_ (.I0(\mem[15][0] ),
    .I1(_177_),
    .S(_197_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _446_ (.I0(\mem[15][1] ),
    .I1(_182_),
    .S(_197_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _447_ (.I0(\mem[15][2] ),
    .I1(_183_),
    .S(_197_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _448_ (.I0(\mem[15][3] ),
    .I1(_184_),
    .S(_197_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _449_ (.I0(\mem[15][4] ),
    .I1(_185_),
    .S(_197_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _450_ (.I0(\mem[15][5] ),
    .I1(_186_),
    .S(_197_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _451_ (.I0(\mem[15][6] ),
    .I1(_187_),
    .S(_197_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _452_ (.I0(\mem[15][7] ),
    .I1(_188_),
    .S(_197_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _453_ (.A1(_336_),
    .A2(_180_),
    .Z(_198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _454_ (.I0(\mem[1][0] ),
    .I1(_177_),
    .S(_198_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _455_ (.I0(\mem[1][1] ),
    .I1(_182_),
    .S(_198_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _456_ (.I0(\mem[1][2] ),
    .I1(_183_),
    .S(_198_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _457_ (.I0(\mem[1][3] ),
    .I1(_184_),
    .S(_198_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _458_ (.I0(\mem[1][4] ),
    .I1(_185_),
    .S(_198_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _459_ (.I0(\mem[1][5] ),
    .I1(_186_),
    .S(_198_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _460_ (.I0(\mem[1][6] ),
    .I1(_187_),
    .S(_198_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _461_ (.I0(\mem[1][7] ),
    .I1(_188_),
    .S(_198_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _462_ (.A1(_334_),
    .A2(_180_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _463_ (.I0(\mem[2][0] ),
    .I1(_177_),
    .S(_199_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _464_ (.I0(\mem[2][1] ),
    .I1(_182_),
    .S(_199_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _465_ (.I0(\mem[2][2] ),
    .I1(_183_),
    .S(_199_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _466_ (.I0(\mem[2][3] ),
    .I1(_184_),
    .S(_199_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _467_ (.I0(\mem[2][4] ),
    .I1(_185_),
    .S(_199_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _468_ (.I0(\mem[2][5] ),
    .I1(_186_),
    .S(_199_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _469_ (.I0(\mem[2][6] ),
    .I1(_187_),
    .S(_199_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _470_ (.I0(\mem[2][7] ),
    .I1(_188_),
    .S(_199_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _471_ (.A1(_338_),
    .A2(_180_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _472_ (.I0(\mem[3][0] ),
    .I1(_177_),
    .S(_200_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _473_ (.I0(\mem[3][1] ),
    .I1(_182_),
    .S(_200_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _474_ (.I0(\mem[3][2] ),
    .I1(_183_),
    .S(_200_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _475_ (.I0(\mem[3][3] ),
    .I1(_184_),
    .S(_200_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _476_ (.I0(\mem[3][4] ),
    .I1(_185_),
    .S(_200_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _477_ (.I0(\mem[3][5] ),
    .I1(_186_),
    .S(_200_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _478_ (.I0(\mem[3][6] ),
    .I1(_187_),
    .S(_200_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _479_ (.I0(\mem[3][7] ),
    .I1(_188_),
    .S(_200_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _480_ (.A1(net12),
    .A2(_178_),
    .A3(\wr_addr[2] ),
    .A4(_156_),
    .Z(_201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _481_ (.A1(_333_),
    .A2(_201_),
    .Z(_202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _482_ (.I0(\mem[4][0] ),
    .I1(net4),
    .S(_202_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _483_ (.I0(\mem[4][1] ),
    .I1(net5),
    .S(_202_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _484_ (.I0(\mem[4][2] ),
    .I1(net6),
    .S(_202_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _485_ (.I0(\mem[4][3] ),
    .I1(net7),
    .S(_202_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _486_ (.I0(\mem[4][4] ),
    .I1(net8),
    .S(_202_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _487_ (.I0(\mem[4][5] ),
    .I1(net9),
    .S(_202_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _488_ (.I0(\mem[4][6] ),
    .I1(net10),
    .S(_202_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _489_ (.I0(\mem[4][7] ),
    .I1(net11),
    .S(_202_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _490_ (.A1(_336_),
    .A2(_201_),
    .Z(_203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _491_ (.I0(\mem[5][0] ),
    .I1(net4),
    .S(_203_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _492_ (.I0(\mem[5][1] ),
    .I1(net5),
    .S(_203_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _493_ (.I0(\mem[5][2] ),
    .I1(net6),
    .S(_203_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _494_ (.I0(\mem[5][3] ),
    .I1(net7),
    .S(_203_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _495_ (.I0(\mem[5][4] ),
    .I1(net8),
    .S(_203_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _496_ (.I0(\mem[5][5] ),
    .I1(net9),
    .S(_203_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _497_ (.I0(\mem[5][6] ),
    .I1(net10),
    .S(_203_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _498_ (.I0(\mem[5][7] ),
    .I1(net11),
    .S(_203_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _499_ (.A1(_334_),
    .A2(_201_),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _500_ (.I0(\mem[6][0] ),
    .I1(net4),
    .S(_204_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _501_ (.I0(\mem[6][1] ),
    .I1(net5),
    .S(_204_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _502_ (.I0(\mem[6][2] ),
    .I1(net6),
    .S(_204_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _503_ (.I0(\mem[6][3] ),
    .I1(net7),
    .S(_204_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _504_ (.I0(\mem[6][4] ),
    .I1(net8),
    .S(_204_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _505_ (.I0(\mem[6][5] ),
    .I1(net9),
    .S(_204_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _506_ (.I0(\mem[6][6] ),
    .I1(net10),
    .S(_204_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _507_ (.I0(\mem[6][7] ),
    .I1(net11),
    .S(_204_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _508_ (.A1(_338_),
    .A2(_201_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _509_ (.I0(\mem[7][0] ),
    .I1(net4),
    .S(_205_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _510_ (.I0(\mem[7][1] ),
    .I1(net5),
    .S(_205_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _511_ (.I0(\mem[7][2] ),
    .I1(net6),
    .S(_205_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _512_ (.I0(\mem[7][3] ),
    .I1(net7),
    .S(_205_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _513_ (.I0(\mem[7][4] ),
    .I1(net8),
    .S(_205_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _514_ (.I0(\mem[7][5] ),
    .I1(net9),
    .S(_205_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _515_ (.I0(\mem[7][6] ),
    .I1(net10),
    .S(_205_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _516_ (.I0(\mem[7][7] ),
    .I1(net11),
    .S(_205_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _517_ (.A1(_333_),
    .A2(_189_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _518_ (.I0(\mem[8][0] ),
    .I1(net4),
    .S(_206_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _519_ (.I0(\mem[8][1] ),
    .I1(net5),
    .S(_206_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _520_ (.I0(\mem[8][2] ),
    .I1(net6),
    .S(_206_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _521_ (.I0(\mem[8][3] ),
    .I1(net7),
    .S(_206_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _522_ (.I0(\mem[8][4] ),
    .I1(net8),
    .S(_206_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _523_ (.I0(\mem[8][5] ),
    .I1(net9),
    .S(_206_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _524_ (.I0(\mem[8][6] ),
    .I1(net10),
    .S(_206_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _525_ (.I0(\mem[8][7] ),
    .I1(net11),
    .S(_206_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _526_ (.A1(_336_),
    .A2(_189_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _527_ (.I0(\mem[9][0] ),
    .I1(net4),
    .S(_207_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _528_ (.I0(\mem[9][1] ),
    .I1(net5),
    .S(_207_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _529_ (.I0(\mem[9][2] ),
    .I1(net6),
    .S(_207_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _530_ (.I0(\mem[9][3] ),
    .I1(net7),
    .S(_207_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _531_ (.I0(\mem[9][4] ),
    .I1(net8),
    .S(_207_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _532_ (.I0(\mem[9][5] ),
    .I1(net9),
    .S(_207_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _533_ (.I0(\mem[9][6] ),
    .I1(net10),
    .S(_207_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _534_ (.I0(\mem[9][7] ),
    .I1(net11),
    .S(_207_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _535_ (.I(_158_),
    .Z(_208_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _536_ (.I(\rd_addr[2] ),
    .Z(_209_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _537_ (.I0(\mem[1][0] ),
    .I1(\mem[3][0] ),
    .I2(\mem[5][0] ),
    .I3(\mem[7][0] ),
    .S0(_208_),
    .S1(_209_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _538_ (.I(\rd_addr[0] ),
    .Z(_211_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _539_ (.A1(_211_),
    .A2(_323_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _540_ (.I(\rd_addr[0] ),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _541_ (.I(_213_),
    .Z(_214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _542_ (.A1(_214_),
    .A2(_323_),
    .Z(_215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _543_ (.I0(\mem[0][0] ),
    .I1(\mem[2][0] ),
    .I2(\mem[4][0] ),
    .I3(\mem[6][0] ),
    .S0(_158_),
    .S1(\rd_addr[2] ),
    .Z(_216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _544_ (.A1(_210_),
    .A2(_212_),
    .B1(_215_),
    .B2(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _545_ (.A1(\rd_addr[2] ),
    .A2(\rd_addr[3] ),
    .Z(_218_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _546_ (.I(_218_),
    .Z(_219_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _547_ (.A1(\rd_addr[0] ),
    .A2(_219_),
    .Z(_220_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _548_ (.I(_158_),
    .Z(_221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _549_ (.I0(\mem[13][0] ),
    .I1(\mem[15][0] ),
    .S(_221_),
    .Z(_222_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _550_ (.A1(_213_),
    .A2(_161_),
    .A3(_160_),
    .Z(_223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _551_ (.I0(\mem[8][0] ),
    .I1(\mem[10][0] ),
    .S(_221_),
    .Z(_224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _552_ (.A1(_220_),
    .A2(_222_),
    .B1(_223_),
    .B2(_224_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _553_ (.I0(\mem[12][0] ),
    .I1(\mem[14][0] ),
    .S(_221_),
    .Z(_226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _554_ (.A1(_214_),
    .A2(_219_),
    .A3(_226_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _555_ (.I0(\mem[9][0] ),
    .I1(\mem[11][0] ),
    .S(_208_),
    .Z(_228_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _556_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_228_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _557_ (.A1(_217_),
    .A2(_225_),
    .A3(_227_),
    .A4(_229_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _558_ (.I0(\rd_data_reg[0] ),
    .I1(_230_),
    .S(_000_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _559_ (.I0(\mem[1][1] ),
    .I1(\mem[3][1] ),
    .I2(\mem[5][1] ),
    .I3(\mem[7][1] ),
    .S0(_208_),
    .S1(_209_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _560_ (.I(_158_),
    .Z(_232_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _561_ (.I0(\mem[0][1] ),
    .I1(\mem[2][1] ),
    .I2(\mem[4][1] ),
    .I3(\mem[6][1] ),
    .S0(_232_),
    .S1(_209_),
    .Z(_233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _562_ (.A1(_212_),
    .A2(_231_),
    .B1(_233_),
    .B2(_215_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _563_ (.I0(\mem[12][1] ),
    .I1(\mem[14][1] ),
    .S(_159_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _564_ (.A1(_214_),
    .A2(_219_),
    .A3(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _565_ (.I(_158_),
    .Z(_237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _566_ (.I0(\mem[9][1] ),
    .I1(\mem[11][1] ),
    .S(_237_),
    .Z(_238_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _567_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_238_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _568_ (.I0(\mem[8][1] ),
    .I1(\mem[10][1] ),
    .S(_221_),
    .Z(_240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _569_ (.I0(\mem[13][1] ),
    .I1(\mem[15][1] ),
    .S(_237_),
    .Z(_241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _570_ (.A1(_223_),
    .A2(_240_),
    .B1(_241_),
    .B2(_220_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _571_ (.A1(_234_),
    .A2(_236_),
    .A3(_239_),
    .A4(_242_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _572_ (.I0(\rd_data_reg[1] ),
    .I1(_243_),
    .S(_000_),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _573_ (.I0(\mem[1][2] ),
    .I1(\mem[3][2] ),
    .I2(\mem[5][2] ),
    .I3(\mem[7][2] ),
    .S0(_208_),
    .S1(_209_),
    .Z(_244_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _574_ (.I0(\mem[0][2] ),
    .I1(\mem[2][2] ),
    .I2(\mem[4][2] ),
    .I3(\mem[6][2] ),
    .S0(_232_),
    .S1(\rd_addr[2] ),
    .Z(_245_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _575_ (.A1(_212_),
    .A2(_244_),
    .B1(_245_),
    .B2(_215_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _576_ (.I0(\mem[12][2] ),
    .I1(\mem[14][2] ),
    .S(_159_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _577_ (.A1(_214_),
    .A2(_219_),
    .A3(_247_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _578_ (.I0(\mem[9][2] ),
    .I1(\mem[11][2] ),
    .S(_237_),
    .Z(_249_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _579_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_249_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _580_ (.I0(\mem[8][2] ),
    .I1(\mem[10][2] ),
    .S(_221_),
    .Z(_251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _581_ (.I0(\mem[13][2] ),
    .I1(\mem[15][2] ),
    .S(_237_),
    .Z(_252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _582_ (.A1(_223_),
    .A2(_251_),
    .B1(_252_),
    .B2(_220_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _583_ (.A1(_246_),
    .A2(_248_),
    .A3(_250_),
    .A4(_253_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _584_ (.I0(\rd_data_reg[2] ),
    .I1(_254_),
    .S(_000_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _585_ (.I0(\mem[1][3] ),
    .I1(\mem[3][3] ),
    .I2(\mem[5][3] ),
    .I3(\mem[7][3] ),
    .S0(_208_),
    .S1(_209_),
    .Z(_255_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _586_ (.I0(\mem[0][3] ),
    .I1(\mem[2][3] ),
    .I2(\mem[4][3] ),
    .I3(\mem[6][3] ),
    .S0(_232_),
    .S1(\rd_addr[2] ),
    .Z(_256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _587_ (.A1(_212_),
    .A2(_255_),
    .B1(_256_),
    .B2(_215_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _588_ (.I0(\mem[12][3] ),
    .I1(\mem[14][3] ),
    .S(_159_),
    .Z(_258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _589_ (.A1(_214_),
    .A2(_219_),
    .A3(_258_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _590_ (.I0(\mem[9][3] ),
    .I1(\mem[11][3] ),
    .S(_237_),
    .Z(_260_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _591_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_260_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _592_ (.I0(\mem[8][3] ),
    .I1(\mem[10][3] ),
    .S(_221_),
    .Z(_262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _593_ (.I0(\mem[13][3] ),
    .I1(\mem[15][3] ),
    .S(_237_),
    .Z(_263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _594_ (.A1(_223_),
    .A2(_262_),
    .B1(_263_),
    .B2(_220_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _595_ (.A1(_257_),
    .A2(_259_),
    .A3(_261_),
    .A4(_264_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _596_ (.I0(\rd_data_reg[3] ),
    .I1(_265_),
    .S(_000_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _597_ (.I0(\mem[1][4] ),
    .I1(\mem[3][4] ),
    .I2(\mem[5][4] ),
    .I3(\mem[7][4] ),
    .S0(_208_),
    .S1(_209_),
    .Z(_266_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _598_ (.I0(\mem[0][4] ),
    .I1(\mem[2][4] ),
    .I2(\mem[4][4] ),
    .I3(\mem[6][4] ),
    .S0(_232_),
    .S1(\rd_addr[2] ),
    .Z(_267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _599_ (.A1(_212_),
    .A2(_266_),
    .B1(_267_),
    .B2(_215_),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _600_ (.I0(\mem[12][4] ),
    .I1(\mem[14][4] ),
    .S(_159_),
    .Z(_269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _601_ (.A1(_214_),
    .A2(_219_),
    .A3(_269_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _602_ (.I0(\mem[9][4] ),
    .I1(\mem[11][4] ),
    .S(_237_),
    .Z(_271_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _603_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_271_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _604_ (.I0(\mem[8][4] ),
    .I1(\mem[10][4] ),
    .S(_221_),
    .Z(_273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _605_ (.I0(\mem[13][4] ),
    .I1(\mem[15][4] ),
    .S(_208_),
    .Z(_274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _606_ (.A1(_223_),
    .A2(_273_),
    .B1(_274_),
    .B2(_220_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _607_ (.A1(_268_),
    .A2(_270_),
    .A3(_272_),
    .A4(_275_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _608_ (.I0(\rd_data_reg[4] ),
    .I1(_276_),
    .S(_000_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _609_ (.I0(\mem[1][5] ),
    .I1(\mem[3][5] ),
    .I2(\mem[5][5] ),
    .I3(\mem[7][5] ),
    .S0(_232_),
    .S1(_209_),
    .Z(_277_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _610_ (.I0(\mem[0][5] ),
    .I1(\mem[2][5] ),
    .I2(\mem[4][5] ),
    .I3(\mem[6][5] ),
    .S0(_232_),
    .S1(\rd_addr[2] ),
    .Z(_278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _611_ (.A1(_212_),
    .A2(_277_),
    .B1(_278_),
    .B2(_215_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _612_ (.I0(\mem[12][5] ),
    .I1(\mem[14][5] ),
    .S(_159_),
    .Z(_280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _613_ (.A1(_214_),
    .A2(_219_),
    .A3(_280_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _614_ (.I0(\mem[9][5] ),
    .I1(\mem[11][5] ),
    .S(_237_),
    .Z(_282_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _615_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_282_),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _616_ (.I0(\mem[8][5] ),
    .I1(\mem[10][5] ),
    .S(_221_),
    .Z(_284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _617_ (.I0(\mem[13][5] ),
    .I1(\mem[15][5] ),
    .S(_208_),
    .Z(_285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _618_ (.A1(_223_),
    .A2(_284_),
    .B1(_285_),
    .B2(_220_),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _619_ (.A1(_279_),
    .A2(_281_),
    .A3(_283_),
    .A4(_286_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _620_ (.I0(\rd_data_reg[5] ),
    .I1(_287_),
    .S(_000_),
    .Z(_139_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _621_ (.I0(\mem[1][6] ),
    .I1(\mem[3][6] ),
    .I2(\mem[5][6] ),
    .I3(\mem[7][6] ),
    .S0(_232_),
    .S1(_209_),
    .Z(_288_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _622_ (.I0(\mem[0][6] ),
    .I1(\mem[2][6] ),
    .I2(\mem[4][6] ),
    .I3(\mem[6][6] ),
    .S0(_232_),
    .S1(\rd_addr[2] ),
    .Z(_289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _623_ (.A1(_212_),
    .A2(_288_),
    .B1(_289_),
    .B2(_215_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _624_ (.I0(\mem[12][6] ),
    .I1(\mem[14][6] ),
    .S(_159_),
    .Z(_291_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _625_ (.A1(_214_),
    .A2(_219_),
    .A3(_291_),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _626_ (.I0(\mem[9][6] ),
    .I1(\mem[11][6] ),
    .S(_237_),
    .Z(_293_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _627_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_293_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _628_ (.I0(\mem[8][6] ),
    .I1(\mem[10][6] ),
    .S(_221_),
    .Z(_295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _629_ (.I0(\mem[13][6] ),
    .I1(\mem[15][6] ),
    .S(_208_),
    .Z(_296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _630_ (.A1(_223_),
    .A2(_295_),
    .B1(_296_),
    .B2(_220_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _631_ (.A1(_290_),
    .A2(_292_),
    .A3(_294_),
    .A4(_297_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _632_ (.I0(\rd_data_reg[6] ),
    .I1(_298_),
    .S(_000_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _633_ (.I0(\mem[1][7] ),
    .I1(\mem[3][7] ),
    .I2(\mem[5][7] ),
    .I3(\mem[7][7] ),
    .S0(_232_),
    .S1(_209_),
    .Z(_299_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _634_ (.I0(\mem[0][7] ),
    .I1(\mem[2][7] ),
    .I2(\mem[4][7] ),
    .I3(\mem[6][7] ),
    .S0(_232_),
    .S1(\rd_addr[2] ),
    .Z(_300_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _635_ (.A1(_212_),
    .A2(_299_),
    .B1(_300_),
    .B2(_215_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _636_ (.I0(\mem[12][7] ),
    .I1(\mem[14][7] ),
    .S(_159_),
    .Z(_302_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _637_ (.A1(_214_),
    .A2(_219_),
    .A3(_302_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _638_ (.I0(\mem[9][7] ),
    .I1(\mem[11][7] ),
    .S(_237_),
    .Z(_304_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _639_ (.A1(_211_),
    .A2(_326_),
    .A3(_160_),
    .A4(_304_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _640_ (.I0(\mem[8][7] ),
    .I1(\mem[10][7] ),
    .S(_221_),
    .Z(_306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _641_ (.I0(\mem[13][7] ),
    .I1(\mem[15][7] ),
    .S(_208_),
    .Z(_307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _642_ (.A1(_223_),
    .A2(_306_),
    .B1(_307_),
    .B2(_220_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _643_ (.A1(_301_),
    .A2(_303_),
    .A3(_305_),
    .A4(_308_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _644_ (.I0(\rd_data_reg[7] ),
    .I1(_309_),
    .S(_000_),
    .Z(_141_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _645_ (.A1(_214_),
    .A2(_157_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _646_ (.I0(_159_),
    .I1(_001_),
    .S(_000_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _647_ (.A1(_331_),
    .A2(_157_),
    .Z(_310_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _648_ (.A1(_326_),
    .A2(_310_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _649_ (.A1(_211_),
    .A2(_159_),
    .A3(_209_),
    .A4(_157_),
    .Z(_311_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _650_ (.A1(_323_),
    .A2(_311_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _651_ (.A1(_331_),
    .A2(_157_),
    .A3(_219_),
    .Z(_312_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _652_ (.A1(\rd_ptr[4] ),
    .A2(_312_),
    .Z(_146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _653_ (.A1(net12),
    .A2(_156_),
    .ZN(_313_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _654_ (.A1(\wr_addr[0] ),
    .A2(_313_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _655_ (.I0(_003_),
    .I1(\wr_addr[1] ),
    .S(_313_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _656_ (.A1(net12),
    .A2(_338_),
    .A3(_156_),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _657_ (.A1(\wr_addr[2] ),
    .A2(_314_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _658_ (.A1(net12),
    .A2(\wr_addr[0] ),
    .Z(_315_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _659_ (.A1(\wr_addr[2] ),
    .A2(\wr_addr[1] ),
    .A3(_156_),
    .A4(_315_),
    .Z(_316_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _660_ (.A1(_178_),
    .A2(_316_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _661_ (.A1(\wr_ptr[4] ),
    .A2(_197_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _662_ (.A1(\rd_data_reg[0] ),
    .A2(rd_valid),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _663_ (.A1(\rd_data_reg[1] ),
    .A2(rd_valid),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _664_ (.A1(\rd_data_reg[2] ),
    .A2(rd_valid),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _665_ (.A1(\rd_data_reg[3] ),
    .A2(rd_valid),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _666_ (.A1(\rd_data_reg[4] ),
    .A2(rd_valid),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _667_ (.A1(\rd_data_reg[5] ),
    .A2(rd_valid),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _668_ (.A1(\rd_data_reg[6] ),
    .A2(rd_valid),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _669_ (.A1(\rd_data_reg[7] ),
    .A2(rd_valid),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _670_ (.A(_317_),
    .B(\wr_addr[1] ),
    .CI(_318_),
    .CO(_319_),
    .S(_320_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _671_ (.A(_317_),
    .B(\wr_addr[1] ),
    .CO(_321_),
    .S(_322_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _672_ (.A(_323_),
    .B(\wr_addr[3] ),
    .CO(_324_),
    .S(_325_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _673_ (.A(_326_),
    .B(\wr_addr[2] ),
    .CO(_327_),
    .S(_328_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _674_ (.A(\rd_addr[0] ),
    .B(_002_),
    .CO(_329_),
    .S(_330_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _675_ (.A(\rd_addr[0] ),
    .B(\rd_addr[1] ),
    .CO(_331_),
    .S(_001_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _676_ (.A(_002_),
    .B(_332_),
    .CO(_333_),
    .S(_003_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _677_ (.A(_002_),
    .B(\wr_addr[1] ),
    .CO(_334_),
    .S(_335_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _678_ (.A(\wr_addr[0] ),
    .B(_332_),
    .CO(_336_),
    .S(_337_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _679_ (.A(\wr_addr[0] ),
    .B(\wr_addr[1] ),
    .CO(_338_),
    .S(_339_));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \almost_empty_reg$_DFFE_PN1P_  (.D(_004_),
    .SETN(net3),
    .CLK(clknet_4_4_0_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \almost_full_reg$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][0]$_DFFE_PP_  (.D(_006_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][1]$_DFFE_PP_  (.D(_007_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][2]$_DFFE_PP_  (.D(_008_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][3]$_DFFE_PP_  (.D(_009_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][4]$_DFFE_PP_  (.D(_010_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][5]$_DFFE_PP_  (.D(_011_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][6]$_DFFE_PP_  (.D(_012_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][7]$_DFFE_PP_  (.D(_013_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][0]$_DFFE_PP_  (.D(_014_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[10][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][1]$_DFFE_PP_  (.D(_015_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[10][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][2]$_DFFE_PP_  (.D(_016_),
    .CLK(clknet_4_6_0_clk),
    .Q(\mem[10][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][3]$_DFFE_PP_  (.D(_017_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[10][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][4]$_DFFE_PP_  (.D(_018_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[10][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][5]$_DFFE_PP_  (.D(_019_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[10][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][6]$_DFFE_PP_  (.D(_020_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[10][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][7]$_DFFE_PP_  (.D(_021_),
    .CLK(clknet_4_6_0_clk),
    .Q(\mem[10][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][0]$_DFFE_PP_  (.D(_022_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[11][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][1]$_DFFE_PP_  (.D(_023_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[11][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][2]$_DFFE_PP_  (.D(_024_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[11][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][3]$_DFFE_PP_  (.D(_025_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[11][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][4]$_DFFE_PP_  (.D(_026_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[11][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][5]$_DFFE_PP_  (.D(_027_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[11][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][6]$_DFFE_PP_  (.D(_028_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[11][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][7]$_DFFE_PP_  (.D(_029_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[11][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][0]$_DFFE_PP_  (.D(_030_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[12][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][1]$_DFFE_PP_  (.D(_031_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[12][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][2]$_DFFE_PP_  (.D(_032_),
    .CLK(clknet_4_5_0_clk),
    .Q(\mem[12][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][3]$_DFFE_PP_  (.D(_033_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[12][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][4]$_DFFE_PP_  (.D(_034_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[12][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][5]$_DFFE_PP_  (.D(_035_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[12][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][6]$_DFFE_PP_  (.D(_036_),
    .CLK(clknet_4_5_0_clk),
    .Q(\mem[12][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][7]$_DFFE_PP_  (.D(_037_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[12][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][0]$_DFFE_PP_  (.D(_038_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[13][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][1]$_DFFE_PP_  (.D(_039_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[13][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][2]$_DFFE_PP_  (.D(_040_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[13][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][3]$_DFFE_PP_  (.D(_041_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[13][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][4]$_DFFE_PP_  (.D(_042_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[13][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][5]$_DFFE_PP_  (.D(_043_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[13][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][6]$_DFFE_PP_  (.D(_044_),
    .CLK(clknet_4_6_0_clk),
    .Q(\mem[13][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][7]$_DFFE_PP_  (.D(_045_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[13][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][0]$_DFFE_PP_  (.D(_046_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[14][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][1]$_DFFE_PP_  (.D(_047_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[14][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][2]$_DFFE_PP_  (.D(_048_),
    .CLK(clknet_4_5_0_clk),
    .Q(\mem[14][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][3]$_DFFE_PP_  (.D(_049_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[14][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][4]$_DFFE_PP_  (.D(_050_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[14][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][5]$_DFFE_PP_  (.D(_051_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[14][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][6]$_DFFE_PP_  (.D(_052_),
    .CLK(clknet_4_5_0_clk),
    .Q(\mem[14][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][7]$_DFFE_PP_  (.D(_053_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[14][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][0]$_DFFE_PP_  (.D(_054_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[15][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][1]$_DFFE_PP_  (.D(_055_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[15][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][2]$_DFFE_PP_  (.D(_056_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[15][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][3]$_DFFE_PP_  (.D(_057_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[15][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][4]$_DFFE_PP_  (.D(_058_),
    .CLK(clknet_4_15_0_clk),
    .Q(\mem[15][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][5]$_DFFE_PP_  (.D(_059_),
    .CLK(clknet_4_7_0_clk),
    .Q(\mem[15][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][6]$_DFFE_PP_  (.D(_060_),
    .CLK(clknet_4_6_0_clk),
    .Q(\mem[15][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][7]$_DFFE_PP_  (.D(_061_),
    .CLK(clknet_4_13_0_clk),
    .Q(\mem[15][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][0]$_DFFE_PP_  (.D(_062_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][1]$_DFFE_PP_  (.D(_063_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][2]$_DFFE_PP_  (.D(_064_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][3]$_DFFE_PP_  (.D(_065_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][4]$_DFFE_PP_  (.D(_066_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][5]$_DFFE_PP_  (.D(_067_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][6]$_DFFE_PP_  (.D(_068_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][7]$_DFFE_PP_  (.D(_069_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][0]$_DFFE_PP_  (.D(_070_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][1]$_DFFE_PP_  (.D(_071_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][2]$_DFFE_PP_  (.D(_072_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][3]$_DFFE_PP_  (.D(_073_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][4]$_DFFE_PP_  (.D(_074_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][5]$_DFFE_PP_  (.D(_075_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][6]$_DFFE_PP_  (.D(_076_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][7]$_DFFE_PP_  (.D(_077_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][0]$_DFFE_PP_  (.D(_078_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][1]$_DFFE_PP_  (.D(_079_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][2]$_DFFE_PP_  (.D(_080_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][3]$_DFFE_PP_  (.D(_081_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][4]$_DFFE_PP_  (.D(_082_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][5]$_DFFE_PP_  (.D(_083_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][6]$_DFFE_PP_  (.D(_084_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][7]$_DFFE_PP_  (.D(_085_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][0]$_DFFE_PP_  (.D(_086_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][1]$_DFFE_PP_  (.D(_087_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][2]$_DFFE_PP_  (.D(_088_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][3]$_DFFE_PP_  (.D(_089_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][4]$_DFFE_PP_  (.D(_090_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][5]$_DFFE_PP_  (.D(_091_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][6]$_DFFE_PP_  (.D(_092_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][7]$_DFFE_PP_  (.D(_093_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][0]$_DFFE_PP_  (.D(_094_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][1]$_DFFE_PP_  (.D(_095_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][2]$_DFFE_PP_  (.D(_096_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][3]$_DFFE_PP_  (.D(_097_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][4]$_DFFE_PP_  (.D(_098_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][5]$_DFFE_PP_  (.D(_099_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][6]$_DFFE_PP_  (.D(_100_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][7]$_DFFE_PP_  (.D(_101_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][0]$_DFFE_PP_  (.D(_102_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][1]$_DFFE_PP_  (.D(_103_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][2]$_DFFE_PP_  (.D(_104_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][3]$_DFFE_PP_  (.D(_105_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][4]$_DFFE_PP_  (.D(_106_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][5]$_DFFE_PP_  (.D(_107_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][6]$_DFFE_PP_  (.D(_108_),
    .CLK(clknet_4_0_0_clk),
    .Q(\mem[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][7]$_DFFE_PP_  (.D(_109_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][0]$_DFFE_PP_  (.D(_110_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][1]$_DFFE_PP_  (.D(_111_),
    .CLK(clknet_4_11_0_clk),
    .Q(\mem[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][2]$_DFFE_PP_  (.D(_112_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][3]$_DFFE_PP_  (.D(_113_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][4]$_DFFE_PP_  (.D(_114_),
    .CLK(clknet_4_10_0_clk),
    .Q(\mem[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][5]$_DFFE_PP_  (.D(_115_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][6]$_DFFE_PP_  (.D(_116_),
    .CLK(clknet_4_2_0_clk),
    .Q(\mem[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][7]$_DFFE_PP_  (.D(_117_),
    .CLK(clknet_4_8_0_clk),
    .Q(\mem[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][0]$_DFFE_PP_  (.D(_118_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[8][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][1]$_DFFE_PP_  (.D(_119_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[8][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][2]$_DFFE_PP_  (.D(_120_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[8][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][3]$_DFFE_PP_  (.D(_121_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[8][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][4]$_DFFE_PP_  (.D(_122_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[8][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][5]$_DFFE_PP_  (.D(_123_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[8][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][6]$_DFFE_PP_  (.D(_124_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[8][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][7]$_DFFE_PP_  (.D(_125_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[8][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][0]$_DFFE_PP_  (.D(_126_),
    .CLK(clknet_4_12_0_clk),
    .Q(\mem[9][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][1]$_DFFE_PP_  (.D(_127_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[9][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][2]$_DFFE_PP_  (.D(_128_),
    .CLK(clknet_4_1_0_clk),
    .Q(\mem[9][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][3]$_DFFE_PP_  (.D(_129_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[9][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][4]$_DFFE_PP_  (.D(_130_),
    .CLK(clknet_4_14_0_clk),
    .Q(\mem[9][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][5]$_DFFE_PP_  (.D(_131_),
    .CLK(clknet_4_9_0_clk),
    .Q(\mem[9][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][6]$_DFFE_PP_  (.D(_132_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[9][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][7]$_DFFE_PP_  (.D(_133_),
    .CLK(clknet_4_3_0_clk),
    .Q(\mem[9][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[0]$_DFFE_PN0P_  (.D(_134_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\rd_data_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[1]$_DFFE_PN0P_  (.D(_135_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\rd_data_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[2]$_DFFE_PN0P_  (.D(_136_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\rd_data_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[3]$_DFFE_PN0P_  (.D(_137_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\rd_data_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[4]$_DFFE_PN0P_  (.D(_138_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\rd_data_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[5]$_DFFE_PN0P_  (.D(_139_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\rd_data_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[6]$_DFFE_PN0P_  (.D(_140_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\rd_data_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_reg[7]$_DFFE_PN0P_  (.D(_141_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\rd_data_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[0]$_DFFE_PN0P_  (.D(_142_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\rd_addr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[1]$_DFFE_PN0P_  (.D(_143_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\rd_addr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \rd_ptr[2]$_DFFE_PN0P_  (.D(_144_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\rd_addr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[3]$_DFFE_PN0P_  (.D(_145_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\rd_addr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[4]$_DFFE_PN0P_  (.D(_146_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\rd_ptr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \rd_valid$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(rd_valid));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[0]$_DFFE_PN0P_  (.D(_147_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\wr_addr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_148_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\wr_addr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[2]$_DFFE_PN0P_  (.D(_149_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\wr_addr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[3]$_DFFE_PN0P_  (.D(_150_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\wr_addr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[4]$_DFFE_PN0P_  (.D(_151_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\wr_ptr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 hold1 (.I(net3),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Right_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Right_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Right_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Right_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Right_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Right_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Right_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Right_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Right_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Right_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Right_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Right_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Right_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Right_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Right_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Right_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Right_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Right_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Right_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Right_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Right_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Right_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Right_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Right_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Right_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Right_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Right_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Right_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Right_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Right_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Right_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Right_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Right_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Right_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Right_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Right_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Right_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Right_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Right_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Right_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Right_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Right_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Right_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Right_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Right_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Right_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Right_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Right_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Right_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Right_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Right_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Right_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Right_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Right_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Right_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Right_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Right_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Right_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Right_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Right_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Right_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Right_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Right_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_309_Right_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_310_Right_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_311_Right_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_312_Right_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_313_Right_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_314_Right_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_315_Right_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_316_Right_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_317_Right_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_318_Right_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_319_Right_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_320_Right_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_321_Right_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_322_Right_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_323_Right_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_324_Right_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_325_Right_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_326_Right_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_327_Right_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_328_Right_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_329_Right_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_330_Right_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_331_Right_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_332_Right_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_333_Right_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_334_Right_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_335_Right_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_336_Right_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_337_Right_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_338_Right_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_339_Right_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_340_Right_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_341_Right_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_342_Right_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_343_Right_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_344_Right_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_345_Right_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_346_Right_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_347_Right_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_348_Right_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_349_Right_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_350_Right_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_351_Right_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_352_Right_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_353_Right_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_354_Right_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_355_Right_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_356_Right_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_357_Right_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_358_Right_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_359_Right_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_360_Right_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_361_Right_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_362_Right_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_363_Right_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_364_Right_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_365_Right_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_366_Right_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_367_Right_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_368_Right_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_369_Right_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_370_Right_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_371_Right_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_372_Right_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_373_Right_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_374_Right_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_375_Right_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_376_Right_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_377_Right_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_378_Right_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_379_Right_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_380_Right_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_381_Right_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_382_Right_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_383_Right_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_384_Right_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_385_Right_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_386_Right_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_387_Right_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_388_Right_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_389_Right_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_390_Right_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_391_Right_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_392_Right_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_393_Right_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_394_Right_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_395_Right_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_396_Right_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_397_Right_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_398_Right_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_399_Right_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_400_Right_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_401_Right_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_402_Right_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_403_Right_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_404_Right_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_405_Right_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_406_Right_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_407_Right_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_408_Right_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_409_Right_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_410_Right_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_411_Right_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_412_Right_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_413_Right_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_414_Right_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_415_Right_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_416_Right_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_417_Right_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_418_Right_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_419_Right_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_420_Right_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_421_Right_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_422_Right_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_423_Right_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_424_Right_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_425_Right_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_426_Right_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_427_Right_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_428_Right_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_429_Right_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_430_Right_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_431_Right_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_432_Right_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_433_Right_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_434_Right_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_435_Right_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_436_Right_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_437_Right_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_438_Right_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_439_Right_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_440_Right_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_441_Right_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_442_Right_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_469 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_470 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_471 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_472 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_473 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_474 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_475 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_476 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_477 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_478 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_479 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_480 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_481 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_482 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_483 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_484 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_485 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_486 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_487 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_488 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_489 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_490 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_491 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_492 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_493 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_494 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_495 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_496 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_497 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_498 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_499 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_500 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_501 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_502 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_503 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_504 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_505 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_506 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_507 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_508 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_509 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_510 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_511 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_512 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_513 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_514 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_515 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_516 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_517 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_518 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_519 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_520 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_521 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_522 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_523 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_524 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_525 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_526 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_527 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_528 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_529 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_530 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_531 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_532 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_533 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_534 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_535 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_536 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_537 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_538 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_539 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_540 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_541 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_542 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_543 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_544 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_545 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_546 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_547 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_548 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_549 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_550 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_551 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_552 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_553 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_554 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_555 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_556 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_557 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_558 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_559 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_560 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_561 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_562 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_563 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_564 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_565 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_566 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_567 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_568 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_569 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_570 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_571 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_572 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_573 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_574 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_575 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_576 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_577 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_578 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_579 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_580 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_581 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_582 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_583 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_584 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_585 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_586 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_587 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_588 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_589 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_590 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_591 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_592 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_593 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_594 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_595 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_596 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_597 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_598 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_599 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_600 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_601 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_602 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_603 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_604 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_605 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_606 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_607 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_608 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_609 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_610 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_611 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_612 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_613 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_614 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_615 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_616 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_617 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_618 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_619 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_620 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_621 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_622 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_623 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_624 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_625 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_626 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_627 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_628 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_629 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_630 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_631 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_632 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_633 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_634 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_635 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_636 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_637 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_638 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_639 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_640 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_641 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_642 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_643 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_644 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_645 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_646 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_647 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_648 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_649 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_650 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_651 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_652 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_653 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_654 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_655 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_656 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_657 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_658 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_659 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_660 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_661 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_662 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_663 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_664 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_665 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_666 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_667 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_668 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_669 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_670 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_671 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_672 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_673 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_674 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_675 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_676 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_677 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_678 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_679 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_680 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_681 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_682 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_683 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_684 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_685 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_686 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_687 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_688 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Left_689 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Left_690 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Left_691 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Left_692 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Left_693 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Left_694 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Left_695 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Left_696 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Left_697 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Left_698 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Left_699 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Left_700 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Left_701 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Left_702 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Left_703 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Left_704 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Left_705 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Left_706 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Left_707 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Left_708 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Left_709 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Left_710 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Left_711 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Left_712 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Left_713 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Left_714 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Left_715 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Left_716 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Left_717 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Left_718 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Left_719 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Left_720 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Left_721 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Left_722 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Left_723 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Left_724 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Left_725 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Left_726 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Left_727 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Left_728 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Left_729 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Left_730 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Left_731 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Left_732 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Left_733 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Left_734 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Left_735 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Left_736 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Left_737 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Left_738 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Left_739 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Left_740 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Left_741 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Left_742 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Left_743 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Left_744 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Left_745 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Left_746 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Left_747 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Left_748 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Left_749 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Left_750 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Left_751 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_309_Left_752 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_310_Left_753 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_311_Left_754 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_312_Left_755 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_313_Left_756 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_314_Left_757 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_315_Left_758 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_316_Left_759 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_317_Left_760 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_318_Left_761 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_319_Left_762 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_320_Left_763 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_321_Left_764 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_322_Left_765 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_323_Left_766 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_324_Left_767 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_325_Left_768 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_326_Left_769 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_327_Left_770 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_328_Left_771 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_329_Left_772 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_330_Left_773 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_331_Left_774 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_332_Left_775 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_333_Left_776 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_334_Left_777 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_335_Left_778 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_336_Left_779 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_337_Left_780 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_338_Left_781 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_339_Left_782 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_340_Left_783 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_341_Left_784 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_342_Left_785 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_343_Left_786 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_344_Left_787 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_345_Left_788 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_346_Left_789 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_347_Left_790 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_348_Left_791 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_349_Left_792 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_350_Left_793 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_351_Left_794 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_352_Left_795 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_353_Left_796 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_354_Left_797 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_355_Left_798 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_356_Left_799 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_357_Left_800 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_358_Left_801 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_359_Left_802 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_360_Left_803 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_361_Left_804 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_362_Left_805 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_363_Left_806 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_364_Left_807 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_365_Left_808 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_366_Left_809 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_367_Left_810 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_368_Left_811 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_369_Left_812 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_370_Left_813 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_371_Left_814 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_372_Left_815 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_373_Left_816 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_374_Left_817 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_375_Left_818 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_376_Left_819 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_377_Left_820 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_378_Left_821 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_379_Left_822 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_380_Left_823 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_381_Left_824 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_382_Left_825 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_383_Left_826 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_384_Left_827 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_385_Left_828 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_386_Left_829 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_387_Left_830 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_388_Left_831 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_389_Left_832 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_390_Left_833 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_391_Left_834 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_392_Left_835 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_393_Left_836 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_394_Left_837 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_395_Left_838 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_396_Left_839 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_397_Left_840 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_398_Left_841 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_399_Left_842 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_400_Left_843 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_401_Left_844 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_402_Left_845 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_403_Left_846 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_404_Left_847 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_405_Left_848 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_406_Left_849 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_407_Left_850 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_408_Left_851 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_409_Left_852 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_410_Left_853 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_411_Left_854 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_412_Left_855 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_413_Left_856 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_414_Left_857 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_415_Left_858 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_416_Left_859 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_417_Left_860 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_418_Left_861 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_419_Left_862 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_420_Left_863 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_421_Left_864 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_422_Left_865 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_423_Left_866 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_424_Left_867 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_425_Left_868 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_426_Left_869 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_427_Left_870 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_428_Left_871 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_429_Left_872 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_430_Left_873 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_431_Left_874 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_432_Left_875 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_433_Left_876 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_434_Left_877 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_435_Left_878 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_436_Left_879 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_437_Left_880 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_438_Left_881 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_439_Left_882 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_440_Left_883 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_441_Left_884 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_442_Left_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_2645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_2678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_2689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_2700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_2711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_2722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_2733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_2744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_2755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_2766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_2777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_2799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_2810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_2821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_2843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_2854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_2865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_2876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_2887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_2898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_2909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_3525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_3536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_3547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_3569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_3580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_3591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_3602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_3613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_3624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_3635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_3646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_3657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_3668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_3679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_3701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_3712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_3723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_3734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_3745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_3756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_3767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_3778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_3789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_3800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_3811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_3822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_3833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_3844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_3855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_3866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_3877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_3888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_3899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_3910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_3921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_3943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_3954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_3965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_3976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_3987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_3998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_3999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_4405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_4427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_4438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_4449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_4460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_4471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_4482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_4493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_4504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_4515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_4526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_4537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_4570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_4581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_4592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_4603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_4614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_4625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_4636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_4647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_4658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_4669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_4680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_4691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_4702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_4713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_4724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_4735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_4746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_4757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_4768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_4779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_4790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_4801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_4812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_4823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_4834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_4845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_4856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_4867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_4878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_4889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_4900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_4911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_4922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_4933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_4944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_4955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_4966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_4977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_4988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_4999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_5285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_5296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_5307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_5318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_5329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_5340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_5351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_5362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_5373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_5384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_5395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_5406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_5417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_5428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_5439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_5450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_5461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_5472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_5483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_5494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_5505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_5516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_5527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_5538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_5549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_5560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_5571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_5582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_5593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_5604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_5615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_5626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_5637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_5648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_5659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_5670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_5681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_5692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_5703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_5714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_5725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_5736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_5747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_5758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_5780 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(rd_en),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input2 (.I(net25),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input3 (.I(wr_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input4 (.I(wr_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input5 (.I(wr_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input6 (.I(wr_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input7 (.I(wr_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input8 (.I(wr_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input9 (.I(wr_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input10 (.I(wr_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input11 (.I(wr_en),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(almost_empty));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(almost_full));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(empty));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(full));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rd_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rd_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rd_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rd_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rd_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(rd_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(rd_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(rd_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload0 (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload1 (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload2 (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload3 (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload4 (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload5 (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload6 (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload7 (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload8 (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload9 (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload10 (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload11 (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload12 (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload13 (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 clkload14 (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net4));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net4));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net4));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_4 (.I(net4));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_5 (.I(net6));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_6 (.I(net13));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_7 (.I(net13));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_2473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_2304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_2289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_3957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_3989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_3934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_3942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_3948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_3979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_3965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_3981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_3989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_236_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_246_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_247_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_256_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_256_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_259_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_260_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_262_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_266_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_266_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_268_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_272_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_275_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_276_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_278_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_279_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_280_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_281_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_281_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_282_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_282_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_283_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_284_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_284_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_284_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_285_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_285_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_286_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_286_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_286_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_287_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_287_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_287_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_288_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_288_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_289_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_289_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_290_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_290_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_291_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_291_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_291_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_292_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_292_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_292_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_293_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_293_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_293_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_294_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_294_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_294_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_294_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_294_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_295_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_295_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_295_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_296_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_296_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_296_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_296_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_296_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_297_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_297_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_297_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_298_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_298_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_298_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_298_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_298_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_299_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_299_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_299_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_300_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_300_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_300_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_300_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_300_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_301_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_301_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_301_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_302_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_302_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_302_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_302_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_302_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_303_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_303_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_303_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_304_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_304_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_304_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_304_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_304_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_305_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_305_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_305_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_306_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_306_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_306_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_306_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_306_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_307_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_307_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_307_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_308_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_309_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_309_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_309_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_310_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_310_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_310_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_310_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_310_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_311_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_311_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_311_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_312_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_312_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_312_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_312_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_312_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_313_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_313_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_313_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_314_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_314_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_314_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_314_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_314_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_315_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_315_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_315_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_316_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_316_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_316_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_316_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_316_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_317_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_317_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_317_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_318_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_318_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_318_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_318_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_318_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_319_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_319_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_319_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_320_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_320_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_320_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_320_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_320_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_321_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_321_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_321_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_322_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_322_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_322_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_322_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_322_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_323_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_323_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_323_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_324_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_324_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_324_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_324_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_324_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_325_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_325_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_325_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_326_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_326_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_326_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_326_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_326_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_327_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_327_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_327_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_328_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_328_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_328_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_328_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_328_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_329_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_329_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_329_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_330_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_330_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_330_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_330_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_330_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_331_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_331_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_331_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_332_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_332_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_332_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_332_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_332_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_333_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_333_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_333_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_334_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_334_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_334_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_334_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_334_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_335_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_335_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_335_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_336_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_336_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_336_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_336_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_336_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_337_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_337_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_337_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_338_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_338_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_338_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_338_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_338_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_339_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_339_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_339_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_340_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_340_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_340_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_340_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_340_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_341_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_341_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_341_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_342_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_342_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_342_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_342_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_342_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_343_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_343_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_343_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_344_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_344_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_344_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_344_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_344_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_345_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_345_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_345_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_346_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_346_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_346_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_346_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_346_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_347_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_347_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_347_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_348_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_348_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_348_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_348_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_348_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_349_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_349_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_349_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_350_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_350_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_350_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_350_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_350_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_351_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_351_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_351_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_352_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_352_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_352_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_352_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_352_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_353_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_353_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_353_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_354_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_354_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_354_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_354_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_354_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_355_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_355_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_355_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_356_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_356_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_356_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_356_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_356_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_357_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_357_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_357_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_358_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_358_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_358_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_358_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_358_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_359_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_359_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_359_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_360_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_360_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_360_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_360_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_360_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_361_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_361_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_361_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_362_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_362_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_362_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_362_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_362_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_363_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_363_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_363_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_364_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_364_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_364_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_364_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_364_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_365_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_365_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_365_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_366_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_366_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_366_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_366_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_366_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_367_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_367_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_367_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_368_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_368_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_368_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_368_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_368_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_369_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_369_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_369_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_370_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_370_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_370_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_370_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_370_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_371_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_371_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_371_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_372_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_372_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_372_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_372_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_372_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_373_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_373_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_373_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_374_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_374_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_374_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_374_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_374_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_375_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_375_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_375_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_376_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_376_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_376_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_376_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_376_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_377_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_377_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_377_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_378_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_378_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_378_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_378_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_378_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_379_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_379_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_379_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_380_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_380_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_380_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_380_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_380_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_381_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_381_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_381_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_382_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_382_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_382_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_382_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_382_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_383_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_383_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_383_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_384_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_384_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_384_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_384_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_384_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_385_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_385_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_385_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_386_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_386_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_386_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_386_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_386_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_387_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_387_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_387_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_388_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_388_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_388_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_388_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_388_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_389_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_389_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_389_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_390_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_390_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_390_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_390_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_390_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_391_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_391_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_391_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_392_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_392_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_392_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_392_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_392_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_393_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_393_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_393_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_394_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_394_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_394_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_394_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_394_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_395_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_395_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_395_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_396_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_396_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_396_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_396_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_396_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_397_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_397_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_397_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_398_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_398_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_398_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_398_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_398_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_399_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_399_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_399_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_400_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_400_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_400_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_400_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_400_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_401_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_401_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_401_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_402_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_402_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_402_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_402_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_402_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_403_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_403_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_403_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_404_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_404_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_404_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_404_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_404_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_405_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_405_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_405_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_406_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_406_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_406_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_406_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_406_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_407_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_407_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_407_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_408_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_408_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_408_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_408_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_408_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_409_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_409_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_409_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_410_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_410_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_410_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_410_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_410_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_411_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_411_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_411_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_412_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_412_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_412_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_412_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_412_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_413_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_413_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_413_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_414_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_414_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_414_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_414_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_414_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_415_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_415_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_415_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_416_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_416_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_416_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_416_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_416_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_417_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_417_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_417_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_418_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_418_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_418_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_418_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_418_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_419_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_419_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_419_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_420_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_420_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_420_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_420_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_420_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_421_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_421_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_421_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_422_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_422_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_422_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_422_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_422_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_423_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_423_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_423_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_424_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_424_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_424_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_424_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_424_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_425_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_425_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_425_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_426_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_426_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_426_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_426_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_426_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_427_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_427_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_427_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_428_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_428_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_428_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_428_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_428_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_429_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_429_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_429_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_430_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_430_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_430_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_430_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_430_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_431_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_431_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_431_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_432_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_432_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_432_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_432_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_432_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_433_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_433_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_433_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_434_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_434_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_434_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_434_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_434_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_435_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_435_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_435_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_436_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_436_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_436_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_436_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_436_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_437_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_437_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_437_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_438_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_438_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_438_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_438_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_438_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_439_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_439_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_439_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_440_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_440_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_440_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_440_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_440_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_440_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_440_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_440_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_440_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_440_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_441_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_441_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_441_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_441_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_441_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_441_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_442_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_442_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_442_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_3010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_3188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_3366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_3544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_3722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_3900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_442_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_442_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_442_3994 ();
endmodule
