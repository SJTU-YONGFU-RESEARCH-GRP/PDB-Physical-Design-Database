module mesh_router (clk,
    east_in_ready,
    east_in_valid,
    east_out_ready,
    east_out_valid,
    local_in_ready,
    local_in_valid,
    local_out_ready,
    local_out_valid,
    north_in_ready,
    north_in_valid,
    north_out_ready,
    north_out_valid,
    rst_n,
    south_in_ready,
    south_in_valid,
    south_out_ready,
    south_out_valid,
    west_in_ready,
    west_in_valid,
    west_out_ready,
    west_out_valid,
    east_in_data,
    east_out_data,
    local_in_data,
    local_out_data,
    north_in_data,
    north_out_data,
    south_in_data,
    south_out_data,
    west_in_data,
    west_out_data);
 input clk;
 output east_in_ready;
 input east_in_valid;
 input east_out_ready;
 output east_out_valid;
 output local_in_ready;
 input local_in_valid;
 input local_out_ready;
 output local_out_valid;
 output north_in_ready;
 input north_in_valid;
 input north_out_ready;
 output north_out_valid;
 input rst_n;
 output south_in_ready;
 input south_in_valid;
 input south_out_ready;
 output south_out_valid;
 output west_in_ready;
 input west_in_valid;
 input west_out_ready;
 output west_out_valid;
 input [31:0] east_in_data;
 output [31:0] east_out_data;
 input [31:0] local_in_data;
 output [31:0] local_out_data;
 input [31:0] north_in_data;
 output [31:0] north_out_data;
 input [31:0] south_in_data;
 output [31:0] south_out_data;
 input [31:0] west_in_data;
 output [31:0] west_out_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire clknet_0_clk;
 wire \dest_id[0][0] ;
 wire \dest_id[0][1] ;
 wire \dest_id[0][2] ;
 wire \dest_id[0][3] ;
 wire \dest_id[0][4] ;
 wire \dest_id[0][5] ;
 wire \dest_id[0][6] ;
 wire \dest_id[0][7] ;
 wire \dest_id[1][0] ;
 wire \dest_id[1][1] ;
 wire \dest_id[1][2] ;
 wire \dest_id[1][3] ;
 wire \dest_id[1][4] ;
 wire \dest_id[1][5] ;
 wire \dest_id[1][6] ;
 wire \dest_id[1][7] ;
 wire \dest_id[2][0] ;
 wire \dest_id[2][1] ;
 wire \dest_id[2][2] ;
 wire \dest_id[2][3] ;
 wire \dest_id[2][4] ;
 wire \dest_id[2][5] ;
 wire \dest_id[2][6] ;
 wire \dest_id[2][7] ;
 wire \dest_id[3][0] ;
 wire \dest_id[3][1] ;
 wire \dest_id[3][2] ;
 wire \dest_id[3][3] ;
 wire \dest_id[3][4] ;
 wire \dest_id[3][5] ;
 wire \dest_id[3][6] ;
 wire \dest_id[3][7] ;
 wire \dest_id[4][0] ;
 wire \dest_id[4][1] ;
 wire \dest_id[4][2] ;
 wire \dest_id[4][3] ;
 wire \dest_id[4][4] ;
 wire \dest_id[4][5] ;
 wire \dest_id[4][6] ;
 wire \dest_id[4][7] ;
 wire \input_buffer[0][0] ;
 wire \input_buffer[0][10] ;
 wire \input_buffer[0][11] ;
 wire \input_buffer[0][12] ;
 wire \input_buffer[0][13] ;
 wire \input_buffer[0][14] ;
 wire \input_buffer[0][15] ;
 wire \input_buffer[0][16] ;
 wire \input_buffer[0][17] ;
 wire \input_buffer[0][18] ;
 wire \input_buffer[0][19] ;
 wire \input_buffer[0][1] ;
 wire \input_buffer[0][20] ;
 wire \input_buffer[0][21] ;
 wire \input_buffer[0][22] ;
 wire \input_buffer[0][23] ;
 wire \input_buffer[0][2] ;
 wire \input_buffer[0][3] ;
 wire \input_buffer[0][4] ;
 wire \input_buffer[0][5] ;
 wire \input_buffer[0][6] ;
 wire \input_buffer[0][7] ;
 wire \input_buffer[0][8] ;
 wire \input_buffer[0][9] ;
 wire \input_buffer[1][0] ;
 wire \input_buffer[1][10] ;
 wire \input_buffer[1][11] ;
 wire \input_buffer[1][12] ;
 wire \input_buffer[1][13] ;
 wire \input_buffer[1][14] ;
 wire \input_buffer[1][15] ;
 wire \input_buffer[1][16] ;
 wire \input_buffer[1][17] ;
 wire \input_buffer[1][18] ;
 wire \input_buffer[1][19] ;
 wire \input_buffer[1][1] ;
 wire \input_buffer[1][20] ;
 wire \input_buffer[1][21] ;
 wire \input_buffer[1][22] ;
 wire \input_buffer[1][23] ;
 wire \input_buffer[1][2] ;
 wire \input_buffer[1][3] ;
 wire \input_buffer[1][4] ;
 wire \input_buffer[1][5] ;
 wire \input_buffer[1][6] ;
 wire \input_buffer[1][7] ;
 wire \input_buffer[1][8] ;
 wire \input_buffer[1][9] ;
 wire \input_buffer[2][0] ;
 wire \input_buffer[2][10] ;
 wire \input_buffer[2][11] ;
 wire \input_buffer[2][12] ;
 wire \input_buffer[2][13] ;
 wire \input_buffer[2][14] ;
 wire \input_buffer[2][15] ;
 wire \input_buffer[2][16] ;
 wire \input_buffer[2][17] ;
 wire \input_buffer[2][18] ;
 wire \input_buffer[2][19] ;
 wire \input_buffer[2][1] ;
 wire \input_buffer[2][20] ;
 wire \input_buffer[2][21] ;
 wire \input_buffer[2][22] ;
 wire \input_buffer[2][23] ;
 wire \input_buffer[2][2] ;
 wire \input_buffer[2][3] ;
 wire \input_buffer[2][4] ;
 wire \input_buffer[2][5] ;
 wire \input_buffer[2][6] ;
 wire \input_buffer[2][7] ;
 wire \input_buffer[2][8] ;
 wire \input_buffer[2][9] ;
 wire \input_buffer[3][0] ;
 wire \input_buffer[3][10] ;
 wire \input_buffer[3][11] ;
 wire \input_buffer[3][12] ;
 wire \input_buffer[3][13] ;
 wire \input_buffer[3][14] ;
 wire \input_buffer[3][15] ;
 wire \input_buffer[3][16] ;
 wire \input_buffer[3][17] ;
 wire \input_buffer[3][18] ;
 wire \input_buffer[3][19] ;
 wire \input_buffer[3][1] ;
 wire \input_buffer[3][20] ;
 wire \input_buffer[3][21] ;
 wire \input_buffer[3][22] ;
 wire \input_buffer[3][23] ;
 wire \input_buffer[3][2] ;
 wire \input_buffer[3][3] ;
 wire \input_buffer[3][4] ;
 wire \input_buffer[3][5] ;
 wire \input_buffer[3][6] ;
 wire \input_buffer[3][7] ;
 wire \input_buffer[3][8] ;
 wire \input_buffer[3][9] ;
 wire \input_buffer[4][0] ;
 wire \input_buffer[4][10] ;
 wire \input_buffer[4][11] ;
 wire \input_buffer[4][12] ;
 wire \input_buffer[4][13] ;
 wire \input_buffer[4][14] ;
 wire \input_buffer[4][15] ;
 wire \input_buffer[4][16] ;
 wire \input_buffer[4][17] ;
 wire \input_buffer[4][18] ;
 wire \input_buffer[4][19] ;
 wire \input_buffer[4][1] ;
 wire \input_buffer[4][20] ;
 wire \input_buffer[4][21] ;
 wire \input_buffer[4][22] ;
 wire \input_buffer[4][23] ;
 wire \input_buffer[4][2] ;
 wire \input_buffer[4][3] ;
 wire \input_buffer[4][4] ;
 wire \input_buffer[4][5] ;
 wire \input_buffer[4][6] ;
 wire \input_buffer[4][7] ;
 wire \input_buffer[4][8] ;
 wire \input_buffer[4][9] ;
 wire \input_buffer_valid[0] ;
 wire \input_buffer_valid[1] ;
 wire \input_buffer_valid[2] ;
 wire \input_buffer_valid[3] ;
 wire \input_buffer_valid[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;

 sky130_fd_sc_hd__inv_1 _1163_ (.A(\input_buffer_valid[4] ),
    .Y(net203));
 sky130_fd_sc_hd__and3_4 _1164_ (.A(net203),
    .B(net68),
    .C(net104),
    .X(_0005_));
 sky130_fd_sc_hd__buf_4 _1165_ (.A(\input_buffer_valid[3] ),
    .X(_0597_));
 sky130_fd_sc_hd__clkinv_2 _1166_ (.A(_0597_),
    .Y(net301));
 sky130_fd_sc_hd__and3_4 _1167_ (.A(net104),
    .B(net301),
    .C(net171),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _1168_ (.A(\input_buffer_valid[2] ),
    .X(_0598_));
 sky130_fd_sc_hd__buf_2 _1169_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__inv_1 _1170_ (.A(_0599_),
    .Y(net271));
 sky130_fd_sc_hd__and3_4 _1171_ (.A(net104),
    .B(net271),
    .C(net137),
    .X(_0007_));
 sky130_fd_sc_hd__buf_4 _1172_ (.A(\input_buffer_valid[1] ),
    .X(_0600_));
 sky130_fd_sc_hd__buf_2 _1173_ (.A(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__buf_2 _1174_ (.A(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__inv_1 _1175_ (.A(_0602_),
    .Y(net173));
 sky130_fd_sc_hd__and3_4 _1176_ (.A(net104),
    .B(net173),
    .C(net34),
    .X(_0008_));
 sky130_fd_sc_hd__buf_2 _1177_ (.A(\input_buffer_valid[0] ),
    .X(_0603_));
 sky130_fd_sc_hd__clkinvlp_4 _1178_ (.A(_0603_),
    .Y(net237));
 sky130_fd_sc_hd__and3_4 _1179_ (.A(net104),
    .B(net237),
    .C(net102),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_4 _1180_ (.A(\dest_id[4][1] ),
    .X(_0604_));
 sky130_fd_sc_hd__buf_4 _1181_ (.A(\dest_id[4][2] ),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_4 _1182_ (.A(\dest_id[4][0] ),
    .X(_0606_));
 sky130_fd_sc_hd__nor3b_2 _1183_ (.A(_0604_),
    .B(_0605_),
    .C_N(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__clkbuf_4 _1184_ (.A(\dest_id[4][3] ),
    .X(_0608_));
 sky130_fd_sc_hd__nor3b_2 _1185_ (.A(_0606_),
    .B(_0608_),
    .C_N(_0605_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor4_2 _1186_ (.A(\dest_id[4][5] ),
    .B(\dest_id[4][4] ),
    .C(\dest_id[4][7] ),
    .D(\dest_id[4][6] ),
    .Y(_0610_));
 sky130_fd_sc_hd__o21ai_2 _1187_ (.A1(_0607_),
    .A2(_0609_),
    .B1(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_1 _1188_ (.A(_0611_),
    .Y(_1159_));
 sky130_fd_sc_hd__or4_1 _1189_ (.A(\dest_id[4][5] ),
    .B(\dest_id[4][4] ),
    .C(\dest_id[4][7] ),
    .D(\dest_id[4][6] ),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_4 _1190_ (.A(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__or3b_1 _1191_ (.A(\dest_id[4][0] ),
    .B(_0608_),
    .C_N(_0605_),
    .X(_0614_));
 sky130_fd_sc_hd__buf_4 _1192_ (.A(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_2 _1193_ (.A(_0613_),
    .B(_0615_),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_1 _1194_ (.A(_1148_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand3b_1 _1195_ (.A_N(_0605_),
    .B(_0608_),
    .C(_0606_),
    .Y(_0616_));
 sky130_fd_sc_hd__a211o_1 _1196_ (.A1(_0615_),
    .A2(_0616_),
    .B1(_0604_),
    .C1(_0613_),
    .X(_1147_));
 sky130_fd_sc_hd__inv_1 _1197_ (.A(_1147_),
    .Y(_1154_));
 sky130_fd_sc_hd__a221oi_1 _1198_ (.A1(net172),
    .A2(_0609_),
    .B1(_1151_),
    .B2(net138),
    .C1(_1147_),
    .Y(_0617_));
 sky130_fd_sc_hd__or3b_1 _1199_ (.A(_0604_),
    .B(_0605_),
    .C_N(\dest_id[4][0] ),
    .X(_0618_));
 sky130_fd_sc_hd__buf_2 _1200_ (.A(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__nand3b_1 _1201_ (.A_N(_0606_),
    .B(_0604_),
    .C(_0605_),
    .Y(_0620_));
 sky130_fd_sc_hd__a211oi_2 _1202_ (.A1(_0619_),
    .A2(_0620_),
    .B1(_0608_),
    .C1(_0613_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2_1 _1203_ (.A(net103),
    .B(_1151_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _1204_ (.A(net35),
    .B(_1148_),
    .Y(_0623_));
 sky130_fd_sc_hd__and3_1 _1205_ (.A(_0621_),
    .B(_0622_),
    .C(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__buf_4 _1206_ (.A(\input_buffer_valid[4] ),
    .X(_0625_));
 sky130_fd_sc_hd__o21ai_0 _1207_ (.A1(net69),
    .A2(_1159_),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__o32a_1 _1208_ (.A1(_0617_),
    .A2(_0624_),
    .A3(_0626_),
    .B1(net68),
    .B2(_0625_),
    .X(_0004_));
 sky130_fd_sc_hd__buf_4 _1209_ (.A(\dest_id[3][1] ),
    .X(_0627_));
 sky130_fd_sc_hd__buf_4 _1210_ (.A(\dest_id[3][2] ),
    .X(_0628_));
 sky130_fd_sc_hd__or3b_2 _1211_ (.A(_0627_),
    .B(_0628_),
    .C_N(\dest_id[3][0] ),
    .X(_0629_));
 sky130_fd_sc_hd__or3b_2 _1212_ (.A(\dest_id[3][0] ),
    .B(\dest_id[3][3] ),
    .C_N(\dest_id[3][2] ),
    .X(_0630_));
 sky130_fd_sc_hd__or4_2 _1213_ (.A(\dest_id[3][5] ),
    .B(\dest_id[3][4] ),
    .C(\dest_id[3][7] ),
    .D(\dest_id[3][6] ),
    .X(_0631_));
 sky130_fd_sc_hd__a21oi_4 _1214_ (.A1(_0629_),
    .A2(_0630_),
    .B1(_0631_),
    .Y(_1144_));
 sky130_fd_sc_hd__nor2_1 _1215_ (.A(_0631_),
    .B(_0630_),
    .Y(_1133_));
 sky130_fd_sc_hd__inv_1 _1216_ (.A(_1133_),
    .Y(_1136_));
 sky130_fd_sc_hd__inv_1 _1217_ (.A(_0627_),
    .Y(_0632_));
 sky130_fd_sc_hd__nor4_4 _1218_ (.A(\dest_id[3][5] ),
    .B(\dest_id[3][4] ),
    .C(\dest_id[3][7] ),
    .D(\dest_id[3][6] ),
    .Y(_0633_));
 sky130_fd_sc_hd__buf_4 _1219_ (.A(\dest_id[3][0] ),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _1220_ (.A(_0634_),
    .B(\dest_id[3][3] ),
    .Y(_0635_));
 sky130_fd_sc_hd__o21ai_0 _1221_ (.A1(_0628_),
    .A2(_0635_),
    .B1(_0630_),
    .Y(_0636_));
 sky130_fd_sc_hd__and3_1 _1222_ (.A(_0632_),
    .B(_0633_),
    .C(_0636_),
    .X(_1139_));
 sky130_fd_sc_hd__buf_2 _1223_ (.A(_0597_),
    .X(_0637_));
 sky130_fd_sc_hd__nor4_1 _1224_ (.A(_1145_),
    .B(_1134_),
    .C(_1140_),
    .D(_1142_),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_1 _1225_ (.A(net69),
    .B(_1144_),
    .Y(_0639_));
 sky130_fd_sc_hd__a21oi_1 _1226_ (.A1(_1144_),
    .A2(_0638_),
    .B1(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(net138),
    .B(_0630_),
    .Y(_0641_));
 sky130_fd_sc_hd__nor3b_4 _1228_ (.A(_0634_),
    .B(\dest_id[3][3] ),
    .C_N(_0628_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand2_1 _1229_ (.A(net172),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nor2_1 _1230_ (.A(\dest_id[3][3] ),
    .B(_0631_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2b_1 _1231_ (.A_N(_0634_),
    .B(_0628_),
    .Y(_0645_));
 sky130_fd_sc_hd__o32ai_1 _1232_ (.A1(net35),
    .A2(_0632_),
    .A3(_0645_),
    .B1(_0629_),
    .B2(net103),
    .Y(_0646_));
 sky130_fd_sc_hd__a32oi_1 _1233_ (.A1(_1139_),
    .A2(_0641_),
    .A3(_0643_),
    .B1(_0644_),
    .B2(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(_0637_),
    .B(net171),
    .Y(_0648_));
 sky130_fd_sc_hd__a31oi_1 _1235_ (.A1(_0637_),
    .A2(_0640_),
    .A3(_0647_),
    .B1(_0648_),
    .Y(_0003_));
 sky130_fd_sc_hd__buf_4 _1236_ (.A(\dest_id[2][2] ),
    .X(_0649_));
 sky130_fd_sc_hd__buf_4 _1237_ (.A(\dest_id[2][0] ),
    .X(_0650_));
 sky130_fd_sc_hd__nor3b_4 _1238_ (.A(\dest_id[2][1] ),
    .B(_0649_),
    .C_N(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__clkbuf_4 _1239_ (.A(\dest_id[2][3] ),
    .X(_0652_));
 sky130_fd_sc_hd__nor3b_2 _1240_ (.A(_0650_),
    .B(_0652_),
    .C_N(_0649_),
    .Y(_0653_));
 sky130_fd_sc_hd__nor4_4 _1241_ (.A(\dest_id[2][5] ),
    .B(\dest_id[2][4] ),
    .C(\dest_id[2][7] ),
    .D(\dest_id[2][6] ),
    .Y(_0654_));
 sky130_fd_sc_hd__o21ai_4 _1242_ (.A1(_0651_),
    .A2(_0653_),
    .B1(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__inv_1 _1243_ (.A(_0655_),
    .Y(_1129_));
 sky130_fd_sc_hd__or4_4 _1244_ (.A(\dest_id[2][5] ),
    .B(\dest_id[2][4] ),
    .C(\dest_id[2][7] ),
    .D(\dest_id[2][6] ),
    .X(_0656_));
 sky130_fd_sc_hd__or3b_1 _1245_ (.A(\dest_id[2][0] ),
    .B(_0652_),
    .C_N(\dest_id[2][2] ),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_2 _1246_ (.A(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(_0656_),
    .B(_0658_),
    .Y(_1118_));
 sky130_fd_sc_hd__inv_1 _1248_ (.A(_1118_),
    .Y(_1121_));
 sky130_fd_sc_hd__inv_1 _1249_ (.A(\dest_id[2][1] ),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(_0650_),
    .B(_0652_),
    .Y(_0660_));
 sky130_fd_sc_hd__o21ai_0 _1251_ (.A1(_0649_),
    .A2(_0660_),
    .B1(_0658_),
    .Y(_0661_));
 sky130_fd_sc_hd__and3_1 _1252_ (.A(_0659_),
    .B(_0654_),
    .C(_0661_),
    .X(_1124_));
 sky130_fd_sc_hd__nor4_1 _1253_ (.A(_1130_),
    .B(_1119_),
    .C(_1125_),
    .D(_1127_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _1254_ (.A(net69),
    .B(_0655_),
    .Y(_0663_));
 sky130_fd_sc_hd__o21ai_0 _1255_ (.A1(_0655_),
    .A2(_0662_),
    .B1(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _1256_ (.A(net138),
    .B(_0658_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(net172),
    .B(_0653_),
    .Y(_0666_));
 sky130_fd_sc_hd__nor2_1 _1258_ (.A(_0652_),
    .B(_0656_),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2b_1 _1259_ (.A_N(_0650_),
    .B(_0649_),
    .Y(_0668_));
 sky130_fd_sc_hd__or3b_2 _1260_ (.A(\dest_id[2][1] ),
    .B(_0649_),
    .C_N(_0650_),
    .X(_0669_));
 sky130_fd_sc_hd__o32ai_1 _1261_ (.A1(net35),
    .A2(_0659_),
    .A3(_0668_),
    .B1(_0669_),
    .B2(net103),
    .Y(_0670_));
 sky130_fd_sc_hd__a32oi_1 _1262_ (.A1(_1124_),
    .A2(_0665_),
    .A3(_0666_),
    .B1(_0667_),
    .B2(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor2_1 _1263_ (.A(_0599_),
    .B(net137),
    .Y(_0672_));
 sky130_fd_sc_hd__a31oi_1 _1264_ (.A1(_0599_),
    .A2(_0664_),
    .A3(_0671_),
    .B1(_0672_),
    .Y(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _1265_ (.A(\dest_id[1][1] ),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_4 _1266_ (.A(\dest_id[1][2] ),
    .X(_0674_));
 sky130_fd_sc_hd__nor3b_2 _1267_ (.A(_0673_),
    .B(_0674_),
    .C_N(\dest_id[1][0] ),
    .Y(_0675_));
 sky130_fd_sc_hd__clkbuf_4 _1268_ (.A(\dest_id[1][0] ),
    .X(_0676_));
 sky130_fd_sc_hd__buf_4 _1269_ (.A(\dest_id[1][3] ),
    .X(_0677_));
 sky130_fd_sc_hd__nor3b_2 _1270_ (.A(_0676_),
    .B(_0677_),
    .C_N(\dest_id[1][2] ),
    .Y(_0678_));
 sky130_fd_sc_hd__nor4_2 _1271_ (.A(\dest_id[1][5] ),
    .B(\dest_id[1][4] ),
    .C(\dest_id[1][7] ),
    .D(\dest_id[1][6] ),
    .Y(_0679_));
 sky130_fd_sc_hd__o21ai_2 _1272_ (.A1(_0675_),
    .A2(_0678_),
    .B1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__clkbuf_4 _1273_ (.A(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_4 _1274_ (.A(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__inv_1 _1275_ (.A(_0682_),
    .Y(_1114_));
 sky130_fd_sc_hd__buf_4 _1276_ (.A(_0679_),
    .X(_0683_));
 sky130_fd_sc_hd__buf_2 _1277_ (.A(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__buf_4 _1278_ (.A(_0678_),
    .X(_0685_));
 sky130_fd_sc_hd__buf_2 _1279_ (.A(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__nand2_2 _1280_ (.A(_0684_),
    .B(_0686_),
    .Y(_1106_));
 sky130_fd_sc_hd__or3b_1 _1281_ (.A(_0676_),
    .B(_0677_),
    .C_N(_0674_),
    .X(_0687_));
 sky130_fd_sc_hd__nand3b_1 _1282_ (.A_N(_0674_),
    .B(_0677_),
    .C(_0676_),
    .Y(_0688_));
 sky130_fd_sc_hd__or4_2 _1283_ (.A(\dest_id[1][5] ),
    .B(\dest_id[1][4] ),
    .C(\dest_id[1][7] ),
    .D(\dest_id[1][6] ),
    .X(_0689_));
 sky130_fd_sc_hd__a211o_1 _1284_ (.A1(_0687_),
    .A2(_0688_),
    .B1(_0673_),
    .C1(_0689_),
    .X(_1102_));
 sky130_fd_sc_hd__clkinvlp_4 _1285_ (.A(_1102_),
    .Y(_1109_));
 sky130_fd_sc_hd__mux2i_1 _1286_ (.A0(net35),
    .A1(net172),
    .S(_1109_),
    .Y(_0690_));
 sky130_fd_sc_hd__mux2i_1 _1287_ (.A0(net103),
    .A1(net138),
    .S(_1109_),
    .Y(_0691_));
 sky130_fd_sc_hd__mux2i_1 _1288_ (.A0(_0690_),
    .A1(_0691_),
    .S(_1106_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor4_1 _1289_ (.A(_1115_),
    .B(_1104_),
    .C(_1110_),
    .D(_1112_),
    .Y(_0693_));
 sky130_fd_sc_hd__nor3_1 _1290_ (.A(net173),
    .B(_0682_),
    .C(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand3_1 _1291_ (.A(_0602_),
    .B(net69),
    .C(_0682_),
    .Y(_0695_));
 sky130_fd_sc_hd__o21ai_0 _1292_ (.A1(_0602_),
    .A2(net34),
    .B1(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__a21oi_1 _1293_ (.A1(_0692_),
    .A2(_0694_),
    .B1(_0696_),
    .Y(_0001_));
 sky130_fd_sc_hd__clkbuf_4 _1294_ (.A(\dest_id[0][2] ),
    .X(_0697_));
 sky130_fd_sc_hd__nor3b_4 _1295_ (.A(\dest_id[0][0] ),
    .B(\dest_id[0][3] ),
    .C_N(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__inv_1 _1296_ (.A(\dest_id[0][0] ),
    .Y(_0699_));
 sky130_fd_sc_hd__inv_1 _1297_ (.A(\dest_id[0][3] ),
    .Y(_0700_));
 sky130_fd_sc_hd__nor3_1 _1298_ (.A(_0699_),
    .B(_0700_),
    .C(_0697_),
    .Y(_0701_));
 sky130_fd_sc_hd__nor4_4 _1299_ (.A(\dest_id[0][5] ),
    .B(\dest_id[0][4] ),
    .C(\dest_id[0][7] ),
    .D(\dest_id[0][6] ),
    .Y(_0702_));
 sky130_fd_sc_hd__nor2b_2 _1300_ (.A(\dest_id[0][1] ),
    .B_N(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__o21a_2 _1301_ (.A1(_0698_),
    .A2(_0701_),
    .B1(_0703_),
    .X(_1091_));
 sky130_fd_sc_hd__nand2_2 _1302_ (.A(_0702_),
    .B(_0698_),
    .Y(_1094_));
 sky130_fd_sc_hd__mux2i_1 _1303_ (.A0(net35),
    .A1(net103),
    .S(_1094_),
    .Y(_0704_));
 sky130_fd_sc_hd__mux2i_1 _1304_ (.A0(net172),
    .A1(net138),
    .S(_1094_),
    .Y(_0705_));
 sky130_fd_sc_hd__mux2i_1 _1305_ (.A0(_0704_),
    .A1(_0705_),
    .S(_1091_),
    .Y(_0706_));
 sky130_fd_sc_hd__nor3b_4 _1306_ (.A(\dest_id[0][1] ),
    .B(_0697_),
    .C_N(\dest_id[0][0] ),
    .Y(_0707_));
 sky130_fd_sc_hd__o21ai_4 _1307_ (.A1(_0698_),
    .A2(_0707_),
    .B1(_0702_),
    .Y(_0708_));
 sky130_fd_sc_hd__clkbuf_2 _1308_ (.A(_1100_),
    .X(_0709_));
 sky130_fd_sc_hd__buf_4 _1309_ (.A(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__nor4_1 _1310_ (.A(_1089_),
    .B(_1092_),
    .C(_1097_),
    .D(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__nor3_1 _1311_ (.A(net237),
    .B(_0708_),
    .C(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__buf_4 _1312_ (.A(_0603_),
    .X(_0713_));
 sky130_fd_sc_hd__clkbuf_4 _1313_ (.A(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__nand3_1 _1314_ (.A(_0714_),
    .B(net69),
    .C(_0708_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21ai_0 _1315_ (.A1(_0714_),
    .A2(net102),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a21oi_1 _1316_ (.A1(_0706_),
    .A2(_0712_),
    .B1(_0716_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_1 _1317_ (.A(_1094_),
    .Y(_1087_));
 sky130_fd_sc_hd__inv_1 _1318_ (.A(_1124_),
    .Y(_1117_));
 sky130_fd_sc_hd__inv_1 _1319_ (.A(_1139_),
    .Y(_1132_));
 sky130_fd_sc_hd__inv_1 _1320_ (.A(_1091_),
    .Y(_1088_));
 sky130_fd_sc_hd__clkinv_2 _1321_ (.A(_0708_),
    .Y(_1099_));
 sky130_fd_sc_hd__inv_1 _1322_ (.A(_1106_),
    .Y(_1103_));
 sky130_fd_sc_hd__o2111ai_4 _1323_ (.A1(_0651_),
    .A2(_0653_),
    .B1(_0598_),
    .C1(_1119_),
    .D1(_0654_),
    .Y(_0717_));
 sky130_fd_sc_hd__clkbuf_4 _1324_ (.A(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_4 _1325_ (.A(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__o211ai_4 _1326_ (.A1(_0698_),
    .A2(_0707_),
    .B1(_1089_),
    .C1(_0702_),
    .Y(_0720_));
 sky130_fd_sc_hd__clkbuf_4 _1327_ (.A(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__and2_0 _1328_ (.A(_0600_),
    .B(_1104_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_2 _1329_ (.A(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__o211a_1 _1330_ (.A1(_0675_),
    .A2(_0678_),
    .B1(_0723_),
    .C1(_0679_),
    .X(_0724_));
 sky130_fd_sc_hd__buf_2 _1331_ (.A(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__clkbuf_4 _1332_ (.A(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__buf_4 _1333_ (.A(_0603_),
    .X(_0727_));
 sky130_fd_sc_hd__nand2_1 _1334_ (.A(_0727_),
    .B(\input_buffer[0][0] ),
    .Y(_0728_));
 sky130_fd_sc_hd__buf_4 _1335_ (.A(_0718_),
    .X(_0729_));
 sky130_fd_sc_hd__buf_4 _1336_ (.A(_0675_),
    .X(_0730_));
 sky130_fd_sc_hd__buf_2 _1337_ (.A(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_4 _1338_ (.A(_0723_),
    .X(_0732_));
 sky130_fd_sc_hd__o2111ai_1 _1339_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][0] ),
    .Y(_0733_));
 sky130_fd_sc_hd__o311ai_1 _1340_ (.A1(_0721_),
    .A2(_0726_),
    .A3(_0728_),
    .B1(_0729_),
    .C1(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__nor3b_4 _1341_ (.A(_0627_),
    .B(_0628_),
    .C_N(_0634_),
    .Y(_0735_));
 sky130_fd_sc_hd__o2111ai_4 _1342_ (.A1(_0735_),
    .A2(_0642_),
    .B1(_0597_),
    .C1(_1134_),
    .D1(_0633_),
    .Y(_0736_));
 sky130_fd_sc_hd__clkbuf_4 _1343_ (.A(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__o211ai_1 _1344_ (.A1(\input_buffer[2][0] ),
    .A2(_0719_),
    .B1(_0734_),
    .C1(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__o2111ai_4 _1345_ (.A1(_0607_),
    .A2(_0609_),
    .B1(_0625_),
    .C1(_1149_),
    .D1(_0610_),
    .Y(_0739_));
 sky130_fd_sc_hd__buf_4 _1346_ (.A(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__buf_4 _1347_ (.A(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__and3_1 _1348_ (.A(_0597_),
    .B(_1134_),
    .C(_1144_),
    .X(_0742_));
 sky130_fd_sc_hd__buf_4 _1349_ (.A(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__buf_6 _1350_ (.A(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(\input_buffer[3][0] ),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__nor2_1 _1352_ (.A(\input_buffer[4][0] ),
    .B(_0741_),
    .Y(_0746_));
 sky130_fd_sc_hd__a31oi_2 _1353_ (.A1(_0738_),
    .A2(_0741_),
    .A3(_0745_),
    .B1(_0746_),
    .Y(net174));
 sky130_fd_sc_hd__clkbuf_4 _1354_ (.A(_0740_),
    .X(_0747_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(_0727_),
    .B(\input_buffer[0][10] ),
    .Y(_0748_));
 sky130_fd_sc_hd__o2111ai_1 _1356_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][10] ),
    .Y(_0749_));
 sky130_fd_sc_hd__o311ai_1 _1357_ (.A1(_0721_),
    .A2(_0726_),
    .A3(_0748_),
    .B1(_0749_),
    .C1(_0729_),
    .Y(_0750_));
 sky130_fd_sc_hd__o211ai_1 _1358_ (.A1(\input_buffer[2][10] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _1359_ (.A(\input_buffer[3][10] ),
    .B(_0744_),
    .Y(_0752_));
 sky130_fd_sc_hd__nor2_1 _1360_ (.A(\input_buffer[4][10] ),
    .B(_0741_),
    .Y(_0753_));
 sky130_fd_sc_hd__a31oi_1 _1361_ (.A1(_0747_),
    .A2(_0751_),
    .A3(_0752_),
    .B1(_0753_),
    .Y(net175));
 sky130_fd_sc_hd__buf_4 _1362_ (.A(_0603_),
    .X(_0754_));
 sky130_fd_sc_hd__nand2_1 _1363_ (.A(_0754_),
    .B(\input_buffer[0][11] ),
    .Y(_0755_));
 sky130_fd_sc_hd__o2111ai_1 _1364_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][11] ),
    .Y(_0756_));
 sky130_fd_sc_hd__o311ai_2 _1365_ (.A1(_0721_),
    .A2(_0726_),
    .A3(_0755_),
    .B1(_0756_),
    .C1(_0729_),
    .Y(_0757_));
 sky130_fd_sc_hd__o211ai_1 _1366_ (.A1(\input_buffer[2][11] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand2_1 _1367_ (.A(\input_buffer[3][11] ),
    .B(_0744_),
    .Y(_0759_));
 sky130_fd_sc_hd__nor2_1 _1368_ (.A(\input_buffer[4][11] ),
    .B(_0741_),
    .Y(_0760_));
 sky130_fd_sc_hd__a31oi_1 _1369_ (.A1(_0747_),
    .A2(_0758_),
    .A3(_0759_),
    .B1(_0760_),
    .Y(net176));
 sky130_fd_sc_hd__nand2_1 _1370_ (.A(_0727_),
    .B(\input_buffer[0][12] ),
    .Y(_0761_));
 sky130_fd_sc_hd__o2111ai_1 _1371_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][12] ),
    .Y(_0762_));
 sky130_fd_sc_hd__clkbuf_4 _1372_ (.A(_0718_),
    .X(_0763_));
 sky130_fd_sc_hd__o311ai_1 _1373_ (.A1(_0721_),
    .A2(_0726_),
    .A3(_0761_),
    .B1(_0762_),
    .C1(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__o211ai_1 _1374_ (.A1(\input_buffer[2][12] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__nand2_1 _1375_ (.A(\input_buffer[3][12] ),
    .B(_0744_),
    .Y(_0766_));
 sky130_fd_sc_hd__buf_4 _1376_ (.A(_0739_),
    .X(_0767_));
 sky130_fd_sc_hd__nor2_1 _1377_ (.A(\input_buffer[4][12] ),
    .B(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__a31oi_1 _1378_ (.A1(_0747_),
    .A2(_0765_),
    .A3(_0766_),
    .B1(_0768_),
    .Y(net177));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0727_),
    .B(\input_buffer[0][13] ),
    .Y(_0769_));
 sky130_fd_sc_hd__o2111ai_1 _1380_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][13] ),
    .Y(_0770_));
 sky130_fd_sc_hd__o311ai_1 _1381_ (.A1(_0721_),
    .A2(_0726_),
    .A3(_0769_),
    .B1(_0770_),
    .C1(_0763_),
    .Y(_0771_));
 sky130_fd_sc_hd__o211ai_1 _1382_ (.A1(\input_buffer[2][13] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__nand2_1 _1383_ (.A(\input_buffer[3][13] ),
    .B(_0744_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor2_1 _1384_ (.A(\input_buffer[4][13] ),
    .B(_0767_),
    .Y(_0774_));
 sky130_fd_sc_hd__a31oi_1 _1385_ (.A1(_0747_),
    .A2(_0772_),
    .A3(_0773_),
    .B1(_0774_),
    .Y(net178));
 sky130_fd_sc_hd__clkbuf_4 _1386_ (.A(_0724_),
    .X(_0775_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(_0754_),
    .B(\input_buffer[0][14] ),
    .Y(_0776_));
 sky130_fd_sc_hd__o2111ai_1 _1388_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][14] ),
    .Y(_0777_));
 sky130_fd_sc_hd__o311ai_2 _1389_ (.A1(_0721_),
    .A2(_0775_),
    .A3(_0776_),
    .B1(_0777_),
    .C1(_0763_),
    .Y(_0778_));
 sky130_fd_sc_hd__o211ai_1 _1390_ (.A1(\input_buffer[2][14] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(\input_buffer[3][14] ),
    .B(_0744_),
    .Y(_0780_));
 sky130_fd_sc_hd__nor2_1 _1392_ (.A(\input_buffer[4][14] ),
    .B(_0767_),
    .Y(_0781_));
 sky130_fd_sc_hd__a31oi_1 _1393_ (.A1(_0747_),
    .A2(_0779_),
    .A3(_0780_),
    .B1(_0781_),
    .Y(net179));
 sky130_fd_sc_hd__nand2_1 _1394_ (.A(_0754_),
    .B(\input_buffer[0][15] ),
    .Y(_0782_));
 sky130_fd_sc_hd__o2111ai_1 _1395_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][15] ),
    .Y(_0783_));
 sky130_fd_sc_hd__o311ai_0 _1396_ (.A1(_0721_),
    .A2(_0775_),
    .A3(_0782_),
    .B1(_0783_),
    .C1(_0763_),
    .Y(_0784_));
 sky130_fd_sc_hd__o211ai_1 _1397_ (.A1(\input_buffer[2][15] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand2_1 _1398_ (.A(\input_buffer[3][15] ),
    .B(_0744_),
    .Y(_0786_));
 sky130_fd_sc_hd__nor2_1 _1399_ (.A(\input_buffer[4][15] ),
    .B(_0767_),
    .Y(_0787_));
 sky130_fd_sc_hd__a31oi_1 _1400_ (.A1(_0747_),
    .A2(_0785_),
    .A3(_0786_),
    .B1(_0787_),
    .Y(net180));
 sky130_fd_sc_hd__nand2_1 _1401_ (.A(_0754_),
    .B(\input_buffer[0][16] ),
    .Y(_0788_));
 sky130_fd_sc_hd__o2111ai_1 _1402_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][16] ),
    .Y(_0789_));
 sky130_fd_sc_hd__o311ai_0 _1403_ (.A1(_0721_),
    .A2(_0775_),
    .A3(_0788_),
    .B1(_0789_),
    .C1(_0763_),
    .Y(_0790_));
 sky130_fd_sc_hd__o211ai_1 _1404_ (.A1(\input_buffer[2][16] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _1405_ (.A(\input_buffer[3][16] ),
    .B(_0744_),
    .Y(_0792_));
 sky130_fd_sc_hd__nor2_1 _1406_ (.A(\input_buffer[4][16] ),
    .B(_0767_),
    .Y(_0793_));
 sky130_fd_sc_hd__a31oi_1 _1407_ (.A1(_0747_),
    .A2(_0791_),
    .A3(_0792_),
    .B1(_0793_),
    .Y(net181));
 sky130_fd_sc_hd__nand2_1 _1408_ (.A(_0727_),
    .B(\input_buffer[0][17] ),
    .Y(_0794_));
 sky130_fd_sc_hd__o2111ai_1 _1409_ (.A1(_0731_),
    .A2(_0686_),
    .B1(_0732_),
    .C1(_0684_),
    .D1(\input_buffer[1][17] ),
    .Y(_0795_));
 sky130_fd_sc_hd__o311ai_0 _1410_ (.A1(_0721_),
    .A2(_0775_),
    .A3(_0794_),
    .B1(_0795_),
    .C1(_0763_),
    .Y(_0796_));
 sky130_fd_sc_hd__o211ai_1 _1411_ (.A1(\input_buffer[2][17] ),
    .A2(_0719_),
    .B1(_0737_),
    .C1(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_1 _1412_ (.A(\input_buffer[3][17] ),
    .B(_0744_),
    .Y(_0798_));
 sky130_fd_sc_hd__nor2_1 _1413_ (.A(\input_buffer[4][17] ),
    .B(_0767_),
    .Y(_0799_));
 sky130_fd_sc_hd__a31oi_2 _1414_ (.A1(_0747_),
    .A2(_0797_),
    .A3(_0798_),
    .B1(_0799_),
    .Y(net182));
 sky130_fd_sc_hd__clkbuf_4 _1415_ (.A(_0718_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_4 _1416_ (.A(_0736_),
    .X(_0801_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(_0754_),
    .B(\input_buffer[0][18] ),
    .Y(_0802_));
 sky130_fd_sc_hd__buf_2 _1418_ (.A(_0730_),
    .X(_0803_));
 sky130_fd_sc_hd__buf_2 _1419_ (.A(_0685_),
    .X(_0804_));
 sky130_fd_sc_hd__buf_2 _1420_ (.A(_0683_),
    .X(_0805_));
 sky130_fd_sc_hd__o2111ai_1 _1421_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0732_),
    .C1(_0805_),
    .D1(\input_buffer[1][18] ),
    .Y(_0806_));
 sky130_fd_sc_hd__o311ai_0 _1422_ (.A1(_0721_),
    .A2(_0775_),
    .A3(_0802_),
    .B1(_0806_),
    .C1(_0763_),
    .Y(_0807_));
 sky130_fd_sc_hd__o211ai_1 _1423_ (.A1(\input_buffer[2][18] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(\input_buffer[3][18] ),
    .B(_0744_),
    .Y(_0809_));
 sky130_fd_sc_hd__nor2_1 _1425_ (.A(\input_buffer[4][18] ),
    .B(_0767_),
    .Y(_0810_));
 sky130_fd_sc_hd__a31oi_1 _1426_ (.A1(_0747_),
    .A2(_0808_),
    .A3(_0809_),
    .B1(_0810_),
    .Y(net183));
 sky130_fd_sc_hd__buf_2 _1427_ (.A(_0720_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(_0727_),
    .B(\input_buffer[0][19] ),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_4 _1429_ (.A(_0723_),
    .X(_0813_));
 sky130_fd_sc_hd__o2111ai_1 _1430_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][19] ),
    .Y(_0814_));
 sky130_fd_sc_hd__o311ai_1 _1431_ (.A1(_0811_),
    .A2(_0775_),
    .A3(_0812_),
    .B1(_0814_),
    .C1(_0763_),
    .Y(_0815_));
 sky130_fd_sc_hd__o211ai_1 _1432_ (.A1(\input_buffer[2][19] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__buf_6 _1433_ (.A(_0743_),
    .X(_0817_));
 sky130_fd_sc_hd__nand2_1 _1434_ (.A(\input_buffer[3][19] ),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _1435_ (.A(\input_buffer[4][19] ),
    .B(_0767_),
    .Y(_0819_));
 sky130_fd_sc_hd__a31oi_1 _1436_ (.A1(_0747_),
    .A2(_0816_),
    .A3(_0818_),
    .B1(_0819_),
    .Y(net184));
 sky130_fd_sc_hd__buf_4 _1437_ (.A(_0740_),
    .X(_0820_));
 sky130_fd_sc_hd__nand2_1 _1438_ (.A(_0754_),
    .B(\input_buffer[0][1] ),
    .Y(_0821_));
 sky130_fd_sc_hd__o2111ai_1 _1439_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][1] ),
    .Y(_0822_));
 sky130_fd_sc_hd__o311ai_0 _1440_ (.A1(_0811_),
    .A2(_0775_),
    .A3(_0821_),
    .B1(_0822_),
    .C1(_0763_),
    .Y(_0823_));
 sky130_fd_sc_hd__o211ai_1 _1441_ (.A1(\input_buffer[2][1] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__nand2_1 _1442_ (.A(\input_buffer[3][1] ),
    .B(_0817_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _1443_ (.A(\input_buffer[4][1] ),
    .B(_0767_),
    .Y(_0826_));
 sky130_fd_sc_hd__a31oi_1 _1444_ (.A1(_0820_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .Y(net185));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(_0754_),
    .B(\input_buffer[0][20] ),
    .Y(_0827_));
 sky130_fd_sc_hd__o2111ai_1 _1446_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][20] ),
    .Y(_0828_));
 sky130_fd_sc_hd__o311ai_0 _1447_ (.A1(_0811_),
    .A2(_0775_),
    .A3(_0827_),
    .B1(_0828_),
    .C1(_0763_),
    .Y(_0829_));
 sky130_fd_sc_hd__o211ai_1 _1448_ (.A1(\input_buffer[2][20] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_1 _1449_ (.A(\input_buffer[3][20] ),
    .B(_0817_),
    .Y(_0831_));
 sky130_fd_sc_hd__nor2_1 _1450_ (.A(\input_buffer[4][20] ),
    .B(_0767_),
    .Y(_0832_));
 sky130_fd_sc_hd__a31oi_1 _1451_ (.A1(_0820_),
    .A2(_0830_),
    .A3(_0831_),
    .B1(_0832_),
    .Y(net186));
 sky130_fd_sc_hd__nand2_1 _1452_ (.A(_0713_),
    .B(\input_buffer[0][21] ),
    .Y(_0833_));
 sky130_fd_sc_hd__o2111ai_1 _1453_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][21] ),
    .Y(_0834_));
 sky130_fd_sc_hd__buf_2 _1454_ (.A(_0717_),
    .X(_0835_));
 sky130_fd_sc_hd__o311ai_0 _1455_ (.A1(_0811_),
    .A2(_0775_),
    .A3(_0833_),
    .B1(_0834_),
    .C1(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__o211ai_1 _1456_ (.A1(\input_buffer[2][21] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(\input_buffer[3][21] ),
    .B(_0817_),
    .Y(_0838_));
 sky130_fd_sc_hd__buf_4 _1458_ (.A(_0739_),
    .X(_0839_));
 sky130_fd_sc_hd__nor2_1 _1459_ (.A(\input_buffer[4][21] ),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__a31oi_1 _1460_ (.A1(_0820_),
    .A2(_0837_),
    .A3(_0838_),
    .B1(_0840_),
    .Y(net187));
 sky130_fd_sc_hd__nand2_1 _1461_ (.A(_0754_),
    .B(\input_buffer[0][22] ),
    .Y(_0841_));
 sky130_fd_sc_hd__o2111ai_1 _1462_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][22] ),
    .Y(_0842_));
 sky130_fd_sc_hd__o311ai_0 _1463_ (.A1(_0811_),
    .A2(_0775_),
    .A3(_0841_),
    .B1(_0842_),
    .C1(_0835_),
    .Y(_0843_));
 sky130_fd_sc_hd__o211ai_1 _1464_ (.A1(\input_buffer[2][22] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _1465_ (.A(\input_buffer[3][22] ),
    .B(_0817_),
    .Y(_0845_));
 sky130_fd_sc_hd__nor2_1 _1466_ (.A(\input_buffer[4][22] ),
    .B(_0839_),
    .Y(_0846_));
 sky130_fd_sc_hd__a31oi_1 _1467_ (.A1(_0820_),
    .A2(_0844_),
    .A3(_0845_),
    .B1(_0846_),
    .Y(net188));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(_0713_),
    .B(\input_buffer[0][23] ),
    .Y(_0847_));
 sky130_fd_sc_hd__o2111ai_1 _1469_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][23] ),
    .Y(_0848_));
 sky130_fd_sc_hd__o311ai_1 _1470_ (.A1(_0811_),
    .A2(_0725_),
    .A3(_0847_),
    .B1(_0848_),
    .C1(_0835_),
    .Y(_0849_));
 sky130_fd_sc_hd__o211ai_1 _1471_ (.A1(\input_buffer[2][23] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(\input_buffer[3][23] ),
    .B(_0817_),
    .Y(_0851_));
 sky130_fd_sc_hd__nor2_1 _1473_ (.A(\input_buffer[4][23] ),
    .B(_0839_),
    .Y(_0852_));
 sky130_fd_sc_hd__a31oi_2 _1474_ (.A1(_0820_),
    .A2(_0850_),
    .A3(_0851_),
    .B1(_0852_),
    .Y(net189));
 sky130_fd_sc_hd__clkinvlp_4 _1475_ (.A(_1089_),
    .Y(_0853_));
 sky130_fd_sc_hd__buf_4 _1476_ (.A(_0603_),
    .X(_0854_));
 sky130_fd_sc_hd__nand4_4 _1477_ (.A(_0854_),
    .B(\dest_id[0][0] ),
    .C(_0702_),
    .D(_0707_),
    .Y(_0855_));
 sky130_fd_sc_hd__nor3_1 _1478_ (.A(_0853_),
    .B(_0726_),
    .C(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__clkbuf_4 _1479_ (.A(_0601_),
    .X(_0857_));
 sky130_fd_sc_hd__nand3_1 _1480_ (.A(_0857_),
    .B(_0676_),
    .C(_1104_),
    .Y(_0858_));
 sky130_fd_sc_hd__o21ai_0 _1481_ (.A1(_0682_),
    .A2(_0858_),
    .B1(_0729_),
    .Y(_0859_));
 sky130_fd_sc_hd__o21a_1 _1482_ (.A1(_0650_),
    .A2(_0718_),
    .B1(_0736_),
    .X(_0860_));
 sky130_fd_sc_hd__o21ai_0 _1483_ (.A1(_0856_),
    .A2(_0859_),
    .B1(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_1 _1484_ (.A(_0634_),
    .B(_0817_),
    .Y(_0862_));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(_0606_),
    .B(_0839_),
    .Y(_0863_));
 sky130_fd_sc_hd__a31oi_2 _1486_ (.A1(_0820_),
    .A2(_0861_),
    .A3(_0862_),
    .B1(_0863_),
    .Y(net190));
 sky130_fd_sc_hd__nand3_1 _1487_ (.A(_0857_),
    .B(_0673_),
    .C(_1104_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21ai_0 _1488_ (.A1(_0681_),
    .A2(_0864_),
    .B1(_0718_),
    .Y(_0865_));
 sky130_fd_sc_hd__nand2_1 _1489_ (.A(_0854_),
    .B(\dest_id[0][1] ),
    .Y(_0866_));
 sky130_fd_sc_hd__nor4_1 _1490_ (.A(_0853_),
    .B(_0708_),
    .C(_0726_),
    .D(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__o21a_1 _1491_ (.A1(\dest_id[2][1] ),
    .A2(_0718_),
    .B1(_0736_),
    .X(_0868_));
 sky130_fd_sc_hd__o21ai_0 _1492_ (.A1(_0865_),
    .A2(_0867_),
    .B1(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _1493_ (.A(_0627_),
    .B(_0817_),
    .Y(_0870_));
 sky130_fd_sc_hd__nor2_1 _1494_ (.A(_0604_),
    .B(_0839_),
    .Y(_0871_));
 sky130_fd_sc_hd__a31oi_2 _1495_ (.A1(_0820_),
    .A2(_0869_),
    .A3(_0870_),
    .B1(_0871_),
    .Y(net191));
 sky130_fd_sc_hd__nand3_1 _1496_ (.A(_0857_),
    .B(_0674_),
    .C(_1104_),
    .Y(_0872_));
 sky130_fd_sc_hd__o21ai_0 _1497_ (.A1(_0681_),
    .A2(_0872_),
    .B1(_0718_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _1498_ (.A(_0854_),
    .B(_0697_),
    .Y(_0874_));
 sky130_fd_sc_hd__nor4_1 _1499_ (.A(_0853_),
    .B(_0708_),
    .C(_0726_),
    .D(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__o21a_1 _1500_ (.A1(_0649_),
    .A2(_0718_),
    .B1(_0736_),
    .X(_0876_));
 sky130_fd_sc_hd__o21ai_0 _1501_ (.A1(_0873_),
    .A2(_0875_),
    .B1(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(_0628_),
    .B(_0817_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(_0605_),
    .B(_0839_),
    .Y(_0879_));
 sky130_fd_sc_hd__a31oi_2 _1504_ (.A1(_0820_),
    .A2(_0877_),
    .A3(_0878_),
    .B1(_0879_),
    .Y(net192));
 sky130_fd_sc_hd__nand2_1 _1505_ (.A(_0737_),
    .B(_0740_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _1506_ (.A(_0677_),
    .B(_0726_),
    .Y(_0881_));
 sky130_fd_sc_hd__nor4_2 _1507_ (.A(net237),
    .B(_0699_),
    .C(_0700_),
    .D(_0697_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand4b_1 _1508_ (.A_N(_0726_),
    .B(_0882_),
    .C(_1089_),
    .D(_0703_),
    .Y(_0883_));
 sky130_fd_sc_hd__nor2_1 _1509_ (.A(_0652_),
    .B(_0729_),
    .Y(_0884_));
 sky130_fd_sc_hd__a31oi_1 _1510_ (.A1(_0719_),
    .A2(_0881_),
    .A3(_0883_),
    .B1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__inv_1 _1511_ (.A(\dest_id[3][3] ),
    .Y(_0886_));
 sky130_fd_sc_hd__nor2_1 _1512_ (.A(_0608_),
    .B(_0740_),
    .Y(_0887_));
 sky130_fd_sc_hd__a31oi_1 _1513_ (.A1(_0886_),
    .A2(_0743_),
    .A3(_0740_),
    .B1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__o21a_1 _1514_ (.A1(_0880_),
    .A2(_0885_),
    .B1(_0888_),
    .X(net193));
 sky130_fd_sc_hd__nand2_1 _1515_ (.A(_0727_),
    .B(\input_buffer[0][2] ),
    .Y(_0889_));
 sky130_fd_sc_hd__o2111ai_1 _1516_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][2] ),
    .Y(_0890_));
 sky130_fd_sc_hd__o311ai_0 _1517_ (.A1(_0811_),
    .A2(_0725_),
    .A3(_0889_),
    .B1(_0890_),
    .C1(_0835_),
    .Y(_0891_));
 sky130_fd_sc_hd__o211ai_1 _1518_ (.A1(\input_buffer[2][2] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_1 _1519_ (.A(\input_buffer[3][2] ),
    .B(_0817_),
    .Y(_0893_));
 sky130_fd_sc_hd__nor2_1 _1520_ (.A(\input_buffer[4][2] ),
    .B(_0839_),
    .Y(_0894_));
 sky130_fd_sc_hd__a31oi_1 _1521_ (.A1(_0820_),
    .A2(_0892_),
    .A3(_0893_),
    .B1(_0894_),
    .Y(net194));
 sky130_fd_sc_hd__nand2_1 _1522_ (.A(_0713_),
    .B(\input_buffer[0][3] ),
    .Y(_0895_));
 sky130_fd_sc_hd__o2111ai_1 _1523_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][3] ),
    .Y(_0896_));
 sky130_fd_sc_hd__o311ai_0 _1524_ (.A1(_0811_),
    .A2(_0725_),
    .A3(_0895_),
    .B1(_0896_),
    .C1(_0835_),
    .Y(_0897_));
 sky130_fd_sc_hd__o211ai_1 _1525_ (.A1(\input_buffer[2][3] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _1526_ (.A(\input_buffer[3][3] ),
    .B(_0743_),
    .Y(_0899_));
 sky130_fd_sc_hd__nor2_1 _1527_ (.A(\input_buffer[4][3] ),
    .B(_0839_),
    .Y(_0900_));
 sky130_fd_sc_hd__a31oi_1 _1528_ (.A1(_0820_),
    .A2(_0898_),
    .A3(_0899_),
    .B1(_0900_),
    .Y(net195));
 sky130_fd_sc_hd__nand2_1 _1529_ (.A(_0727_),
    .B(\input_buffer[0][4] ),
    .Y(_0901_));
 sky130_fd_sc_hd__o2111ai_1 _1530_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0813_),
    .C1(_0805_),
    .D1(\input_buffer[1][4] ),
    .Y(_0902_));
 sky130_fd_sc_hd__o311ai_0 _1531_ (.A1(_0811_),
    .A2(_0725_),
    .A3(_0901_),
    .B1(_0902_),
    .C1(_0835_),
    .Y(_0903_));
 sky130_fd_sc_hd__o211ai_1 _1532_ (.A1(\input_buffer[2][4] ),
    .A2(_0800_),
    .B1(_0801_),
    .C1(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(\input_buffer[3][4] ),
    .B(_0743_),
    .Y(_0905_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(\input_buffer[4][4] ),
    .B(_0839_),
    .Y(_0906_));
 sky130_fd_sc_hd__a31oi_1 _1535_ (.A1(_0741_),
    .A2(_0904_),
    .A3(_0905_),
    .B1(_0906_),
    .Y(net196));
 sky130_fd_sc_hd__nand2_1 _1536_ (.A(_0727_),
    .B(\input_buffer[0][5] ),
    .Y(_0907_));
 sky130_fd_sc_hd__o2111ai_1 _1537_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0813_),
    .C1(_0683_),
    .D1(\input_buffer[1][5] ),
    .Y(_0908_));
 sky130_fd_sc_hd__o311ai_0 _1538_ (.A1(_0811_),
    .A2(_0725_),
    .A3(_0907_),
    .B1(_0908_),
    .C1(_0835_),
    .Y(_0909_));
 sky130_fd_sc_hd__o211ai_1 _1539_ (.A1(\input_buffer[2][5] ),
    .A2(_0729_),
    .B1(_0736_),
    .C1(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2_1 _1540_ (.A(\input_buffer[3][5] ),
    .B(_0743_),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_1 _1541_ (.A(\input_buffer[4][5] ),
    .B(_0839_),
    .Y(_0912_));
 sky130_fd_sc_hd__a31oi_1 _1542_ (.A1(_0741_),
    .A2(_0910_),
    .A3(_0911_),
    .B1(_0912_),
    .Y(net197));
 sky130_fd_sc_hd__nand2_1 _1543_ (.A(_0713_),
    .B(\input_buffer[0][6] ),
    .Y(_0913_));
 sky130_fd_sc_hd__o2111ai_1 _1544_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0723_),
    .C1(_0683_),
    .D1(\input_buffer[1][6] ),
    .Y(_0914_));
 sky130_fd_sc_hd__o311ai_1 _1545_ (.A1(_0720_),
    .A2(_0725_),
    .A3(_0913_),
    .B1(_0914_),
    .C1(_0835_),
    .Y(_0915_));
 sky130_fd_sc_hd__o211ai_1 _1546_ (.A1(\input_buffer[2][6] ),
    .A2(_0729_),
    .B1(_0736_),
    .C1(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(\input_buffer[3][6] ),
    .B(_0743_),
    .Y(_0917_));
 sky130_fd_sc_hd__nor2_1 _1548_ (.A(\input_buffer[4][6] ),
    .B(_0740_),
    .Y(_0918_));
 sky130_fd_sc_hd__a31oi_1 _1549_ (.A1(_0741_),
    .A2(_0916_),
    .A3(_0917_),
    .B1(_0918_),
    .Y(net198));
 sky130_fd_sc_hd__nand2_1 _1550_ (.A(_0713_),
    .B(\input_buffer[0][7] ),
    .Y(_0919_));
 sky130_fd_sc_hd__o2111ai_1 _1551_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0723_),
    .C1(_0683_),
    .D1(\input_buffer[1][7] ),
    .Y(_0920_));
 sky130_fd_sc_hd__o311ai_0 _1552_ (.A1(_0720_),
    .A2(_0725_),
    .A3(_0919_),
    .B1(_0920_),
    .C1(_0835_),
    .Y(_0921_));
 sky130_fd_sc_hd__o211ai_1 _1553_ (.A1(\input_buffer[2][7] ),
    .A2(_0729_),
    .B1(_0736_),
    .C1(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__nand2_1 _1554_ (.A(\input_buffer[3][7] ),
    .B(_0743_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_1 _1555_ (.A(\input_buffer[4][7] ),
    .B(_0740_),
    .Y(_0924_));
 sky130_fd_sc_hd__a31oi_2 _1556_ (.A1(_0741_),
    .A2(_0922_),
    .A3(_0923_),
    .B1(_0924_),
    .Y(net199));
 sky130_fd_sc_hd__nand2_1 _1557_ (.A(_0713_),
    .B(\input_buffer[0][8] ),
    .Y(_0925_));
 sky130_fd_sc_hd__o2111ai_1 _1558_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0723_),
    .C1(_0683_),
    .D1(\input_buffer[1][8] ),
    .Y(_0926_));
 sky130_fd_sc_hd__o311ai_0 _1559_ (.A1(_0720_),
    .A2(_0725_),
    .A3(_0925_),
    .B1(_0926_),
    .C1(_0835_),
    .Y(_0927_));
 sky130_fd_sc_hd__o211ai_1 _1560_ (.A1(\input_buffer[2][8] ),
    .A2(_0729_),
    .B1(_0736_),
    .C1(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _1561_ (.A(\input_buffer[3][8] ),
    .B(_0743_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _1562_ (.A(\input_buffer[4][8] ),
    .B(_0740_),
    .Y(_0930_));
 sky130_fd_sc_hd__a31oi_2 _1563_ (.A1(_0741_),
    .A2(_0928_),
    .A3(_0929_),
    .B1(_0930_),
    .Y(net200));
 sky130_fd_sc_hd__nand2_1 _1564_ (.A(_0727_),
    .B(\input_buffer[0][9] ),
    .Y(_0931_));
 sky130_fd_sc_hd__o2111ai_1 _1565_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0723_),
    .C1(_0683_),
    .D1(\input_buffer[1][9] ),
    .Y(_0932_));
 sky130_fd_sc_hd__o311ai_1 _1566_ (.A1(_0720_),
    .A2(_0725_),
    .A3(_0931_),
    .B1(_0932_),
    .C1(_0718_),
    .Y(_0933_));
 sky130_fd_sc_hd__o211ai_1 _1567_ (.A1(\input_buffer[2][9] ),
    .A2(_0729_),
    .B1(_0736_),
    .C1(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _1568_ (.A(\input_buffer[3][9] ),
    .B(_0743_),
    .Y(_0935_));
 sky130_fd_sc_hd__nor2_1 _1569_ (.A(\input_buffer[4][9] ),
    .B(_0740_),
    .Y(_0936_));
 sky130_fd_sc_hd__a31oi_2 _1570_ (.A1(_0741_),
    .A2(_0934_),
    .A3(_0935_),
    .B1(_0936_),
    .Y(net201));
 sky130_fd_sc_hd__nand2_1 _1571_ (.A(_0714_),
    .B(_1101_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand3_1 _1572_ (.A(_0599_),
    .B(_1131_),
    .C(_1119_),
    .Y(_0938_));
 sky130_fd_sc_hd__nand3_1 _1573_ (.A(_0637_),
    .B(_1146_),
    .C(_1134_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _1574_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__a31oi_1 _1575_ (.A1(_0602_),
    .A2(_1116_),
    .A3(_1104_),
    .B1(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand3_1 _1576_ (.A(_0625_),
    .B(_1161_),
    .C(_1149_),
    .Y(_0942_));
 sky130_fd_sc_hd__o211ai_2 _1577_ (.A1(_0853_),
    .A2(_0937_),
    .B1(_0941_),
    .C1(_0942_),
    .Y(net202));
 sky130_fd_sc_hd__and2_0 _1578_ (.A(_0600_),
    .B(_0680_),
    .X(_0943_));
 sky130_fd_sc_hd__buf_4 _1579_ (.A(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__a21oi_4 _1580_ (.A1(_0600_),
    .A2(_0680_),
    .B1(_1099_),
    .Y(_0945_));
 sky130_fd_sc_hd__inv_1 _1581_ (.A(_0728_),
    .Y(_0946_));
 sky130_fd_sc_hd__and2_0 _1582_ (.A(_0598_),
    .B(_0655_),
    .X(_0947_));
 sky130_fd_sc_hd__buf_2 _1583_ (.A(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__buf_6 _1584_ (.A(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__a221oi_1 _1585_ (.A1(\input_buffer[1][0] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0946_),
    .C1(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__o22ai_1 _1586_ (.A1(net203),
    .A2(_1159_),
    .B1(_1144_),
    .B2(net301),
    .Y(_0951_));
 sky130_fd_sc_hd__buf_4 _1587_ (.A(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__nand2_8 _1588_ (.A(_0598_),
    .B(_0655_),
    .Y(_0953_));
 sky130_fd_sc_hd__clkbuf_4 _1589_ (.A(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__nor2_1 _1590_ (.A(\input_buffer[2][0] ),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__nor2_1 _1591_ (.A(net203),
    .B(_1159_),
    .Y(_0956_));
 sky130_fd_sc_hd__buf_4 _1592_ (.A(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_4 _1593_ (.A(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a211oi_4 _1594_ (.A1(_0625_),
    .A2(_0611_),
    .B1(_1144_),
    .C1(net301),
    .Y(_0959_));
 sky130_fd_sc_hd__clkbuf_4 _1595_ (.A(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__a22oi_1 _1596_ (.A1(\input_buffer[4][0] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][0] ),
    .Y(_0961_));
 sky130_fd_sc_hd__o31ai_1 _1597_ (.A1(_0950_),
    .A2(_0952_),
    .A3(_0955_),
    .B1(_0961_),
    .Y(net204));
 sky130_fd_sc_hd__buf_4 _1598_ (.A(_0944_),
    .X(_0962_));
 sky130_fd_sc_hd__buf_4 _1599_ (.A(_0945_),
    .X(_0963_));
 sky130_fd_sc_hd__inv_1 _1600_ (.A(_0748_),
    .Y(_0964_));
 sky130_fd_sc_hd__buf_4 _1601_ (.A(_0948_),
    .X(_0965_));
 sky130_fd_sc_hd__a221oi_1 _1602_ (.A1(\input_buffer[1][10] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0964_),
    .C1(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__nor2_1 _1603_ (.A(\input_buffer[2][10] ),
    .B(_0954_),
    .Y(_0967_));
 sky130_fd_sc_hd__a22oi_1 _1604_ (.A1(\input_buffer[4][10] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][10] ),
    .Y(_0968_));
 sky130_fd_sc_hd__o31ai_1 _1605_ (.A1(_0952_),
    .A2(_0966_),
    .A3(_0967_),
    .B1(_0968_),
    .Y(net205));
 sky130_fd_sc_hd__and2_0 _1606_ (.A(_0713_),
    .B(\input_buffer[0][11] ),
    .X(_0969_));
 sky130_fd_sc_hd__a221oi_1 _1607_ (.A1(\input_buffer[1][11] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0969_),
    .C1(_0965_),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_1 _1608_ (.A(\input_buffer[2][11] ),
    .B(_0954_),
    .Y(_0971_));
 sky130_fd_sc_hd__a22oi_1 _1609_ (.A1(\input_buffer[4][11] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][11] ),
    .Y(_0972_));
 sky130_fd_sc_hd__o31ai_1 _1610_ (.A1(_0952_),
    .A2(_0970_),
    .A3(_0971_),
    .B1(_0972_),
    .Y(net206));
 sky130_fd_sc_hd__inv_1 _1611_ (.A(_0761_),
    .Y(_0973_));
 sky130_fd_sc_hd__a221oi_1 _1612_ (.A1(\input_buffer[1][12] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0973_),
    .C1(_0965_),
    .Y(_0974_));
 sky130_fd_sc_hd__nor2_1 _1613_ (.A(\input_buffer[2][12] ),
    .B(_0954_),
    .Y(_0975_));
 sky130_fd_sc_hd__a22oi_1 _1614_ (.A1(\input_buffer[4][12] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][12] ),
    .Y(_0976_));
 sky130_fd_sc_hd__o31ai_1 _1615_ (.A1(_0952_),
    .A2(_0974_),
    .A3(_0975_),
    .B1(_0976_),
    .Y(net207));
 sky130_fd_sc_hd__inv_1 _1616_ (.A(_0769_),
    .Y(_0977_));
 sky130_fd_sc_hd__a221oi_1 _1617_ (.A1(\input_buffer[1][13] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0977_),
    .C1(_0965_),
    .Y(_0978_));
 sky130_fd_sc_hd__nor2_1 _1618_ (.A(\input_buffer[2][13] ),
    .B(_0954_),
    .Y(_0979_));
 sky130_fd_sc_hd__a22oi_1 _1619_ (.A1(\input_buffer[4][13] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][13] ),
    .Y(_0980_));
 sky130_fd_sc_hd__o31ai_1 _1620_ (.A1(_0952_),
    .A2(_0978_),
    .A3(_0979_),
    .B1(_0980_),
    .Y(net208));
 sky130_fd_sc_hd__and2_0 _1621_ (.A(_0713_),
    .B(\input_buffer[0][14] ),
    .X(_0981_));
 sky130_fd_sc_hd__a221oi_1 _1622_ (.A1(\input_buffer[1][14] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0981_),
    .C1(_0965_),
    .Y(_0982_));
 sky130_fd_sc_hd__nor2_1 _1623_ (.A(\input_buffer[2][14] ),
    .B(_0954_),
    .Y(_0983_));
 sky130_fd_sc_hd__a22oi_1 _1624_ (.A1(\input_buffer[4][14] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][14] ),
    .Y(_0984_));
 sky130_fd_sc_hd__o31ai_1 _1625_ (.A1(_0952_),
    .A2(_0982_),
    .A3(_0983_),
    .B1(_0984_),
    .Y(net209));
 sky130_fd_sc_hd__clkbuf_4 _1626_ (.A(_0603_),
    .X(_0985_));
 sky130_fd_sc_hd__and2_0 _1627_ (.A(_0985_),
    .B(\input_buffer[0][15] ),
    .X(_0986_));
 sky130_fd_sc_hd__a221oi_1 _1628_ (.A1(\input_buffer[1][15] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0986_),
    .C1(_0965_),
    .Y(_0987_));
 sky130_fd_sc_hd__nor2_1 _1629_ (.A(\input_buffer[2][15] ),
    .B(_0954_),
    .Y(_0988_));
 sky130_fd_sc_hd__a22oi_1 _1630_ (.A1(\input_buffer[4][15] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][15] ),
    .Y(_0989_));
 sky130_fd_sc_hd__o31ai_1 _1631_ (.A1(_0952_),
    .A2(_0987_),
    .A3(_0988_),
    .B1(_0989_),
    .Y(net210));
 sky130_fd_sc_hd__and2_0 _1632_ (.A(_0985_),
    .B(\input_buffer[0][16] ),
    .X(_0990_));
 sky130_fd_sc_hd__a221oi_1 _1633_ (.A1(\input_buffer[1][16] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0990_),
    .C1(_0965_),
    .Y(_0991_));
 sky130_fd_sc_hd__nor2_1 _1634_ (.A(\input_buffer[2][16] ),
    .B(_0954_),
    .Y(_0992_));
 sky130_fd_sc_hd__a22oi_1 _1635_ (.A1(\input_buffer[4][16] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][16] ),
    .Y(_0993_));
 sky130_fd_sc_hd__o31ai_1 _1636_ (.A1(_0952_),
    .A2(_0991_),
    .A3(_0992_),
    .B1(_0993_),
    .Y(net211));
 sky130_fd_sc_hd__buf_4 _1637_ (.A(_0944_),
    .X(_0994_));
 sky130_fd_sc_hd__inv_1 _1638_ (.A(_0794_),
    .Y(_0995_));
 sky130_fd_sc_hd__a221oi_1 _1639_ (.A1(\input_buffer[1][17] ),
    .A2(_0994_),
    .B1(_0963_),
    .B2(_0995_),
    .C1(_0965_),
    .Y(_0996_));
 sky130_fd_sc_hd__nor2_1 _1640_ (.A(\input_buffer[2][17] ),
    .B(_0954_),
    .Y(_0997_));
 sky130_fd_sc_hd__a22oi_1 _1641_ (.A1(\input_buffer[4][17] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][17] ),
    .Y(_0998_));
 sky130_fd_sc_hd__o31ai_2 _1642_ (.A1(_0952_),
    .A2(_0996_),
    .A3(_0997_),
    .B1(_0998_),
    .Y(net212));
 sky130_fd_sc_hd__buf_4 _1643_ (.A(_0951_),
    .X(_0999_));
 sky130_fd_sc_hd__buf_6 _1644_ (.A(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__and2_0 _1645_ (.A(_0985_),
    .B(\input_buffer[0][18] ),
    .X(_1001_));
 sky130_fd_sc_hd__buf_4 _1646_ (.A(_0948_),
    .X(_1002_));
 sky130_fd_sc_hd__a221oi_1 _1647_ (.A1(\input_buffer[1][18] ),
    .A2(_0994_),
    .B1(_0963_),
    .B2(_1001_),
    .C1(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__nor2_1 _1648_ (.A(\input_buffer[2][18] ),
    .B(_0954_),
    .Y(_1004_));
 sky130_fd_sc_hd__a22oi_1 _1649_ (.A1(\input_buffer[4][18] ),
    .A2(_0958_),
    .B1(_0960_),
    .B2(\input_buffer[3][18] ),
    .Y(_1005_));
 sky130_fd_sc_hd__o31ai_1 _1650_ (.A1(_1000_),
    .A2(_1003_),
    .A3(_1004_),
    .B1(_1005_),
    .Y(net213));
 sky130_fd_sc_hd__clkbuf_4 _1651_ (.A(_0945_),
    .X(_1006_));
 sky130_fd_sc_hd__inv_1 _1652_ (.A(_0812_),
    .Y(_1007_));
 sky130_fd_sc_hd__a221oi_1 _1653_ (.A1(\input_buffer[1][19] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1007_),
    .C1(_1002_),
    .Y(_1008_));
 sky130_fd_sc_hd__clkbuf_4 _1654_ (.A(_0953_),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _1655_ (.A(\input_buffer[2][19] ),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__buf_4 _1656_ (.A(_0956_),
    .X(_1011_));
 sky130_fd_sc_hd__buf_4 _1657_ (.A(_0959_),
    .X(_1012_));
 sky130_fd_sc_hd__a22oi_1 _1658_ (.A1(\input_buffer[4][19] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][19] ),
    .Y(_1013_));
 sky130_fd_sc_hd__o31ai_1 _1659_ (.A1(_1000_),
    .A2(_1008_),
    .A3(_1010_),
    .B1(_1013_),
    .Y(net214));
 sky130_fd_sc_hd__and2_0 _1660_ (.A(_0985_),
    .B(\input_buffer[0][1] ),
    .X(_1014_));
 sky130_fd_sc_hd__a221oi_1 _1661_ (.A1(\input_buffer[1][1] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1014_),
    .C1(_1002_),
    .Y(_1015_));
 sky130_fd_sc_hd__nor2_1 _1662_ (.A(\input_buffer[2][1] ),
    .B(_1009_),
    .Y(_1016_));
 sky130_fd_sc_hd__a22oi_1 _1663_ (.A1(\input_buffer[4][1] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][1] ),
    .Y(_1017_));
 sky130_fd_sc_hd__o31ai_1 _1664_ (.A1(_1000_),
    .A2(_1015_),
    .A3(_1016_),
    .B1(_1017_),
    .Y(net215));
 sky130_fd_sc_hd__and2_0 _1665_ (.A(_0985_),
    .B(\input_buffer[0][20] ),
    .X(_1018_));
 sky130_fd_sc_hd__a221oi_1 _1666_ (.A1(\input_buffer[1][20] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1018_),
    .C1(_1002_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _1667_ (.A(\input_buffer[2][20] ),
    .B(_1009_),
    .Y(_1020_));
 sky130_fd_sc_hd__a22oi_1 _1668_ (.A1(\input_buffer[4][20] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][20] ),
    .Y(_1021_));
 sky130_fd_sc_hd__o31ai_1 _1669_ (.A1(_1000_),
    .A2(_1019_),
    .A3(_1020_),
    .B1(_1021_),
    .Y(net216));
 sky130_fd_sc_hd__inv_1 _1670_ (.A(_0833_),
    .Y(_1022_));
 sky130_fd_sc_hd__a221oi_1 _1671_ (.A1(\input_buffer[1][21] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1022_),
    .C1(_1002_),
    .Y(_1023_));
 sky130_fd_sc_hd__nor2_1 _1672_ (.A(\input_buffer[2][21] ),
    .B(_1009_),
    .Y(_1024_));
 sky130_fd_sc_hd__a22oi_1 _1673_ (.A1(\input_buffer[4][21] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][21] ),
    .Y(_1025_));
 sky130_fd_sc_hd__o31ai_1 _1674_ (.A1(_1000_),
    .A2(_1023_),
    .A3(_1024_),
    .B1(_1025_),
    .Y(net217));
 sky130_fd_sc_hd__and2_0 _1675_ (.A(_0985_),
    .B(\input_buffer[0][22] ),
    .X(_1026_));
 sky130_fd_sc_hd__a221oi_1 _1676_ (.A1(\input_buffer[1][22] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1026_),
    .C1(_1002_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_1 _1677_ (.A(\input_buffer[2][22] ),
    .B(_1009_),
    .Y(_1028_));
 sky130_fd_sc_hd__a22oi_1 _1678_ (.A1(\input_buffer[4][22] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][22] ),
    .Y(_1029_));
 sky130_fd_sc_hd__o31ai_1 _1679_ (.A1(_1000_),
    .A2(_1027_),
    .A3(_1028_),
    .B1(_1029_),
    .Y(net218));
 sky130_fd_sc_hd__inv_1 _1680_ (.A(_0847_),
    .Y(_1030_));
 sky130_fd_sc_hd__a221oi_1 _1681_ (.A1(\input_buffer[1][23] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1030_),
    .C1(_1002_),
    .Y(_1031_));
 sky130_fd_sc_hd__nor2_1 _1682_ (.A(\input_buffer[2][23] ),
    .B(_1009_),
    .Y(_1032_));
 sky130_fd_sc_hd__a22oi_1 _1683_ (.A1(\input_buffer[4][23] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][23] ),
    .Y(_1033_));
 sky130_fd_sc_hd__o31ai_2 _1684_ (.A1(_1000_),
    .A2(_1031_),
    .A3(_1032_),
    .B1(_1033_),
    .Y(net219));
 sky130_fd_sc_hd__a311oi_1 _1685_ (.A1(_0602_),
    .A2(_0676_),
    .A3(_0682_),
    .B1(_0957_),
    .C1(_0965_),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_1 _1686_ (.A(net301),
    .B(_1144_),
    .Y(_1035_));
 sky130_fd_sc_hd__a32oi_1 _1687_ (.A1(_0714_),
    .A2(\dest_id[0][0] ),
    .A3(_0963_),
    .B1(_1035_),
    .B2(_0634_),
    .Y(_1036_));
 sky130_fd_sc_hd__nor3_1 _1688_ (.A(_0650_),
    .B(_0953_),
    .C(_0999_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand2b_4 _1689_ (.A_N(_1144_),
    .B(_0597_),
    .Y(_1038_));
 sky130_fd_sc_hd__nor2_1 _1690_ (.A(_0608_),
    .B(_0613_),
    .Y(_1039_));
 sky130_fd_sc_hd__a211o_1 _1691_ (.A1(_0605_),
    .A2(_1039_),
    .B1(net203),
    .C1(_0606_),
    .X(_1040_));
 sky130_fd_sc_hd__o31ai_1 _1692_ (.A1(_0634_),
    .A2(_0957_),
    .A3(_1038_),
    .B1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__a211oi_1 _1693_ (.A1(_1034_),
    .A2(_1036_),
    .B1(_1037_),
    .C1(_1041_),
    .Y(net220));
 sky130_fd_sc_hd__a211oi_1 _1694_ (.A1(_0857_),
    .A2(_0681_),
    .B1(_1099_),
    .C1(_0866_),
    .Y(_1042_));
 sky130_fd_sc_hd__a211oi_1 _1695_ (.A1(_0673_),
    .A2(_0962_),
    .B1(_0949_),
    .C1(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__nor2_1 _1696_ (.A(\dest_id[2][1] ),
    .B(_1009_),
    .Y(_1044_));
 sky130_fd_sc_hd__a22oi_1 _1697_ (.A1(_0604_),
    .A2(_1011_),
    .B1(_1012_),
    .B2(_0627_),
    .Y(_1045_));
 sky130_fd_sc_hd__o31ai_2 _1698_ (.A1(_1000_),
    .A2(_1043_),
    .A3(_1044_),
    .B1(_1045_),
    .Y(net221));
 sky130_fd_sc_hd__a211oi_1 _1699_ (.A1(_0857_),
    .A2(_0681_),
    .B1(_1099_),
    .C1(_0874_),
    .Y(_1046_));
 sky130_fd_sc_hd__a211oi_1 _1700_ (.A1(_0674_),
    .A2(_0962_),
    .B1(_0949_),
    .C1(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__nor2_1 _1701_ (.A(_0649_),
    .B(_1009_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22oi_2 _1702_ (.A1(_0605_),
    .A2(_1011_),
    .B1(_1012_),
    .B2(_0628_),
    .Y(_1049_));
 sky130_fd_sc_hd__o31ai_4 _1703_ (.A1(_1000_),
    .A2(_1047_),
    .A3(_1048_),
    .B1(_1049_),
    .Y(net222));
 sky130_fd_sc_hd__and2_0 _1704_ (.A(_0985_),
    .B(\dest_id[0][3] ),
    .X(_1050_));
 sky130_fd_sc_hd__a221oi_1 _1705_ (.A1(_0677_),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1050_),
    .C1(_1002_),
    .Y(_1051_));
 sky130_fd_sc_hd__nor2_1 _1706_ (.A(_0652_),
    .B(_1009_),
    .Y(_1052_));
 sky130_fd_sc_hd__a22oi_1 _1707_ (.A1(_0608_),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\dest_id[3][3] ),
    .Y(_1053_));
 sky130_fd_sc_hd__o31ai_2 _1708_ (.A1(_1000_),
    .A2(_1051_),
    .A3(_1052_),
    .B1(_1053_),
    .Y(net223));
 sky130_fd_sc_hd__nand2_2 _1709_ (.A(_0625_),
    .B(_0611_),
    .Y(_1054_));
 sky130_fd_sc_hd__nand2_1 _1710_ (.A(_0854_),
    .B(\dest_id[0][4] ),
    .Y(_1055_));
 sky130_fd_sc_hd__a21oi_1 _1711_ (.A1(_0857_),
    .A2(_0681_),
    .B1(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__and2_0 _1712_ (.A(_0601_),
    .B(\dest_id[1][4] ),
    .X(_1057_));
 sky130_fd_sc_hd__nand3b_1 _1713_ (.A_N(\dest_id[2][4] ),
    .B(_0655_),
    .C(_0599_),
    .Y(_1058_));
 sky130_fd_sc_hd__o311ai_4 _1714_ (.A1(_0949_),
    .A2(_1056_),
    .A3(_1057_),
    .B1(_1058_),
    .C1(_1038_),
    .Y(_1059_));
 sky130_fd_sc_hd__nand2_1 _1715_ (.A(_0637_),
    .B(\dest_id[3][4] ),
    .Y(_1060_));
 sky130_fd_sc_hd__nor2_1 _1716_ (.A(\dest_id[4][4] ),
    .B(_1054_),
    .Y(_1061_));
 sky130_fd_sc_hd__a31oi_1 _1717_ (.A1(_1054_),
    .A2(_1059_),
    .A3(_1060_),
    .B1(_1061_),
    .Y(net224));
 sky130_fd_sc_hd__nand2_1 _1718_ (.A(_0854_),
    .B(\dest_id[0][5] ),
    .Y(_1062_));
 sky130_fd_sc_hd__a21oi_1 _1719_ (.A1(_0601_),
    .A2(_0681_),
    .B1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__and2_0 _1720_ (.A(_0601_),
    .B(\dest_id[1][5] ),
    .X(_1064_));
 sky130_fd_sc_hd__nand3b_1 _1721_ (.A_N(\dest_id[2][5] ),
    .B(_0655_),
    .C(_0599_),
    .Y(_1065_));
 sky130_fd_sc_hd__o311ai_4 _1722_ (.A1(_0948_),
    .A2(_1063_),
    .A3(_1064_),
    .B1(_1065_),
    .C1(_1038_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2_1 _1723_ (.A(_0637_),
    .B(\dest_id[3][5] ),
    .Y(_1067_));
 sky130_fd_sc_hd__nor2_1 _1724_ (.A(\dest_id[4][5] ),
    .B(_1054_),
    .Y(_1068_));
 sky130_fd_sc_hd__a31oi_1 _1725_ (.A1(_1054_),
    .A2(_1066_),
    .A3(_1067_),
    .B1(_1068_),
    .Y(net225));
 sky130_fd_sc_hd__and2_0 _1726_ (.A(_0985_),
    .B(\input_buffer[0][2] ),
    .X(_1069_));
 sky130_fd_sc_hd__a221oi_1 _1727_ (.A1(\input_buffer[1][2] ),
    .A2(_0994_),
    .B1(_1006_),
    .B2(_1069_),
    .C1(_1002_),
    .Y(_1070_));
 sky130_fd_sc_hd__nor2_1 _1728_ (.A(\input_buffer[2][2] ),
    .B(_1009_),
    .Y(_1071_));
 sky130_fd_sc_hd__a22oi_1 _1729_ (.A1(\input_buffer[4][2] ),
    .A2(_1011_),
    .B1(_1012_),
    .B2(\input_buffer[3][2] ),
    .Y(_1072_));
 sky130_fd_sc_hd__o31ai_1 _1730_ (.A1(_0999_),
    .A2(_1070_),
    .A3(_1071_),
    .B1(_1072_),
    .Y(net226));
 sky130_fd_sc_hd__nand2_1 _1731_ (.A(_0754_),
    .B(\dest_id[0][6] ),
    .Y(_1073_));
 sky130_fd_sc_hd__a21oi_1 _1732_ (.A1(_0601_),
    .A2(_0681_),
    .B1(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__and2_0 _1733_ (.A(_0601_),
    .B(\dest_id[1][6] ),
    .X(_1075_));
 sky130_fd_sc_hd__nand3b_1 _1734_ (.A_N(\dest_id[2][6] ),
    .B(_0655_),
    .C(_0599_),
    .Y(_1076_));
 sky130_fd_sc_hd__o311ai_2 _1735_ (.A1(_0948_),
    .A2(_1074_),
    .A3(_1075_),
    .B1(_1076_),
    .C1(_1038_),
    .Y(_1077_));
 sky130_fd_sc_hd__nand2_1 _1736_ (.A(_0637_),
    .B(\dest_id[3][6] ),
    .Y(_1078_));
 sky130_fd_sc_hd__nor2_1 _1737_ (.A(\dest_id[4][6] ),
    .B(_1054_),
    .Y(_1079_));
 sky130_fd_sc_hd__a31oi_1 _1738_ (.A1(_1054_),
    .A2(_1077_),
    .A3(_1078_),
    .B1(_1079_),
    .Y(net227));
 sky130_fd_sc_hd__nand2_1 _1739_ (.A(_0754_),
    .B(\dest_id[0][7] ),
    .Y(_1080_));
 sky130_fd_sc_hd__a21oi_1 _1740_ (.A1(_0601_),
    .A2(_0681_),
    .B1(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__and2_0 _1741_ (.A(_0601_),
    .B(\dest_id[1][7] ),
    .X(_1082_));
 sky130_fd_sc_hd__nand3b_1 _1742_ (.A_N(\dest_id[2][7] ),
    .B(_0655_),
    .C(_0599_),
    .Y(_1083_));
 sky130_fd_sc_hd__o311ai_2 _1743_ (.A1(_0948_),
    .A2(_1081_),
    .A3(_1082_),
    .B1(_1083_),
    .C1(_1038_),
    .Y(_1084_));
 sky130_fd_sc_hd__nand2_1 _1744_ (.A(_0637_),
    .B(\dest_id[3][7] ),
    .Y(_1085_));
 sky130_fd_sc_hd__nor2_1 _1745_ (.A(\dest_id[4][7] ),
    .B(_1054_),
    .Y(_1086_));
 sky130_fd_sc_hd__a31oi_1 _1746_ (.A1(_1054_),
    .A2(_1084_),
    .A3(_1085_),
    .B1(_1086_),
    .Y(net228));
 sky130_fd_sc_hd__inv_1 _1747_ (.A(_0895_),
    .Y(_0010_));
 sky130_fd_sc_hd__a221oi_1 _1748_ (.A1(\input_buffer[1][3] ),
    .A2(_0944_),
    .B1(_1006_),
    .B2(_0010_),
    .C1(_1002_),
    .Y(_0011_));
 sky130_fd_sc_hd__nor2_1 _1749_ (.A(\input_buffer[2][3] ),
    .B(_0953_),
    .Y(_0012_));
 sky130_fd_sc_hd__a22oi_1 _1750_ (.A1(\input_buffer[4][3] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][3] ),
    .Y(_0013_));
 sky130_fd_sc_hd__o31ai_1 _1751_ (.A1(_0999_),
    .A2(_0011_),
    .A3(_0012_),
    .B1(_0013_),
    .Y(net229));
 sky130_fd_sc_hd__and2_0 _1752_ (.A(_0985_),
    .B(\input_buffer[0][4] ),
    .X(_0014_));
 sky130_fd_sc_hd__a221oi_1 _1753_ (.A1(\input_buffer[1][4] ),
    .A2(_0944_),
    .B1(_1006_),
    .B2(_0014_),
    .C1(_0949_),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_1 _1754_ (.A(\input_buffer[2][4] ),
    .B(_0953_),
    .Y(_0016_));
 sky130_fd_sc_hd__a22oi_1 _1755_ (.A1(\input_buffer[4][4] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][4] ),
    .Y(_0017_));
 sky130_fd_sc_hd__o31ai_1 _1756_ (.A1(_0999_),
    .A2(_0015_),
    .A3(_0016_),
    .B1(_0017_),
    .Y(net230));
 sky130_fd_sc_hd__and2_0 _1757_ (.A(_0985_),
    .B(\input_buffer[0][5] ),
    .X(_0018_));
 sky130_fd_sc_hd__a221oi_1 _1758_ (.A1(\input_buffer[1][5] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0018_),
    .C1(_0949_),
    .Y(_0019_));
 sky130_fd_sc_hd__nor2_1 _1759_ (.A(\input_buffer[2][5] ),
    .B(_0953_),
    .Y(_0020_));
 sky130_fd_sc_hd__a22oi_1 _1760_ (.A1(\input_buffer[4][5] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][5] ),
    .Y(_0021_));
 sky130_fd_sc_hd__o31ai_1 _1761_ (.A1(_0999_),
    .A2(_0019_),
    .A3(_0020_),
    .B1(_0021_),
    .Y(net231));
 sky130_fd_sc_hd__inv_1 _1762_ (.A(_0913_),
    .Y(_0022_));
 sky130_fd_sc_hd__a221oi_1 _1763_ (.A1(\input_buffer[1][6] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0022_),
    .C1(_0949_),
    .Y(_0023_));
 sky130_fd_sc_hd__nor2_1 _1764_ (.A(\input_buffer[2][6] ),
    .B(_0953_),
    .Y(_0024_));
 sky130_fd_sc_hd__a22oi_1 _1765_ (.A1(\input_buffer[4][6] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][6] ),
    .Y(_0025_));
 sky130_fd_sc_hd__o31ai_1 _1766_ (.A1(_0999_),
    .A2(_0023_),
    .A3(_0024_),
    .B1(_0025_),
    .Y(net232));
 sky130_fd_sc_hd__inv_1 _1767_ (.A(_0919_),
    .Y(_0026_));
 sky130_fd_sc_hd__a221oi_1 _1768_ (.A1(\input_buffer[1][7] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0026_),
    .C1(_0949_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(\input_buffer[2][7] ),
    .B(_0953_),
    .Y(_0028_));
 sky130_fd_sc_hd__a22oi_1 _1770_ (.A1(\input_buffer[4][7] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][7] ),
    .Y(_0029_));
 sky130_fd_sc_hd__o31ai_1 _1771_ (.A1(_0999_),
    .A2(_0027_),
    .A3(_0028_),
    .B1(_0029_),
    .Y(net233));
 sky130_fd_sc_hd__inv_1 _1772_ (.A(_0925_),
    .Y(_0030_));
 sky130_fd_sc_hd__a221oi_1 _1773_ (.A1(\input_buffer[1][8] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0030_),
    .C1(_0949_),
    .Y(_0031_));
 sky130_fd_sc_hd__nor2_1 _1774_ (.A(\input_buffer[2][8] ),
    .B(_0953_),
    .Y(_0032_));
 sky130_fd_sc_hd__a22oi_1 _1775_ (.A1(\input_buffer[4][8] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][8] ),
    .Y(_0033_));
 sky130_fd_sc_hd__o31ai_1 _1776_ (.A1(_0999_),
    .A2(_0031_),
    .A3(_0032_),
    .B1(_0033_),
    .Y(net234));
 sky130_fd_sc_hd__and2_0 _1777_ (.A(_0603_),
    .B(\input_buffer[0][9] ),
    .X(_0034_));
 sky130_fd_sc_hd__a221oi_1 _1778_ (.A1(\input_buffer[1][9] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0034_),
    .C1(_0949_),
    .Y(_0035_));
 sky130_fd_sc_hd__nor2_1 _1779_ (.A(\input_buffer[2][9] ),
    .B(_0953_),
    .Y(_0036_));
 sky130_fd_sc_hd__a22oi_1 _1780_ (.A1(\input_buffer[4][9] ),
    .A2(_0957_),
    .B1(_0959_),
    .B2(\input_buffer[3][9] ),
    .Y(_0037_));
 sky130_fd_sc_hd__o31ai_1 _1781_ (.A1(_0999_),
    .A2(_0035_),
    .A3(_0036_),
    .B1(_0037_),
    .Y(net235));
 sky130_fd_sc_hd__nor3_1 _1782_ (.A(_0962_),
    .B(_0965_),
    .C(_0952_),
    .Y(_0038_));
 sky130_fd_sc_hd__o21ai_1 _1783_ (.A1(net237),
    .A2(_1099_),
    .B1(_0038_),
    .Y(net236));
 sky130_fd_sc_hd__nand2_8 _1784_ (.A(_0625_),
    .B(_1160_),
    .Y(_0039_));
 sky130_fd_sc_hd__clkbuf_4 _1785_ (.A(_0039_),
    .X(_0040_));
 sky130_fd_sc_hd__and2_0 _1786_ (.A(_0597_),
    .B(_1145_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_4 _1787_ (.A(_0041_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _1788_ (.A(_0042_),
    .X(_0043_));
 sky130_fd_sc_hd__nand2_8 _1789_ (.A(_0598_),
    .B(_1130_),
    .Y(_0044_));
 sky130_fd_sc_hd__clkbuf_4 _1790_ (.A(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_0 _1791_ (.A(_0600_),
    .B(_1115_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_2 _1792_ (.A(_0046_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_4 _1793_ (.A(_0047_),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_1 _1794_ (.A(\input_buffer[1][0] ),
    .B(_0048_),
    .Y(_0049_));
 sky130_fd_sc_hd__clkbuf_4 _1795_ (.A(_0713_),
    .X(_0050_));
 sky130_fd_sc_hd__buf_4 _1796_ (.A(_0709_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_2 _1797_ (.A(_0600_),
    .B(_1115_),
    .Y(_0052_));
 sky130_fd_sc_hd__buf_4 _1798_ (.A(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__nand4_1 _1799_ (.A(_0050_),
    .B(\input_buffer[0][0] ),
    .C(_0051_),
    .D(_0053_),
    .Y(_0054_));
 sky130_fd_sc_hd__buf_4 _1800_ (.A(_0044_),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_1 _1801_ (.A(\input_buffer[2][0] ),
    .B(_0055_),
    .Y(_0056_));
 sky130_fd_sc_hd__buf_4 _1802_ (.A(_0042_),
    .X(_0057_));
 sky130_fd_sc_hd__a311oi_1 _1803_ (.A1(_0045_),
    .A2(_0049_),
    .A3(_0054_),
    .B1(_0056_),
    .C1(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__a21oi_1 _1804_ (.A1(\input_buffer[3][0] ),
    .A2(_0043_),
    .B1(_0058_),
    .Y(_0059_));
 sky130_fd_sc_hd__buf_4 _1805_ (.A(_0039_),
    .X(_0060_));
 sky130_fd_sc_hd__nor2_1 _1806_ (.A(\input_buffer[4][0] ),
    .B(_0060_),
    .Y(_0061_));
 sky130_fd_sc_hd__a21oi_1 _1807_ (.A1(_0040_),
    .A2(_0059_),
    .B1(_0061_),
    .Y(net238));
 sky130_fd_sc_hd__nand2_1 _1808_ (.A(\input_buffer[1][10] ),
    .B(_0048_),
    .Y(_0062_));
 sky130_fd_sc_hd__nand4_1 _1809_ (.A(_0050_),
    .B(\input_buffer[0][10] ),
    .C(_0051_),
    .D(_0053_),
    .Y(_0063_));
 sky130_fd_sc_hd__nor2_1 _1810_ (.A(\input_buffer[2][10] ),
    .B(_0055_),
    .Y(_0064_));
 sky130_fd_sc_hd__a311oi_1 _1811_ (.A1(_0045_),
    .A2(_0062_),
    .A3(_0063_),
    .B1(_0064_),
    .C1(_0057_),
    .Y(_0065_));
 sky130_fd_sc_hd__a21oi_1 _1812_ (.A1(\input_buffer[3][10] ),
    .A2(_0043_),
    .B1(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__nor2_1 _1813_ (.A(\input_buffer[4][10] ),
    .B(_0060_),
    .Y(_0067_));
 sky130_fd_sc_hd__a21oi_1 _1814_ (.A1(_0040_),
    .A2(_0066_),
    .B1(_0067_),
    .Y(net239));
 sky130_fd_sc_hd__nand2_1 _1815_ (.A(\input_buffer[1][11] ),
    .B(_0048_),
    .Y(_0068_));
 sky130_fd_sc_hd__clkbuf_4 _1816_ (.A(_0052_),
    .X(_0069_));
 sky130_fd_sc_hd__nand3_1 _1817_ (.A(_0710_),
    .B(_0969_),
    .C(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__nor2_1 _1818_ (.A(\input_buffer[2][11] ),
    .B(_0055_),
    .Y(_0071_));
 sky130_fd_sc_hd__a311oi_1 _1819_ (.A1(_0045_),
    .A2(_0068_),
    .A3(_0070_),
    .B1(_0071_),
    .C1(_0057_),
    .Y(_0072_));
 sky130_fd_sc_hd__a21oi_1 _1820_ (.A1(\input_buffer[3][11] ),
    .A2(_0043_),
    .B1(_0072_),
    .Y(_0073_));
 sky130_fd_sc_hd__nor2_1 _1821_ (.A(\input_buffer[4][11] ),
    .B(_0060_),
    .Y(_0074_));
 sky130_fd_sc_hd__a21oi_1 _1822_ (.A1(_0040_),
    .A2(_0073_),
    .B1(_0074_),
    .Y(net240));
 sky130_fd_sc_hd__nand2_1 _1823_ (.A(\input_buffer[1][12] ),
    .B(_0048_),
    .Y(_0075_));
 sky130_fd_sc_hd__clkbuf_4 _1824_ (.A(_0709_),
    .X(_0076_));
 sky130_fd_sc_hd__nand4_1 _1825_ (.A(_0050_),
    .B(\input_buffer[0][12] ),
    .C(_0076_),
    .D(_0053_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor2_1 _1826_ (.A(\input_buffer[2][12] ),
    .B(_0055_),
    .Y(_0078_));
 sky130_fd_sc_hd__a311oi_1 _1827_ (.A1(_0045_),
    .A2(_0075_),
    .A3(_0077_),
    .B1(_0078_),
    .C1(_0057_),
    .Y(_0079_));
 sky130_fd_sc_hd__a21oi_1 _1828_ (.A1(\input_buffer[3][12] ),
    .A2(_0043_),
    .B1(_0079_),
    .Y(_0080_));
 sky130_fd_sc_hd__nor2_1 _1829_ (.A(\input_buffer[4][12] ),
    .B(_0060_),
    .Y(_0081_));
 sky130_fd_sc_hd__a21oi_1 _1830_ (.A1(_0040_),
    .A2(_0080_),
    .B1(_0081_),
    .Y(net241));
 sky130_fd_sc_hd__nand2_1 _1831_ (.A(\input_buffer[1][13] ),
    .B(_0048_),
    .Y(_0082_));
 sky130_fd_sc_hd__buf_4 _1832_ (.A(_0052_),
    .X(_0083_));
 sky130_fd_sc_hd__nand4_1 _1833_ (.A(_0050_),
    .B(\input_buffer[0][13] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__nor2_1 _1834_ (.A(\input_buffer[2][13] ),
    .B(_0055_),
    .Y(_0085_));
 sky130_fd_sc_hd__a311oi_1 _1835_ (.A1(_0045_),
    .A2(_0082_),
    .A3(_0084_),
    .B1(_0085_),
    .C1(_0057_),
    .Y(_0086_));
 sky130_fd_sc_hd__a21oi_1 _1836_ (.A1(\input_buffer[3][13] ),
    .A2(_0043_),
    .B1(_0086_),
    .Y(_0087_));
 sky130_fd_sc_hd__nor2_1 _1837_ (.A(\input_buffer[4][13] ),
    .B(_0060_),
    .Y(_0088_));
 sky130_fd_sc_hd__a21oi_1 _1838_ (.A1(_0040_),
    .A2(_0087_),
    .B1(_0088_),
    .Y(net242));
 sky130_fd_sc_hd__nand2_1 _1839_ (.A(\input_buffer[1][14] ),
    .B(_0048_),
    .Y(_0089_));
 sky130_fd_sc_hd__nand3_1 _1840_ (.A(_0710_),
    .B(_0981_),
    .C(_0069_),
    .Y(_0090_));
 sky130_fd_sc_hd__nor2_1 _1841_ (.A(\input_buffer[2][14] ),
    .B(_0055_),
    .Y(_0091_));
 sky130_fd_sc_hd__a311oi_1 _1842_ (.A1(_0045_),
    .A2(_0089_),
    .A3(_0090_),
    .B1(_0091_),
    .C1(_0057_),
    .Y(_0092_));
 sky130_fd_sc_hd__a21oi_1 _1843_ (.A1(\input_buffer[3][14] ),
    .A2(_0043_),
    .B1(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__nor2_1 _1844_ (.A(\input_buffer[4][14] ),
    .B(_0060_),
    .Y(_0094_));
 sky130_fd_sc_hd__a21oi_1 _1845_ (.A1(_0040_),
    .A2(_0093_),
    .B1(_0094_),
    .Y(net243));
 sky130_fd_sc_hd__nand2_1 _1846_ (.A(\input_buffer[1][15] ),
    .B(_0048_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand3_1 _1847_ (.A(_0710_),
    .B(_0986_),
    .C(_0069_),
    .Y(_0096_));
 sky130_fd_sc_hd__nor2_1 _1848_ (.A(\input_buffer[2][15] ),
    .B(_0055_),
    .Y(_0097_));
 sky130_fd_sc_hd__a311oi_1 _1849_ (.A1(_0045_),
    .A2(_0095_),
    .A3(_0096_),
    .B1(_0097_),
    .C1(_0057_),
    .Y(_0098_));
 sky130_fd_sc_hd__a21oi_1 _1850_ (.A1(\input_buffer[3][15] ),
    .A2(_0043_),
    .B1(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__nor2_1 _1851_ (.A(\input_buffer[4][15] ),
    .B(_0060_),
    .Y(_0100_));
 sky130_fd_sc_hd__a21oi_1 _1852_ (.A1(_0040_),
    .A2(_0099_),
    .B1(_0100_),
    .Y(net244));
 sky130_fd_sc_hd__nand2_1 _1853_ (.A(\input_buffer[1][16] ),
    .B(_0048_),
    .Y(_0101_));
 sky130_fd_sc_hd__nand3_1 _1854_ (.A(_0710_),
    .B(_0990_),
    .C(_0069_),
    .Y(_0102_));
 sky130_fd_sc_hd__nor2_1 _1855_ (.A(\input_buffer[2][16] ),
    .B(_0055_),
    .Y(_0103_));
 sky130_fd_sc_hd__a311oi_1 _1856_ (.A1(_0045_),
    .A2(_0101_),
    .A3(_0102_),
    .B1(_0103_),
    .C1(_0057_),
    .Y(_0104_));
 sky130_fd_sc_hd__a21oi_1 _1857_ (.A1(\input_buffer[3][16] ),
    .A2(_0043_),
    .B1(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__nor2_1 _1858_ (.A(\input_buffer[4][16] ),
    .B(_0060_),
    .Y(_0106_));
 sky130_fd_sc_hd__a21oi_1 _1859_ (.A1(_0040_),
    .A2(_0105_),
    .B1(_0106_),
    .Y(net245));
 sky130_fd_sc_hd__nand2_1 _1860_ (.A(\input_buffer[1][17] ),
    .B(_0048_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand4_1 _1861_ (.A(_0050_),
    .B(\input_buffer[0][17] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0108_));
 sky130_fd_sc_hd__clkbuf_4 _1862_ (.A(_0044_),
    .X(_0109_));
 sky130_fd_sc_hd__nor2_1 _1863_ (.A(\input_buffer[2][17] ),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__clkbuf_4 _1864_ (.A(_0042_),
    .X(_0111_));
 sky130_fd_sc_hd__a311oi_1 _1865_ (.A1(_0045_),
    .A2(_0107_),
    .A3(_0108_),
    .B1(_0110_),
    .C1(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__a21oi_1 _1866_ (.A1(\input_buffer[3][17] ),
    .A2(_0043_),
    .B1(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__clkbuf_4 _1867_ (.A(_0039_),
    .X(_0114_));
 sky130_fd_sc_hd__nor2_1 _1868_ (.A(\input_buffer[4][17] ),
    .B(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__a21oi_1 _1869_ (.A1(_0040_),
    .A2(_0113_),
    .B1(_0115_),
    .Y(net246));
 sky130_fd_sc_hd__nand2_1 _1870_ (.A(\input_buffer[1][18] ),
    .B(_0048_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand3_1 _1871_ (.A(_0710_),
    .B(_1001_),
    .C(_0069_),
    .Y(_0117_));
 sky130_fd_sc_hd__nor2_1 _1872_ (.A(\input_buffer[2][18] ),
    .B(_0109_),
    .Y(_0118_));
 sky130_fd_sc_hd__a311oi_1 _1873_ (.A1(_0045_),
    .A2(_0116_),
    .A3(_0117_),
    .B1(_0118_),
    .C1(_0111_),
    .Y(_0119_));
 sky130_fd_sc_hd__a21oi_1 _1874_ (.A1(\input_buffer[3][18] ),
    .A2(_0043_),
    .B1(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__nor2_1 _1875_ (.A(\input_buffer[4][18] ),
    .B(_0114_),
    .Y(_0121_));
 sky130_fd_sc_hd__a21oi_1 _1876_ (.A1(_0040_),
    .A2(_0120_),
    .B1(_0121_),
    .Y(net247));
 sky130_fd_sc_hd__clkbuf_4 _1877_ (.A(_0039_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_4 _1878_ (.A(_0042_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_4 _1879_ (.A(_0044_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _1880_ (.A(_0047_),
    .X(_0125_));
 sky130_fd_sc_hd__nand2_1 _1881_ (.A(\input_buffer[1][19] ),
    .B(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand4_1 _1882_ (.A(_0050_),
    .B(\input_buffer[0][19] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0127_));
 sky130_fd_sc_hd__nor2_1 _1883_ (.A(\input_buffer[2][19] ),
    .B(_0109_),
    .Y(_0128_));
 sky130_fd_sc_hd__a311oi_1 _1884_ (.A1(_0124_),
    .A2(_0126_),
    .A3(_0127_),
    .B1(_0128_),
    .C1(_0111_),
    .Y(_0129_));
 sky130_fd_sc_hd__a21oi_1 _1885_ (.A1(\input_buffer[3][19] ),
    .A2(_0123_),
    .B1(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__nor2_1 _1886_ (.A(\input_buffer[4][19] ),
    .B(_0114_),
    .Y(_0131_));
 sky130_fd_sc_hd__a21oi_1 _1887_ (.A1(_0122_),
    .A2(_0130_),
    .B1(_0131_),
    .Y(net248));
 sky130_fd_sc_hd__nand2_1 _1888_ (.A(\input_buffer[1][1] ),
    .B(_0125_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand3_1 _1889_ (.A(_0710_),
    .B(_1014_),
    .C(_0069_),
    .Y(_0133_));
 sky130_fd_sc_hd__nor2_1 _1890_ (.A(\input_buffer[2][1] ),
    .B(_0109_),
    .Y(_0134_));
 sky130_fd_sc_hd__a311oi_1 _1891_ (.A1(_0124_),
    .A2(_0132_),
    .A3(_0133_),
    .B1(_0134_),
    .C1(_0111_),
    .Y(_0135_));
 sky130_fd_sc_hd__a21oi_1 _1892_ (.A1(\input_buffer[3][1] ),
    .A2(_0123_),
    .B1(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__nor2_1 _1893_ (.A(\input_buffer[4][1] ),
    .B(_0114_),
    .Y(_0137_));
 sky130_fd_sc_hd__a21oi_1 _1894_ (.A1(_0122_),
    .A2(_0136_),
    .B1(_0137_),
    .Y(net249));
 sky130_fd_sc_hd__nand2_1 _1895_ (.A(\input_buffer[1][20] ),
    .B(_0125_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand3_1 _1896_ (.A(_0710_),
    .B(_1018_),
    .C(_0069_),
    .Y(_0139_));
 sky130_fd_sc_hd__nor2_1 _1897_ (.A(\input_buffer[2][20] ),
    .B(_0109_),
    .Y(_0140_));
 sky130_fd_sc_hd__a311oi_1 _1898_ (.A1(_0124_),
    .A2(_0138_),
    .A3(_0139_),
    .B1(_0140_),
    .C1(_0111_),
    .Y(_0141_));
 sky130_fd_sc_hd__a21oi_1 _1899_ (.A1(\input_buffer[3][20] ),
    .A2(_0123_),
    .B1(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__nor2_1 _1900_ (.A(\input_buffer[4][20] ),
    .B(_0114_),
    .Y(_0143_));
 sky130_fd_sc_hd__a21oi_1 _1901_ (.A1(_0122_),
    .A2(_0142_),
    .B1(_0143_),
    .Y(net250));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(\input_buffer[1][21] ),
    .B(_0125_),
    .Y(_0144_));
 sky130_fd_sc_hd__nand4_1 _1903_ (.A(_0050_),
    .B(\input_buffer[0][21] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0145_));
 sky130_fd_sc_hd__nor2_1 _1904_ (.A(\input_buffer[2][21] ),
    .B(_0109_),
    .Y(_0146_));
 sky130_fd_sc_hd__a311oi_1 _1905_ (.A1(_0124_),
    .A2(_0144_),
    .A3(_0145_),
    .B1(_0146_),
    .C1(_0111_),
    .Y(_0147_));
 sky130_fd_sc_hd__a21oi_1 _1906_ (.A1(\input_buffer[3][21] ),
    .A2(_0123_),
    .B1(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__nor2_1 _1907_ (.A(\input_buffer[4][21] ),
    .B(_0114_),
    .Y(_0149_));
 sky130_fd_sc_hd__a21oi_1 _1908_ (.A1(_0122_),
    .A2(_0148_),
    .B1(_0149_),
    .Y(net251));
 sky130_fd_sc_hd__nand2_1 _1909_ (.A(\input_buffer[1][22] ),
    .B(_0125_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand3_1 _1910_ (.A(_0710_),
    .B(_1026_),
    .C(_0069_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor2_1 _1911_ (.A(\input_buffer[2][22] ),
    .B(_0109_),
    .Y(_0152_));
 sky130_fd_sc_hd__a311oi_1 _1912_ (.A1(_0124_),
    .A2(_0150_),
    .A3(_0151_),
    .B1(_0152_),
    .C1(_0111_),
    .Y(_0153_));
 sky130_fd_sc_hd__a21oi_1 _1913_ (.A1(\input_buffer[3][22] ),
    .A2(_0123_),
    .B1(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2_1 _1914_ (.A(\input_buffer[4][22] ),
    .B(_0114_),
    .Y(_0155_));
 sky130_fd_sc_hd__a21oi_1 _1915_ (.A1(_0122_),
    .A2(_0154_),
    .B1(_0155_),
    .Y(net252));
 sky130_fd_sc_hd__nand2_1 _1916_ (.A(\input_buffer[1][23] ),
    .B(_0125_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand4_1 _1917_ (.A(_0050_),
    .B(\input_buffer[0][23] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0157_));
 sky130_fd_sc_hd__nor2_1 _1918_ (.A(\input_buffer[2][23] ),
    .B(_0109_),
    .Y(_0158_));
 sky130_fd_sc_hd__a311oi_1 _1919_ (.A1(_0124_),
    .A2(_0156_),
    .A3(_0157_),
    .B1(_0158_),
    .C1(_0111_),
    .Y(_0159_));
 sky130_fd_sc_hd__a21oi_1 _1920_ (.A1(\input_buffer[3][23] ),
    .A2(_0123_),
    .B1(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__nor2_1 _1921_ (.A(\input_buffer[4][23] ),
    .B(_0114_),
    .Y(_0161_));
 sky130_fd_sc_hd__a21oi_1 _1922_ (.A1(_0122_),
    .A2(_0160_),
    .B1(_0161_),
    .Y(net253));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(_0676_),
    .B(_0125_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand4_1 _1924_ (.A(_0050_),
    .B(\dest_id[0][0] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_1 _1925_ (.A(_0650_),
    .B(_0109_),
    .Y(_0164_));
 sky130_fd_sc_hd__a311oi_1 _1926_ (.A1(_0124_),
    .A2(_0162_),
    .A3(_0163_),
    .B1(_0164_),
    .C1(_0111_),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_1 _1927_ (.A1(_0634_),
    .A2(_0123_),
    .B1(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2_1 _1928_ (.A(_0606_),
    .B(_0114_),
    .Y(_0167_));
 sky130_fd_sc_hd__a21oi_2 _1929_ (.A1(_0122_),
    .A2(_0166_),
    .B1(_0167_),
    .Y(net254));
 sky130_fd_sc_hd__nand2_1 _1930_ (.A(_0673_),
    .B(_0125_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand4_1 _1931_ (.A(_0050_),
    .B(\dest_id[0][1] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0169_));
 sky130_fd_sc_hd__nor2_1 _1932_ (.A(\dest_id[2][1] ),
    .B(_0109_),
    .Y(_0170_));
 sky130_fd_sc_hd__a311oi_1 _1933_ (.A1(_0124_),
    .A2(_0168_),
    .A3(_0169_),
    .B1(_0170_),
    .C1(_0111_),
    .Y(_0171_));
 sky130_fd_sc_hd__a21oi_1 _1934_ (.A1(_0627_),
    .A2(_0123_),
    .B1(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__nor2_1 _1935_ (.A(_0604_),
    .B(_0114_),
    .Y(_0173_));
 sky130_fd_sc_hd__a21oi_1 _1936_ (.A1(_0122_),
    .A2(_0172_),
    .B1(_0173_),
    .Y(net255));
 sky130_fd_sc_hd__nand2_1 _1937_ (.A(_0674_),
    .B(_0125_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand4_1 _1938_ (.A(_0854_),
    .B(_0697_),
    .C(_0076_),
    .D(_0083_),
    .Y(_0175_));
 sky130_fd_sc_hd__clkbuf_4 _1939_ (.A(_0044_),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _1940_ (.A(_0649_),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__buf_4 _1941_ (.A(_0042_),
    .X(_0178_));
 sky130_fd_sc_hd__a311oi_1 _1942_ (.A1(_0124_),
    .A2(_0174_),
    .A3(_0175_),
    .B1(_0177_),
    .C1(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21oi_1 _1943_ (.A1(_0628_),
    .A2(_0123_),
    .B1(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__buf_4 _1944_ (.A(_0039_),
    .X(_0181_));
 sky130_fd_sc_hd__nor2_1 _1945_ (.A(_0605_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__a21oi_2 _1946_ (.A1(_0122_),
    .A2(_0180_),
    .B1(_0182_),
    .Y(net256));
 sky130_fd_sc_hd__nand2_1 _1947_ (.A(_0677_),
    .B(_0125_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand3_1 _1948_ (.A(_0710_),
    .B(_1050_),
    .C(_0069_),
    .Y(_0184_));
 sky130_fd_sc_hd__nor2_1 _1949_ (.A(_0652_),
    .B(_0176_),
    .Y(_0185_));
 sky130_fd_sc_hd__a311oi_1 _1950_ (.A1(_0124_),
    .A2(_0183_),
    .A3(_0184_),
    .B1(_0185_),
    .C1(_0178_),
    .Y(_0186_));
 sky130_fd_sc_hd__a21oi_1 _1951_ (.A1(\dest_id[3][3] ),
    .A2(_0123_),
    .B1(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _1952_ (.A(_0608_),
    .B(_0181_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21oi_1 _1953_ (.A1(_0122_),
    .A2(_0187_),
    .B1(_0188_),
    .Y(net257));
 sky130_fd_sc_hd__buf_4 _1954_ (.A(_0039_),
    .X(_0189_));
 sky130_fd_sc_hd__buf_4 _1955_ (.A(_0042_),
    .X(_0190_));
 sky130_fd_sc_hd__buf_4 _1956_ (.A(_0044_),
    .X(_0191_));
 sky130_fd_sc_hd__nand4_1 _1957_ (.A(_0714_),
    .B(\dest_id[0][4] ),
    .C(_0051_),
    .D(_0053_),
    .Y(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _1958_ (.A(_0047_),
    .X(_0193_));
 sky130_fd_sc_hd__nand2_1 _1959_ (.A(\dest_id[1][4] ),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _1960_ (.A(\dest_id[2][4] ),
    .B(_0176_),
    .Y(_0195_));
 sky130_fd_sc_hd__a311oi_2 _1961_ (.A1(_0191_),
    .A2(_0192_),
    .A3(_0194_),
    .B1(_0195_),
    .C1(_0178_),
    .Y(_0196_));
 sky130_fd_sc_hd__a21oi_1 _1962_ (.A1(\dest_id[3][4] ),
    .A2(_0190_),
    .B1(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _1963_ (.A(\dest_id[4][4] ),
    .B(_0181_),
    .Y(_0198_));
 sky130_fd_sc_hd__a21oi_1 _1964_ (.A1(_0189_),
    .A2(_0197_),
    .B1(_0198_),
    .Y(net258));
 sky130_fd_sc_hd__nand4_1 _1965_ (.A(_0714_),
    .B(\dest_id[0][5] ),
    .C(_0051_),
    .D(_0053_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _1966_ (.A(\dest_id[1][5] ),
    .B(_0193_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _1967_ (.A(\dest_id[2][5] ),
    .B(_0176_),
    .Y(_0201_));
 sky130_fd_sc_hd__a311oi_2 _1968_ (.A1(_0191_),
    .A2(_0199_),
    .A3(_0200_),
    .B1(_0201_),
    .C1(_0178_),
    .Y(_0202_));
 sky130_fd_sc_hd__a21oi_1 _1969_ (.A1(\dest_id[3][5] ),
    .A2(_0190_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_1 _1970_ (.A(\dest_id[4][5] ),
    .B(_0181_),
    .Y(_0204_));
 sky130_fd_sc_hd__a21oi_1 _1971_ (.A1(_0189_),
    .A2(_0203_),
    .B1(_0204_),
    .Y(net259));
 sky130_fd_sc_hd__nand2_1 _1972_ (.A(\input_buffer[1][2] ),
    .B(_0193_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand3_1 _1973_ (.A(_0051_),
    .B(_1069_),
    .C(_0069_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2_1 _1974_ (.A(\input_buffer[2][2] ),
    .B(_0176_),
    .Y(_0207_));
 sky130_fd_sc_hd__a311oi_1 _1975_ (.A1(_0191_),
    .A2(_0205_),
    .A3(_0206_),
    .B1(_0207_),
    .C1(_0178_),
    .Y(_0208_));
 sky130_fd_sc_hd__a21oi_1 _1976_ (.A1(\input_buffer[3][2] ),
    .A2(_0190_),
    .B1(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _1977_ (.A(\input_buffer[4][2] ),
    .B(_0181_),
    .Y(_0210_));
 sky130_fd_sc_hd__a21oi_1 _1978_ (.A1(_0189_),
    .A2(_0209_),
    .B1(_0210_),
    .Y(net260));
 sky130_fd_sc_hd__nand4_1 _1979_ (.A(_0714_),
    .B(\dest_id[0][6] ),
    .C(_0051_),
    .D(_0053_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _1980_ (.A(\dest_id[1][6] ),
    .B(_0047_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _1981_ (.A(\dest_id[2][6] ),
    .B(_0176_),
    .Y(_0213_));
 sky130_fd_sc_hd__a311oi_2 _1982_ (.A1(_0191_),
    .A2(_0211_),
    .A3(_0212_),
    .B1(_0213_),
    .C1(_0178_),
    .Y(_0214_));
 sky130_fd_sc_hd__a21oi_1 _1983_ (.A1(\dest_id[3][6] ),
    .A2(_0190_),
    .B1(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _1984_ (.A(\dest_id[4][6] ),
    .B(_0181_),
    .Y(_0216_));
 sky130_fd_sc_hd__a21oi_1 _1985_ (.A1(_0189_),
    .A2(_0215_),
    .B1(_0216_),
    .Y(net261));
 sky130_fd_sc_hd__nand4_1 _1986_ (.A(_0714_),
    .B(\dest_id[0][7] ),
    .C(_0051_),
    .D(_0053_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1987_ (.A(\dest_id[1][7] ),
    .B(_0047_),
    .Y(_0218_));
 sky130_fd_sc_hd__nor2_1 _1988_ (.A(\dest_id[2][7] ),
    .B(_0176_),
    .Y(_0219_));
 sky130_fd_sc_hd__a311oi_2 _1989_ (.A1(_0191_),
    .A2(_0217_),
    .A3(_0218_),
    .B1(_0219_),
    .C1(_0178_),
    .Y(_0220_));
 sky130_fd_sc_hd__a21oi_1 _1990_ (.A1(\dest_id[3][7] ),
    .A2(_0190_),
    .B1(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__nor2_1 _1991_ (.A(\dest_id[4][7] ),
    .B(_0181_),
    .Y(_0222_));
 sky130_fd_sc_hd__a21oi_1 _1992_ (.A1(_0189_),
    .A2(_0221_),
    .B1(_0222_),
    .Y(net262));
 sky130_fd_sc_hd__nand2_1 _1993_ (.A(\input_buffer[1][3] ),
    .B(_0193_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand4_1 _1994_ (.A(_0854_),
    .B(\input_buffer[0][3] ),
    .C(_0076_),
    .D(_0083_),
    .Y(_0224_));
 sky130_fd_sc_hd__nor2_1 _1995_ (.A(\input_buffer[2][3] ),
    .B(_0176_),
    .Y(_0225_));
 sky130_fd_sc_hd__a311oi_1 _1996_ (.A1(_0191_),
    .A2(_0223_),
    .A3(_0224_),
    .B1(_0225_),
    .C1(_0178_),
    .Y(_0226_));
 sky130_fd_sc_hd__a21oi_1 _1997_ (.A1(\input_buffer[3][3] ),
    .A2(_0190_),
    .B1(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_1 _1998_ (.A(\input_buffer[4][3] ),
    .B(_0181_),
    .Y(_0228_));
 sky130_fd_sc_hd__a21oi_1 _1999_ (.A1(_0189_),
    .A2(_0227_),
    .B1(_0228_),
    .Y(net263));
 sky130_fd_sc_hd__nand2_1 _2000_ (.A(\input_buffer[1][4] ),
    .B(_0193_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand3_1 _2001_ (.A(_0051_),
    .B(_0014_),
    .C(_0053_),
    .Y(_0230_));
 sky130_fd_sc_hd__nor2_1 _2002_ (.A(\input_buffer[2][4] ),
    .B(_0176_),
    .Y(_0231_));
 sky130_fd_sc_hd__a311oi_1 _2003_ (.A1(_0191_),
    .A2(_0229_),
    .A3(_0230_),
    .B1(_0231_),
    .C1(_0178_),
    .Y(_0232_));
 sky130_fd_sc_hd__a21oi_1 _2004_ (.A1(\input_buffer[3][4] ),
    .A2(_0190_),
    .B1(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _2005_ (.A(\input_buffer[4][4] ),
    .B(_0181_),
    .Y(_0234_));
 sky130_fd_sc_hd__a21oi_1 _2006_ (.A1(_0189_),
    .A2(_0233_),
    .B1(_0234_),
    .Y(net264));
 sky130_fd_sc_hd__nand2_1 _2007_ (.A(\input_buffer[1][5] ),
    .B(_0193_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand3_1 _2008_ (.A(_0051_),
    .B(_0018_),
    .C(_0053_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _2009_ (.A(\input_buffer[2][5] ),
    .B(_0176_),
    .Y(_0237_));
 sky130_fd_sc_hd__a311oi_1 _2010_ (.A1(_0191_),
    .A2(_0235_),
    .A3(_0236_),
    .B1(_0237_),
    .C1(_0178_),
    .Y(_0238_));
 sky130_fd_sc_hd__a21oi_1 _2011_ (.A1(\input_buffer[3][5] ),
    .A2(_0190_),
    .B1(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nor2_1 _2012_ (.A(\input_buffer[4][5] ),
    .B(_0181_),
    .Y(_0240_));
 sky130_fd_sc_hd__a21oi_1 _2013_ (.A1(_0189_),
    .A2(_0239_),
    .B1(_0240_),
    .Y(net265));
 sky130_fd_sc_hd__nand2_1 _2014_ (.A(\input_buffer[1][6] ),
    .B(_0193_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand4_1 _2015_ (.A(_0854_),
    .B(\input_buffer[0][6] ),
    .C(_0709_),
    .D(_0083_),
    .Y(_0242_));
 sky130_fd_sc_hd__nor2_1 _2016_ (.A(\input_buffer[2][6] ),
    .B(_0044_),
    .Y(_0243_));
 sky130_fd_sc_hd__a311oi_1 _2017_ (.A1(_0191_),
    .A2(_0241_),
    .A3(_0242_),
    .B1(_0243_),
    .C1(_0042_),
    .Y(_0244_));
 sky130_fd_sc_hd__a21oi_1 _2018_ (.A1(\input_buffer[3][6] ),
    .A2(_0190_),
    .B1(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__nor2_1 _2019_ (.A(\input_buffer[4][6] ),
    .B(_0039_),
    .Y(_0246_));
 sky130_fd_sc_hd__a21oi_1 _2020_ (.A1(_0189_),
    .A2(_0245_),
    .B1(_0246_),
    .Y(net266));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(\input_buffer[1][7] ),
    .B(_0193_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand4_1 _2022_ (.A(_0854_),
    .B(\input_buffer[0][7] ),
    .C(_0709_),
    .D(_0052_),
    .Y(_0248_));
 sky130_fd_sc_hd__nor2_1 _2023_ (.A(\input_buffer[2][7] ),
    .B(_0044_),
    .Y(_0249_));
 sky130_fd_sc_hd__a311oi_1 _2024_ (.A1(_0191_),
    .A2(_0247_),
    .A3(_0248_),
    .B1(_0249_),
    .C1(_0042_),
    .Y(_0250_));
 sky130_fd_sc_hd__a21oi_1 _2025_ (.A1(\input_buffer[3][7] ),
    .A2(_0190_),
    .B1(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__nor2_1 _2026_ (.A(\input_buffer[4][7] ),
    .B(_0039_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21oi_1 _2027_ (.A1(_0189_),
    .A2(_0251_),
    .B1(_0252_),
    .Y(net267));
 sky130_fd_sc_hd__nand2_1 _2028_ (.A(\input_buffer[1][8] ),
    .B(_0193_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand4_1 _2029_ (.A(_0854_),
    .B(\input_buffer[0][8] ),
    .C(_0709_),
    .D(_0052_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_1 _2030_ (.A(\input_buffer[2][8] ),
    .B(_0044_),
    .Y(_0255_));
 sky130_fd_sc_hd__a311oi_1 _2031_ (.A1(_0055_),
    .A2(_0253_),
    .A3(_0254_),
    .B1(_0255_),
    .C1(_0042_),
    .Y(_0256_));
 sky130_fd_sc_hd__a21oi_1 _2032_ (.A1(\input_buffer[3][8] ),
    .A2(_0057_),
    .B1(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__nor2_1 _2033_ (.A(\input_buffer[4][8] ),
    .B(_0039_),
    .Y(_0258_));
 sky130_fd_sc_hd__a21oi_1 _2034_ (.A1(_0060_),
    .A2(_0257_),
    .B1(_0258_),
    .Y(net268));
 sky130_fd_sc_hd__nand2_1 _2035_ (.A(\input_buffer[1][9] ),
    .B(_0193_),
    .Y(_0259_));
 sky130_fd_sc_hd__nand3_1 _2036_ (.A(_0051_),
    .B(_0034_),
    .C(_0053_),
    .Y(_0260_));
 sky130_fd_sc_hd__nor2_1 _2037_ (.A(\input_buffer[2][9] ),
    .B(_0044_),
    .Y(_0261_));
 sky130_fd_sc_hd__a311oi_1 _2038_ (.A1(_0055_),
    .A2(_0259_),
    .A3(_0260_),
    .B1(_0261_),
    .C1(_0042_),
    .Y(_0262_));
 sky130_fd_sc_hd__a21oi_1 _2039_ (.A1(\input_buffer[3][9] ),
    .A2(_0057_),
    .B1(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nor2_1 _2040_ (.A(\input_buffer[4][9] ),
    .B(_0039_),
    .Y(_0264_));
 sky130_fd_sc_hd__a21oi_1 _2041_ (.A1(_0060_),
    .A2(_0263_),
    .B1(_0264_),
    .Y(net269));
 sky130_fd_sc_hd__nand2_1 _2042_ (.A(_0625_),
    .B(_1150_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_1 _2043_ (.A(_1161_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3_1 _2044_ (.A(_1151_),
    .B(_0621_),
    .C(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor2_1 _2045_ (.A(_0677_),
    .B(_0689_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand4b_1 _2046_ (.A_N(_1116_),
    .B(_1105_),
    .C(_0857_),
    .D(_0676_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor3_1 _2047_ (.A(_0673_),
    .B(_0674_),
    .C(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor4b_1 _2048_ (.A(net301),
    .B(_0629_),
    .C(_1146_),
    .D_N(_1135_),
    .Y(_0271_));
 sky130_fd_sc_hd__a22oi_1 _2049_ (.A1(_0268_),
    .A2(_0270_),
    .B1(_0271_),
    .B2(_0644_),
    .Y(_0272_));
 sky130_fd_sc_hd__nor2b_1 _2050_ (.A(_1131_),
    .B_N(_1120_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand4_1 _2051_ (.A(_0599_),
    .B(_0651_),
    .C(_0667_),
    .D(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor4b_1 _2052_ (.A(\dest_id[0][3] ),
    .B(_0697_),
    .C(_1101_),
    .D_N(_1090_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand4_1 _2053_ (.A(_0714_),
    .B(\dest_id[0][0] ),
    .C(_0703_),
    .D(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand4_1 _2054_ (.A(_0267_),
    .B(_0272_),
    .C(_0274_),
    .D(_0276_),
    .Y(net270));
 sky130_fd_sc_hd__o2111a_1 _2055_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0600_),
    .C1(_1112_),
    .D1(_0683_),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_4 _2056_ (.A(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _2057_ (.A(_0598_),
    .B(_1127_),
    .Y(_0279_));
 sky130_fd_sc_hd__nor2_4 _2058_ (.A(_0655_),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__clkbuf_4 _2059_ (.A(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__o211ai_4 _2060_ (.A1(_0698_),
    .A2(_0707_),
    .B1(_1097_),
    .C1(_0702_),
    .Y(_0282_));
 sky130_fd_sc_hd__clkbuf_4 _2061_ (.A(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__buf_4 _2062_ (.A(_0277_),
    .X(_0284_));
 sky130_fd_sc_hd__nor3_1 _2063_ (.A(_0728_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__a211oi_1 _2064_ (.A1(\input_buffer[1][0] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__a211o_2 _2065_ (.A1(_0669_),
    .A2(_0658_),
    .B1(_0279_),
    .C1(_0656_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_4 _2066_ (.A(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__o2111ai_4 _2067_ (.A1(_0735_),
    .A2(_0642_),
    .B1(_0597_),
    .C1(_1142_),
    .D1(_0633_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _2068_ (.A(\input_buffer_valid[4] ),
    .B(_1157_),
    .Y(_0290_));
 sky130_fd_sc_hd__a211o_1 _2069_ (.A1(_0619_),
    .A2(_0615_),
    .B1(_0290_),
    .C1(_0613_),
    .X(_0291_));
 sky130_fd_sc_hd__and2_2 _2070_ (.A(_0289_),
    .B(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_4 _2071_ (.A(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__o21ai_0 _2072_ (.A1(\input_buffer[2][0] ),
    .A2(_0288_),
    .B1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__a211oi_4 _2073_ (.A1(_0619_),
    .A2(_0615_),
    .B1(_0290_),
    .C1(_0613_),
    .Y(_0295_));
 sky130_fd_sc_hd__buf_4 _2074_ (.A(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_8 _2075_ (.A(_0289_),
    .B(_0295_),
    .Y(_0297_));
 sky130_fd_sc_hd__buf_6 _2076_ (.A(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__a22oi_1 _2077_ (.A1(\input_buffer[4][0] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][0] ),
    .Y(_0299_));
 sky130_fd_sc_hd__o21ai_0 _2078_ (.A1(_0286_),
    .A2(_0294_),
    .B1(_0299_),
    .Y(net272));
 sky130_fd_sc_hd__nor3_1 _2079_ (.A(_0748_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0300_));
 sky130_fd_sc_hd__a211oi_1 _2080_ (.A1(\input_buffer[1][10] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__o21ai_0 _2081_ (.A1(\input_buffer[2][10] ),
    .A2(_0288_),
    .B1(_0293_),
    .Y(_0302_));
 sky130_fd_sc_hd__a22oi_1 _2082_ (.A1(\input_buffer[4][10] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][10] ),
    .Y(_0303_));
 sky130_fd_sc_hd__o21ai_0 _2083_ (.A1(_0301_),
    .A2(_0302_),
    .B1(_0303_),
    .Y(net273));
 sky130_fd_sc_hd__nor3_1 _2084_ (.A(_0755_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0304_));
 sky130_fd_sc_hd__a211oi_1 _2085_ (.A1(\input_buffer[1][11] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21ai_0 _2086_ (.A1(\input_buffer[2][11] ),
    .A2(_0288_),
    .B1(_0293_),
    .Y(_0306_));
 sky130_fd_sc_hd__a22oi_1 _2087_ (.A1(\input_buffer[4][11] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][11] ),
    .Y(_0307_));
 sky130_fd_sc_hd__o21ai_0 _2088_ (.A1(_0305_),
    .A2(_0306_),
    .B1(_0307_),
    .Y(net274));
 sky130_fd_sc_hd__nor3_1 _2089_ (.A(_0761_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0308_));
 sky130_fd_sc_hd__a211oi_1 _2090_ (.A1(\input_buffer[1][12] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__o21ai_0 _2091_ (.A1(\input_buffer[2][12] ),
    .A2(_0288_),
    .B1(_0293_),
    .Y(_0310_));
 sky130_fd_sc_hd__a22oi_1 _2092_ (.A1(\input_buffer[4][12] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][12] ),
    .Y(_0311_));
 sky130_fd_sc_hd__o21ai_0 _2093_ (.A1(_0309_),
    .A2(_0310_),
    .B1(_0311_),
    .Y(net275));
 sky130_fd_sc_hd__nor3_1 _2094_ (.A(_0769_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0312_));
 sky130_fd_sc_hd__a211oi_1 _2095_ (.A1(\input_buffer[1][13] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__o21ai_0 _2096_ (.A1(\input_buffer[2][13] ),
    .A2(_0288_),
    .B1(_0293_),
    .Y(_0314_));
 sky130_fd_sc_hd__a22oi_1 _2097_ (.A1(\input_buffer[4][13] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][13] ),
    .Y(_0315_));
 sky130_fd_sc_hd__o21ai_0 _2098_ (.A1(_0313_),
    .A2(_0314_),
    .B1(_0315_),
    .Y(net276));
 sky130_fd_sc_hd__clkbuf_4 _2099_ (.A(_0277_),
    .X(_0316_));
 sky130_fd_sc_hd__nor3_1 _2100_ (.A(_0776_),
    .B(_0283_),
    .C(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__a211oi_1 _2101_ (.A1(\input_buffer[1][14] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__o21ai_0 _2102_ (.A1(\input_buffer[2][14] ),
    .A2(_0288_),
    .B1(_0293_),
    .Y(_0319_));
 sky130_fd_sc_hd__a22oi_1 _2103_ (.A1(\input_buffer[4][14] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][14] ),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_0 _2104_ (.A1(_0318_),
    .A2(_0319_),
    .B1(_0320_),
    .Y(net277));
 sky130_fd_sc_hd__nor3_1 _2105_ (.A(_0782_),
    .B(_0283_),
    .C(_0316_),
    .Y(_0321_));
 sky130_fd_sc_hd__a211oi_1 _2106_ (.A1(\input_buffer[1][15] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__clkbuf_4 _2107_ (.A(_0287_),
    .X(_0323_));
 sky130_fd_sc_hd__o21ai_0 _2108_ (.A1(\input_buffer[2][15] ),
    .A2(_0323_),
    .B1(_0293_),
    .Y(_0324_));
 sky130_fd_sc_hd__buf_6 _2109_ (.A(_0297_),
    .X(_0325_));
 sky130_fd_sc_hd__a22oi_1 _2110_ (.A1(\input_buffer[4][15] ),
    .A2(_0296_),
    .B1(_0325_),
    .B2(\input_buffer[3][15] ),
    .Y(_0326_));
 sky130_fd_sc_hd__o21ai_1 _2111_ (.A1(_0322_),
    .A2(_0324_),
    .B1(_0326_),
    .Y(net278));
 sky130_fd_sc_hd__nor3_1 _2112_ (.A(_0788_),
    .B(_0283_),
    .C(_0316_),
    .Y(_0327_));
 sky130_fd_sc_hd__a211oi_1 _2113_ (.A1(\input_buffer[1][16] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__o21ai_0 _2114_ (.A1(\input_buffer[2][16] ),
    .A2(_0323_),
    .B1(_0293_),
    .Y(_0329_));
 sky130_fd_sc_hd__clkbuf_4 _2115_ (.A(_0295_),
    .X(_0330_));
 sky130_fd_sc_hd__a22oi_1 _2116_ (.A1(\input_buffer[4][16] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][16] ),
    .Y(_0331_));
 sky130_fd_sc_hd__o21ai_1 _2117_ (.A1(_0328_),
    .A2(_0329_),
    .B1(_0331_),
    .Y(net279));
 sky130_fd_sc_hd__nand2_2 _2118_ (.A(_0289_),
    .B(_0291_),
    .Y(_0332_));
 sky130_fd_sc_hd__clkbuf_4 _2119_ (.A(_0277_),
    .X(_0333_));
 sky130_fd_sc_hd__nor3_1 _2120_ (.A(_0794_),
    .B(_0282_),
    .C(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__a211oi_1 _2121_ (.A1(\input_buffer[1][17] ),
    .A2(_0284_),
    .B1(_0280_),
    .C1(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_1 _2122_ (.A(\input_buffer[2][17] ),
    .B(_0288_),
    .Y(_0336_));
 sky130_fd_sc_hd__a22oi_1 _2123_ (.A1(\input_buffer[4][17] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][17] ),
    .Y(_0337_));
 sky130_fd_sc_hd__o31ai_2 _2124_ (.A1(_0332_),
    .A2(_0335_),
    .A3(_0336_),
    .B1(_0337_),
    .Y(net280));
 sky130_fd_sc_hd__nor3_1 _2125_ (.A(_0802_),
    .B(_0283_),
    .C(_0316_),
    .Y(_0338_));
 sky130_fd_sc_hd__a211oi_1 _2126_ (.A1(\input_buffer[1][18] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__o21ai_0 _2127_ (.A1(\input_buffer[2][18] ),
    .A2(_0323_),
    .B1(_0293_),
    .Y(_0340_));
 sky130_fd_sc_hd__a22oi_1 _2128_ (.A1(\input_buffer[4][18] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][18] ),
    .Y(_0341_));
 sky130_fd_sc_hd__o21ai_1 _2129_ (.A1(_0339_),
    .A2(_0340_),
    .B1(_0341_),
    .Y(net281));
 sky130_fd_sc_hd__nor3_1 _2130_ (.A(_0812_),
    .B(_0283_),
    .C(_0316_),
    .Y(_0342_));
 sky130_fd_sc_hd__a211oi_1 _2131_ (.A1(\input_buffer[1][19] ),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__clkbuf_4 _2132_ (.A(_0292_),
    .X(_0344_));
 sky130_fd_sc_hd__o21ai_0 _2133_ (.A1(\input_buffer[2][19] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__a22oi_1 _2134_ (.A1(\input_buffer[4][19] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][19] ),
    .Y(_0346_));
 sky130_fd_sc_hd__o21ai_1 _2135_ (.A1(_0343_),
    .A2(_0345_),
    .B1(_0346_),
    .Y(net282));
 sky130_fd_sc_hd__clkbuf_4 _2136_ (.A(_0277_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_4 _2137_ (.A(_0280_),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_4 _2138_ (.A(_0282_),
    .X(_0349_));
 sky130_fd_sc_hd__nor3_1 _2139_ (.A(_0821_),
    .B(_0349_),
    .C(_0316_),
    .Y(_0350_));
 sky130_fd_sc_hd__a211oi_1 _2140_ (.A1(\input_buffer[1][1] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__o21ai_0 _2141_ (.A1(\input_buffer[2][1] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0352_));
 sky130_fd_sc_hd__a22oi_1 _2142_ (.A1(\input_buffer[4][1] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][1] ),
    .Y(_0353_));
 sky130_fd_sc_hd__o21ai_1 _2143_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0353_),
    .Y(net283));
 sky130_fd_sc_hd__nor3_1 _2144_ (.A(_0827_),
    .B(_0349_),
    .C(_0316_),
    .Y(_0354_));
 sky130_fd_sc_hd__a211oi_1 _2145_ (.A1(\input_buffer[1][20] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__o21ai_0 _2146_ (.A1(\input_buffer[2][20] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0356_));
 sky130_fd_sc_hd__a22oi_1 _2147_ (.A1(\input_buffer[4][20] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][20] ),
    .Y(_0357_));
 sky130_fd_sc_hd__o21ai_0 _2148_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0357_),
    .Y(net284));
 sky130_fd_sc_hd__nor3_1 _2149_ (.A(_0833_),
    .B(_0349_),
    .C(_0316_),
    .Y(_0358_));
 sky130_fd_sc_hd__a211oi_1 _2150_ (.A1(\input_buffer[1][21] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__o21ai_0 _2151_ (.A1(\input_buffer[2][21] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0360_));
 sky130_fd_sc_hd__a22oi_1 _2152_ (.A1(\input_buffer[4][21] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][21] ),
    .Y(_0361_));
 sky130_fd_sc_hd__o21ai_0 _2153_ (.A1(_0359_),
    .A2(_0360_),
    .B1(_0361_),
    .Y(net285));
 sky130_fd_sc_hd__nor3_1 _2154_ (.A(_0841_),
    .B(_0349_),
    .C(_0316_),
    .Y(_0362_));
 sky130_fd_sc_hd__a211oi_1 _2155_ (.A1(\input_buffer[1][22] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__o21ai_0 _2156_ (.A1(\input_buffer[2][22] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0364_));
 sky130_fd_sc_hd__a22oi_1 _2157_ (.A1(\input_buffer[4][22] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][22] ),
    .Y(_0365_));
 sky130_fd_sc_hd__o21ai_0 _2158_ (.A1(_0363_),
    .A2(_0364_),
    .B1(_0365_),
    .Y(net286));
 sky130_fd_sc_hd__nor3_1 _2159_ (.A(_0847_),
    .B(_0282_),
    .C(_0333_),
    .Y(_0366_));
 sky130_fd_sc_hd__a211oi_1 _2160_ (.A1(\input_buffer[1][23] ),
    .A2(_0284_),
    .B1(_0280_),
    .C1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__nor2_1 _2161_ (.A(\input_buffer[2][23] ),
    .B(_0288_),
    .Y(_0368_));
 sky130_fd_sc_hd__a22oi_1 _2162_ (.A1(\input_buffer[4][23] ),
    .A2(_0296_),
    .B1(_0298_),
    .B2(\input_buffer[3][23] ),
    .Y(_0369_));
 sky130_fd_sc_hd__o31ai_2 _2163_ (.A1(_0332_),
    .A2(_0367_),
    .A3(_0368_),
    .B1(_0369_),
    .Y(net287));
 sky130_fd_sc_hd__nor3b_1 _2164_ (.A(_0284_),
    .B(_0855_),
    .C_N(_1097_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand3_1 _2165_ (.A(_0602_),
    .B(_0676_),
    .C(_1112_),
    .Y(_0371_));
 sky130_fd_sc_hd__clkbuf_4 _2166_ (.A(_0287_),
    .X(_0372_));
 sky130_fd_sc_hd__o21ai_0 _2167_ (.A1(_0682_),
    .A2(_0371_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__o221ai_2 _2168_ (.A1(_0650_),
    .A2(_0288_),
    .B1(_0370_),
    .B2(_0373_),
    .C1(_0293_),
    .Y(_0374_));
 sky130_fd_sc_hd__a22oi_1 _2169_ (.A1(_0606_),
    .A2(_0296_),
    .B1(_0298_),
    .B2(_0634_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _2170_ (.A(_0374_),
    .B(_0375_),
    .Y(net288));
 sky130_fd_sc_hd__nor2_1 _2171_ (.A(_0708_),
    .B(_0866_),
    .Y(_0376_));
 sky130_fd_sc_hd__o2111ai_4 _2172_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0601_),
    .C1(_1112_),
    .D1(_0683_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand3_1 _2173_ (.A(_0602_),
    .B(_0673_),
    .C(_1112_),
    .Y(_0378_));
 sky130_fd_sc_hd__o21ai_0 _2174_ (.A1(_0682_),
    .A2(_0378_),
    .B1(_0372_),
    .Y(_0379_));
 sky130_fd_sc_hd__a31oi_1 _2175_ (.A1(_1097_),
    .A2(_0376_),
    .A3(_0377_),
    .B1(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__o21ai_0 _2176_ (.A1(\dest_id[2][1] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0381_));
 sky130_fd_sc_hd__a22oi_1 _2177_ (.A1(_0604_),
    .A2(_0330_),
    .B1(_0325_),
    .B2(_0627_),
    .Y(_0382_));
 sky130_fd_sc_hd__o21ai_2 _2178_ (.A1(_0380_),
    .A2(_0381_),
    .B1(_0382_),
    .Y(net289));
 sky130_fd_sc_hd__nor2_1 _2179_ (.A(_0708_),
    .B(_0874_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_1 _2180_ (.A(_0857_),
    .B(_0674_),
    .C(_1112_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21ai_0 _2181_ (.A1(_0681_),
    .A2(_0384_),
    .B1(_0287_),
    .Y(_0385_));
 sky130_fd_sc_hd__a31oi_1 _2182_ (.A1(_1097_),
    .A2(_0383_),
    .A3(_0377_),
    .B1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__nor2_1 _2183_ (.A(_0649_),
    .B(_0288_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _2184_ (.A(_0606_),
    .B(_0291_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_1 _2185_ (.A1(_0628_),
    .A2(_0298_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__o31ai_2 _2186_ (.A1(_0332_),
    .A2(_0386_),
    .A3(_0387_),
    .B1(_0389_),
    .Y(net290));
 sky130_fd_sc_hd__nand2_1 _2187_ (.A(_0677_),
    .B(_0333_),
    .Y(_0390_));
 sky130_fd_sc_hd__nand4_1 _2188_ (.A(_1097_),
    .B(_0703_),
    .C(_0882_),
    .D(_0377_),
    .Y(_0391_));
 sky130_fd_sc_hd__nor2_1 _2189_ (.A(_0652_),
    .B(_0287_),
    .Y(_0392_));
 sky130_fd_sc_hd__a31oi_1 _2190_ (.A1(_0372_),
    .A2(_0390_),
    .A3(_0391_),
    .B1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_1 _2191_ (.A(_0886_),
    .B(_0297_),
    .Y(_0394_));
 sky130_fd_sc_hd__o221a_1 _2192_ (.A1(_0608_),
    .A2(_0291_),
    .B1(_0332_),
    .B2(_0393_),
    .C1(_0394_),
    .X(net291));
 sky130_fd_sc_hd__nor3_1 _2193_ (.A(_0889_),
    .B(_0349_),
    .C(_0316_),
    .Y(_0395_));
 sky130_fd_sc_hd__a211oi_1 _2194_ (.A1(\input_buffer[1][2] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__o21ai_0 _2195_ (.A1(\input_buffer[2][2] ),
    .A2(_0323_),
    .B1(_0344_),
    .Y(_0397_));
 sky130_fd_sc_hd__a22oi_1 _2196_ (.A1(\input_buffer[4][2] ),
    .A2(_0330_),
    .B1(_0325_),
    .B2(\input_buffer[3][2] ),
    .Y(_0398_));
 sky130_fd_sc_hd__o21ai_0 _2197_ (.A1(_0396_),
    .A2(_0397_),
    .B1(_0398_),
    .Y(net292));
 sky130_fd_sc_hd__nor3_1 _2198_ (.A(_0895_),
    .B(_0349_),
    .C(_0333_),
    .Y(_0399_));
 sky130_fd_sc_hd__a211oi_1 _2199_ (.A1(\input_buffer[1][3] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o21ai_0 _2200_ (.A1(\input_buffer[2][3] ),
    .A2(_0372_),
    .B1(_0344_),
    .Y(_0401_));
 sky130_fd_sc_hd__a22oi_1 _2201_ (.A1(\input_buffer[4][3] ),
    .A2(_0330_),
    .B1(_0297_),
    .B2(\input_buffer[3][3] ),
    .Y(_0402_));
 sky130_fd_sc_hd__o21ai_0 _2202_ (.A1(_0400_),
    .A2(_0401_),
    .B1(_0402_),
    .Y(net293));
 sky130_fd_sc_hd__nor3_1 _2203_ (.A(_0901_),
    .B(_0349_),
    .C(_0333_),
    .Y(_0403_));
 sky130_fd_sc_hd__a211oi_1 _2204_ (.A1(\input_buffer[1][4] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__o21ai_0 _2205_ (.A1(\input_buffer[2][4] ),
    .A2(_0372_),
    .B1(_0344_),
    .Y(_0405_));
 sky130_fd_sc_hd__a22oi_1 _2206_ (.A1(\input_buffer[4][4] ),
    .A2(_0295_),
    .B1(_0297_),
    .B2(\input_buffer[3][4] ),
    .Y(_0406_));
 sky130_fd_sc_hd__o21ai_0 _2207_ (.A1(_0404_),
    .A2(_0405_),
    .B1(_0406_),
    .Y(net294));
 sky130_fd_sc_hd__nor3_1 _2208_ (.A(_0907_),
    .B(_0349_),
    .C(_0333_),
    .Y(_0407_));
 sky130_fd_sc_hd__a211oi_1 _2209_ (.A1(\input_buffer[1][5] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__o21ai_0 _2210_ (.A1(\input_buffer[2][5] ),
    .A2(_0372_),
    .B1(_0344_),
    .Y(_0409_));
 sky130_fd_sc_hd__a22oi_1 _2211_ (.A1(\input_buffer[4][5] ),
    .A2(_0295_),
    .B1(_0297_),
    .B2(\input_buffer[3][5] ),
    .Y(_0410_));
 sky130_fd_sc_hd__o21ai_0 _2212_ (.A1(_0408_),
    .A2(_0409_),
    .B1(_0410_),
    .Y(net295));
 sky130_fd_sc_hd__nor3_1 _2213_ (.A(_0913_),
    .B(_0349_),
    .C(_0333_),
    .Y(_0411_));
 sky130_fd_sc_hd__a211oi_1 _2214_ (.A1(\input_buffer[1][6] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__o21ai_0 _2215_ (.A1(\input_buffer[2][6] ),
    .A2(_0372_),
    .B1(_0292_),
    .Y(_0413_));
 sky130_fd_sc_hd__a22oi_1 _2216_ (.A1(\input_buffer[4][6] ),
    .A2(_0295_),
    .B1(_0297_),
    .B2(\input_buffer[3][6] ),
    .Y(_0414_));
 sky130_fd_sc_hd__o21ai_0 _2217_ (.A1(_0412_),
    .A2(_0413_),
    .B1(_0414_),
    .Y(net296));
 sky130_fd_sc_hd__nor3_1 _2218_ (.A(_0919_),
    .B(_0349_),
    .C(_0333_),
    .Y(_0415_));
 sky130_fd_sc_hd__a211oi_1 _2219_ (.A1(\input_buffer[1][7] ),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__o21ai_0 _2220_ (.A1(\input_buffer[2][7] ),
    .A2(_0372_),
    .B1(_0292_),
    .Y(_0417_));
 sky130_fd_sc_hd__a22oi_1 _2221_ (.A1(\input_buffer[4][7] ),
    .A2(_0295_),
    .B1(_0297_),
    .B2(\input_buffer[3][7] ),
    .Y(_0418_));
 sky130_fd_sc_hd__o21ai_1 _2222_ (.A1(_0416_),
    .A2(_0417_),
    .B1(_0418_),
    .Y(net297));
 sky130_fd_sc_hd__nor3_1 _2223_ (.A(_0925_),
    .B(_0282_),
    .C(_0333_),
    .Y(_0419_));
 sky130_fd_sc_hd__a211oi_1 _2224_ (.A1(\input_buffer[1][8] ),
    .A2(_0284_),
    .B1(_0280_),
    .C1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__o21ai_0 _2225_ (.A1(\input_buffer[2][8] ),
    .A2(_0372_),
    .B1(_0292_),
    .Y(_0421_));
 sky130_fd_sc_hd__a22oi_1 _2226_ (.A1(\input_buffer[4][8] ),
    .A2(_0295_),
    .B1(_0297_),
    .B2(\input_buffer[3][8] ),
    .Y(_0422_));
 sky130_fd_sc_hd__o21ai_1 _2227_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0422_),
    .Y(net298));
 sky130_fd_sc_hd__nor3_1 _2228_ (.A(_0931_),
    .B(_0282_),
    .C(_0333_),
    .Y(_0423_));
 sky130_fd_sc_hd__a211oi_1 _2229_ (.A1(\input_buffer[1][9] ),
    .A2(_0284_),
    .B1(_0280_),
    .C1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21ai_0 _2230_ (.A1(\input_buffer[2][9] ),
    .A2(_0372_),
    .B1(_0292_),
    .Y(_0425_));
 sky130_fd_sc_hd__a22oi_1 _2231_ (.A1(\input_buffer[4][9] ),
    .A2(_0295_),
    .B1(_0297_),
    .B2(\input_buffer[3][9] ),
    .Y(_0426_));
 sky130_fd_sc_hd__o21ai_1 _2232_ (.A1(_0424_),
    .A2(_0425_),
    .B1(_0426_),
    .Y(net299));
 sky130_fd_sc_hd__nand2_1 _2233_ (.A(_0625_),
    .B(_1161_),
    .Y(_0427_));
 sky130_fd_sc_hd__nand2_1 _2234_ (.A(_0629_),
    .B(_0645_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand2_1 _2235_ (.A(_0637_),
    .B(_1146_),
    .Y(_0429_));
 sky130_fd_sc_hd__a211oi_1 _2236_ (.A1(_0644_),
    .A2(_0428_),
    .B1(_0429_),
    .C1(_1135_),
    .Y(_0430_));
 sky130_fd_sc_hd__a21o_1 _2237_ (.A1(_0699_),
    .A2(_0697_),
    .B1(_0707_),
    .X(_0431_));
 sky130_fd_sc_hd__a311oi_2 _2238_ (.A1(_0700_),
    .A2(_0702_),
    .A3(_0431_),
    .B1(_0937_),
    .C1(_1090_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _2239_ (.A(_0669_),
    .B(_0668_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_1 _2240_ (.A(_0598_),
    .B(_1131_),
    .Y(_0434_));
 sky130_fd_sc_hd__a211oi_1 _2241_ (.A1(_0667_),
    .A2(_0433_),
    .B1(_0434_),
    .C1(_1120_),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_1 _2242_ (.A(_0676_),
    .Y(_0436_));
 sky130_fd_sc_hd__a21o_1 _2243_ (.A1(_0436_),
    .A2(_0674_),
    .B1(_0731_),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_1 _2244_ (.A(_0602_),
    .B(_1116_),
    .Y(_0438_));
 sky130_fd_sc_hd__a211oi_1 _2245_ (.A1(_0268_),
    .A2(_0437_),
    .B1(_0438_),
    .C1(_1105_),
    .Y(_0439_));
 sky130_fd_sc_hd__nor4_1 _2246_ (.A(_0430_),
    .B(_0432_),
    .C(_0435_),
    .D(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__o41ai_1 _2247_ (.A1(_1150_),
    .A2(_1148_),
    .A3(_0621_),
    .A4(_0427_),
    .B1(_0440_),
    .Y(net300));
 sky130_fd_sc_hd__nand2_1 _2248_ (.A(_0598_),
    .B(_1125_),
    .Y(_0441_));
 sky130_fd_sc_hd__a211o_2 _2249_ (.A1(_0669_),
    .A2(_0658_),
    .B1(_0441_),
    .C1(_0656_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_4 _2250_ (.A(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__o2111a_2 _2251_ (.A1(_0675_),
    .A2(_0678_),
    .B1(_0600_),
    .C1(_1110_),
    .D1(_0679_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_4 _2252_ (.A(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a211oi_4 _2253_ (.A1(_0669_),
    .A2(_0658_),
    .B1(_0441_),
    .C1(_0656_),
    .Y(_0446_));
 sky130_fd_sc_hd__a21o_1 _2254_ (.A1(\input_buffer[1][0] ),
    .A2(_0445_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__o211ai_4 _2255_ (.A1(_0698_),
    .A2(_0707_),
    .B1(_1092_),
    .C1(_0702_),
    .Y(_0448_));
 sky130_fd_sc_hd__clkbuf_4 _2256_ (.A(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__buf_4 _2257_ (.A(_0444_),
    .X(_0450_));
 sky130_fd_sc_hd__nor3_1 _2258_ (.A(_0728_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand3_2 _2259_ (.A(_0637_),
    .B(_1140_),
    .C(_1144_),
    .Y(_0452_));
 sky130_fd_sc_hd__o221ai_1 _2260_ (.A1(\input_buffer[2][0] ),
    .A2(_0443_),
    .B1(_0447_),
    .B2(_0451_),
    .C1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__and3_1 _2261_ (.A(_0597_),
    .B(_1140_),
    .C(_1144_),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _2262_ (.A(\input_buffer_valid[4] ),
    .B(_1155_),
    .Y(_0455_));
 sky130_fd_sc_hd__a211oi_4 _2263_ (.A1(_0619_),
    .A2(_0615_),
    .B1(_0455_),
    .C1(_0613_),
    .Y(_0456_));
 sky130_fd_sc_hd__clkbuf_4 _2264_ (.A(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__a21oi_1 _2265_ (.A1(\input_buffer[3][0] ),
    .A2(_0454_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__a211o_1 _2266_ (.A1(_0619_),
    .A2(_0615_),
    .B1(_0455_),
    .C1(_0613_),
    .X(_0459_));
 sky130_fd_sc_hd__nor2_1 _2267_ (.A(\input_buffer[4][0] ),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _2268_ (.A1(_0453_),
    .A2(_0458_),
    .B1(_0460_),
    .Y(net302));
 sky130_fd_sc_hd__clkbuf_4 _2269_ (.A(_0444_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_4 _2270_ (.A(_0446_),
    .X(_0462_));
 sky130_fd_sc_hd__nor3_1 _2271_ (.A(_0748_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0463_));
 sky130_fd_sc_hd__a211oi_1 _2272_ (.A1(\input_buffer[1][10] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__clkbuf_4 _2273_ (.A(_0442_),
    .X(_0465_));
 sky130_fd_sc_hd__o2111ai_4 _2274_ (.A1(_0735_),
    .A2(_0642_),
    .B1(_0597_),
    .C1(_1140_),
    .D1(_0633_),
    .Y(_0466_));
 sky130_fd_sc_hd__and2_2 _2275_ (.A(_0459_),
    .B(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_4 _2276_ (.A(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__o21ai_0 _2277_ (.A1(\input_buffer[2][10] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_8 _2278_ (.A(_0456_),
    .B(_0466_),
    .Y(_0470_));
 sky130_fd_sc_hd__buf_6 _2279_ (.A(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a22oi_1 _2280_ (.A1(\input_buffer[4][10] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][10] ),
    .Y(_0472_));
 sky130_fd_sc_hd__o21ai_1 _2281_ (.A1(_0464_),
    .A2(_0469_),
    .B1(_0472_),
    .Y(net303));
 sky130_fd_sc_hd__nor3_1 _2282_ (.A(_0755_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0473_));
 sky130_fd_sc_hd__a211oi_1 _2283_ (.A1(\input_buffer[1][11] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21ai_0 _2284_ (.A1(\input_buffer[2][11] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0475_));
 sky130_fd_sc_hd__a22oi_1 _2285_ (.A1(\input_buffer[4][11] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][11] ),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_1 _2286_ (.A1(_0474_),
    .A2(_0475_),
    .B1(_0476_),
    .Y(net304));
 sky130_fd_sc_hd__nor3_1 _2287_ (.A(_0761_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0477_));
 sky130_fd_sc_hd__a211oi_1 _2288_ (.A1(\input_buffer[1][12] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__o21ai_0 _2289_ (.A1(\input_buffer[2][12] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0479_));
 sky130_fd_sc_hd__a22oi_1 _2290_ (.A1(\input_buffer[4][12] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][12] ),
    .Y(_0480_));
 sky130_fd_sc_hd__o21ai_1 _2291_ (.A1(_0478_),
    .A2(_0479_),
    .B1(_0480_),
    .Y(net305));
 sky130_fd_sc_hd__nor3_1 _2292_ (.A(_0769_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0481_));
 sky130_fd_sc_hd__a21o_1 _2293_ (.A1(\input_buffer[1][13] ),
    .A2(_0445_),
    .B1(_0446_),
    .X(_0482_));
 sky130_fd_sc_hd__o221ai_1 _2294_ (.A1(\input_buffer[2][13] ),
    .A2(_0443_),
    .B1(_0481_),
    .B2(_0482_),
    .C1(_0452_),
    .Y(_0483_));
 sky130_fd_sc_hd__a21oi_1 _2295_ (.A1(\input_buffer[3][13] ),
    .A2(_0454_),
    .B1(_0457_),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_1 _2296_ (.A(\input_buffer[4][13] ),
    .B(_0459_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _2297_ (.A1(_0483_),
    .A2(_0484_),
    .B1(_0485_),
    .Y(net306));
 sky130_fd_sc_hd__nor3_1 _2298_ (.A(_0776_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0486_));
 sky130_fd_sc_hd__a211oi_1 _2299_ (.A1(\input_buffer[1][14] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__o21ai_0 _2300_ (.A1(\input_buffer[2][14] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0488_));
 sky130_fd_sc_hd__a22oi_1 _2301_ (.A1(\input_buffer[4][14] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][14] ),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _2302_ (.A1(_0487_),
    .A2(_0488_),
    .B1(_0489_),
    .Y(net307));
 sky130_fd_sc_hd__nor3_1 _2303_ (.A(_0782_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0490_));
 sky130_fd_sc_hd__a211oi_1 _2304_ (.A1(\input_buffer[1][15] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__o21ai_0 _2305_ (.A1(\input_buffer[2][15] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0492_));
 sky130_fd_sc_hd__a22oi_1 _2306_ (.A1(\input_buffer[4][15] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][15] ),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_1 _2307_ (.A1(_0491_),
    .A2(_0492_),
    .B1(_0493_),
    .Y(net308));
 sky130_fd_sc_hd__nor3_1 _2308_ (.A(_0788_),
    .B(_0449_),
    .C(_0450_),
    .Y(_0494_));
 sky130_fd_sc_hd__a211oi_1 _2309_ (.A1(\input_buffer[1][16] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__o21ai_0 _2310_ (.A1(\input_buffer[2][16] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0496_));
 sky130_fd_sc_hd__a22oi_1 _2311_ (.A1(\input_buffer[4][16] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][16] ),
    .Y(_0497_));
 sky130_fd_sc_hd__o21ai_1 _2312_ (.A1(_0495_),
    .A2(_0496_),
    .B1(_0497_),
    .Y(net309));
 sky130_fd_sc_hd__clkbuf_4 _2313_ (.A(_0444_),
    .X(_0498_));
 sky130_fd_sc_hd__nor3_1 _2314_ (.A(_0794_),
    .B(_0449_),
    .C(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__a211oi_1 _2315_ (.A1(\input_buffer[1][17] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_0 _2316_ (.A1(\input_buffer[2][17] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0501_));
 sky130_fd_sc_hd__a22oi_1 _2317_ (.A1(\input_buffer[4][17] ),
    .A2(_0457_),
    .B1(_0471_),
    .B2(\input_buffer[3][17] ),
    .Y(_0502_));
 sky130_fd_sc_hd__o21ai_1 _2318_ (.A1(_0500_),
    .A2(_0501_),
    .B1(_0502_),
    .Y(net310));
 sky130_fd_sc_hd__nor3_1 _2319_ (.A(_0802_),
    .B(_0449_),
    .C(_0498_),
    .Y(_0503_));
 sky130_fd_sc_hd__a211oi_1 _2320_ (.A1(\input_buffer[1][18] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__o21ai_0 _2321_ (.A1(\input_buffer[2][18] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0505_));
 sky130_fd_sc_hd__buf_4 _2322_ (.A(_0456_),
    .X(_0506_));
 sky130_fd_sc_hd__a22oi_1 _2323_ (.A1(\input_buffer[4][18] ),
    .A2(_0506_),
    .B1(_0471_),
    .B2(\input_buffer[3][18] ),
    .Y(_0507_));
 sky130_fd_sc_hd__o21ai_1 _2324_ (.A1(_0504_),
    .A2(_0505_),
    .B1(_0507_),
    .Y(net311));
 sky130_fd_sc_hd__clkbuf_4 _2325_ (.A(_0448_),
    .X(_0508_));
 sky130_fd_sc_hd__nor3_1 _2326_ (.A(_0812_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0509_));
 sky130_fd_sc_hd__a211oi_1 _2327_ (.A1(\input_buffer[1][19] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21ai_0 _2328_ (.A1(\input_buffer[2][19] ),
    .A2(_0465_),
    .B1(_0468_),
    .Y(_0511_));
 sky130_fd_sc_hd__a22oi_1 _2329_ (.A1(\input_buffer[4][19] ),
    .A2(_0506_),
    .B1(_0471_),
    .B2(\input_buffer[3][19] ),
    .Y(_0512_));
 sky130_fd_sc_hd__o21ai_1 _2330_ (.A1(_0510_),
    .A2(_0511_),
    .B1(_0512_),
    .Y(net312));
 sky130_fd_sc_hd__nor3_1 _2331_ (.A(_0821_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0513_));
 sky130_fd_sc_hd__a211oi_1 _2332_ (.A1(\input_buffer[1][1] ),
    .A2(_0461_),
    .B1(_0462_),
    .C1(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _2333_ (.A(_0467_),
    .X(_0515_));
 sky130_fd_sc_hd__o21ai_0 _2334_ (.A1(\input_buffer[2][1] ),
    .A2(_0465_),
    .B1(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__a22oi_1 _2335_ (.A1(\input_buffer[4][1] ),
    .A2(_0506_),
    .B1(_0471_),
    .B2(\input_buffer[3][1] ),
    .Y(_0517_));
 sky130_fd_sc_hd__o21ai_1 _2336_ (.A1(_0514_),
    .A2(_0516_),
    .B1(_0517_),
    .Y(net313));
 sky130_fd_sc_hd__clkbuf_4 _2337_ (.A(_0444_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_4 _2338_ (.A(_0446_),
    .X(_0519_));
 sky130_fd_sc_hd__nor3_1 _2339_ (.A(_0827_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0520_));
 sky130_fd_sc_hd__a211oi_1 _2340_ (.A1(\input_buffer[1][20] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__clkbuf_4 _2341_ (.A(_0442_),
    .X(_0522_));
 sky130_fd_sc_hd__o21ai_0 _2342_ (.A1(\input_buffer[2][20] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0523_));
 sky130_fd_sc_hd__buf_6 _2343_ (.A(_0470_),
    .X(_0524_));
 sky130_fd_sc_hd__a22oi_1 _2344_ (.A1(\input_buffer[4][20] ),
    .A2(_0506_),
    .B1(_0524_),
    .B2(\input_buffer[3][20] ),
    .Y(_0525_));
 sky130_fd_sc_hd__o21ai_0 _2345_ (.A1(_0521_),
    .A2(_0523_),
    .B1(_0525_),
    .Y(net314));
 sky130_fd_sc_hd__nor3_1 _2346_ (.A(_0833_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0526_));
 sky130_fd_sc_hd__a211oi_1 _2347_ (.A1(\input_buffer[1][21] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21ai_0 _2348_ (.A1(\input_buffer[2][21] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0528_));
 sky130_fd_sc_hd__a22oi_1 _2349_ (.A1(\input_buffer[4][21] ),
    .A2(_0506_),
    .B1(_0524_),
    .B2(\input_buffer[3][21] ),
    .Y(_0529_));
 sky130_fd_sc_hd__o21ai_0 _2350_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0529_),
    .Y(net315));
 sky130_fd_sc_hd__nor3_1 _2351_ (.A(_0841_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0530_));
 sky130_fd_sc_hd__a211oi_1 _2352_ (.A1(\input_buffer[1][22] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__o21ai_0 _2353_ (.A1(\input_buffer[2][22] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0532_));
 sky130_fd_sc_hd__a22oi_1 _2354_ (.A1(\input_buffer[4][22] ),
    .A2(_0506_),
    .B1(_0524_),
    .B2(\input_buffer[3][22] ),
    .Y(_0533_));
 sky130_fd_sc_hd__o21ai_0 _2355_ (.A1(_0531_),
    .A2(_0532_),
    .B1(_0533_),
    .Y(net316));
 sky130_fd_sc_hd__nor3_1 _2356_ (.A(_0847_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0534_));
 sky130_fd_sc_hd__a211oi_1 _2357_ (.A1(\input_buffer[1][23] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_0 _2358_ (.A1(\input_buffer[2][23] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0536_));
 sky130_fd_sc_hd__a22oi_1 _2359_ (.A1(\input_buffer[4][23] ),
    .A2(_0506_),
    .B1(_0524_),
    .B2(\input_buffer[3][23] ),
    .Y(_0537_));
 sky130_fd_sc_hd__o21ai_1 _2360_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_0537_),
    .Y(net317));
 sky130_fd_sc_hd__nor3b_1 _2361_ (.A(_0445_),
    .B(_0855_),
    .C_N(_1092_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand3_1 _2362_ (.A(_0602_),
    .B(_0676_),
    .C(_1110_),
    .Y(_0539_));
 sky130_fd_sc_hd__o21ai_0 _2363_ (.A1(_0682_),
    .A2(_0539_),
    .B1(_0443_),
    .Y(_0540_));
 sky130_fd_sc_hd__o221ai_1 _2364_ (.A1(_0650_),
    .A2(_0443_),
    .B1(_0538_),
    .B2(_0540_),
    .C1(_0452_),
    .Y(_0541_));
 sky130_fd_sc_hd__a21oi_1 _2365_ (.A1(_0634_),
    .A2(_0454_),
    .B1(_0457_),
    .Y(_0542_));
 sky130_fd_sc_hd__nor2_1 _2366_ (.A(_0606_),
    .B(_0459_),
    .Y(_0543_));
 sky130_fd_sc_hd__a21oi_1 _2367_ (.A1(_0541_),
    .A2(_0542_),
    .B1(_0543_),
    .Y(net318));
 sky130_fd_sc_hd__o2111ai_4 _2368_ (.A1(_0730_),
    .A2(_0685_),
    .B1(_0600_),
    .C1(_1110_),
    .D1(_0683_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand3_1 _2369_ (.A(_0857_),
    .B(_0673_),
    .C(_1110_),
    .Y(_0545_));
 sky130_fd_sc_hd__o21ai_1 _2370_ (.A1(_0682_),
    .A2(_0545_),
    .B1(_0443_),
    .Y(_0546_));
 sky130_fd_sc_hd__a31oi_2 _2371_ (.A1(_1092_),
    .A2(_0376_),
    .A3(_0544_),
    .B1(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__o21ai_0 _2372_ (.A1(\dest_id[2][1] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0548_));
 sky130_fd_sc_hd__a22oi_1 _2373_ (.A1(_0604_),
    .A2(_0506_),
    .B1(_0524_),
    .B2(_0627_),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_2 _2374_ (.A1(_0547_),
    .A2(_0548_),
    .B1(_0549_),
    .Y(net319));
 sky130_fd_sc_hd__nand3_1 _2375_ (.A(_0857_),
    .B(_0674_),
    .C(_1110_),
    .Y(_0550_));
 sky130_fd_sc_hd__o21ai_0 _2376_ (.A1(_0682_),
    .A2(_0550_),
    .B1(_0443_),
    .Y(_0551_));
 sky130_fd_sc_hd__a31oi_1 _2377_ (.A1(_1092_),
    .A2(_0383_),
    .A3(_0544_),
    .B1(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__o21ai_1 _2378_ (.A1(_0649_),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0553_));
 sky130_fd_sc_hd__a21oi_1 _2379_ (.A1(_0628_),
    .A2(_0470_),
    .B1(_0543_),
    .Y(_0554_));
 sky130_fd_sc_hd__o21ai_1 _2380_ (.A1(_0552_),
    .A2(_0553_),
    .B1(_0554_),
    .Y(net320));
 sky130_fd_sc_hd__nand2_1 _2381_ (.A(_0677_),
    .B(_0445_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand4_1 _2382_ (.A(_1092_),
    .B(_0703_),
    .C(_0882_),
    .D(_0544_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_1 _2383_ (.A(_0652_),
    .B(_0442_),
    .Y(_0557_));
 sky130_fd_sc_hd__a31o_1 _2384_ (.A1(_0442_),
    .A2(_0555_),
    .A3(_0556_),
    .B1(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _2385_ (.A(_0608_),
    .B(_0459_),
    .Y(_0559_));
 sky130_fd_sc_hd__a221oi_2 _2386_ (.A1(_0886_),
    .A2(_0470_),
    .B1(_0558_),
    .B2(_0468_),
    .C1(_0559_),
    .Y(net321));
 sky130_fd_sc_hd__nor3_1 _2387_ (.A(_0889_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0560_));
 sky130_fd_sc_hd__a211oi_1 _2388_ (.A1(\input_buffer[1][2] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__o21ai_0 _2389_ (.A1(\input_buffer[2][2] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0562_));
 sky130_fd_sc_hd__a22oi_1 _2390_ (.A1(\input_buffer[4][2] ),
    .A2(_0506_),
    .B1(_0524_),
    .B2(\input_buffer[3][2] ),
    .Y(_0563_));
 sky130_fd_sc_hd__o21ai_0 _2391_ (.A1(_0561_),
    .A2(_0562_),
    .B1(_0563_),
    .Y(net322));
 sky130_fd_sc_hd__nor3_1 _2392_ (.A(_0895_),
    .B(_0508_),
    .C(_0498_),
    .Y(_0564_));
 sky130_fd_sc_hd__a211oi_1 _2393_ (.A1(\input_buffer[1][3] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21ai_0 _2394_ (.A1(\input_buffer[2][3] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0566_));
 sky130_fd_sc_hd__a22oi_1 _2395_ (.A1(\input_buffer[4][3] ),
    .A2(_0506_),
    .B1(_0524_),
    .B2(\input_buffer[3][3] ),
    .Y(_0567_));
 sky130_fd_sc_hd__o21ai_0 _2396_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0567_),
    .Y(net323));
 sky130_fd_sc_hd__nor3_1 _2397_ (.A(_0901_),
    .B(_0508_),
    .C(_0445_),
    .Y(_0568_));
 sky130_fd_sc_hd__a211oi_1 _2398_ (.A1(\input_buffer[1][4] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__o21ai_0 _2399_ (.A1(\input_buffer[2][4] ),
    .A2(_0522_),
    .B1(_0515_),
    .Y(_0570_));
 sky130_fd_sc_hd__a22oi_1 _2400_ (.A1(\input_buffer[4][4] ),
    .A2(_0456_),
    .B1(_0524_),
    .B2(\input_buffer[3][4] ),
    .Y(_0571_));
 sky130_fd_sc_hd__o21ai_0 _2401_ (.A1(_0569_),
    .A2(_0570_),
    .B1(_0571_),
    .Y(net324));
 sky130_fd_sc_hd__nor3_1 _2402_ (.A(_0907_),
    .B(_0508_),
    .C(_0445_),
    .Y(_0572_));
 sky130_fd_sc_hd__a211oi_1 _2403_ (.A1(\input_buffer[1][5] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21ai_0 _2404_ (.A1(\input_buffer[2][5] ),
    .A2(_0522_),
    .B1(_0467_),
    .Y(_0574_));
 sky130_fd_sc_hd__a22oi_1 _2405_ (.A1(\input_buffer[4][5] ),
    .A2(_0456_),
    .B1(_0524_),
    .B2(\input_buffer[3][5] ),
    .Y(_0575_));
 sky130_fd_sc_hd__o21ai_0 _2406_ (.A1(_0573_),
    .A2(_0574_),
    .B1(_0575_),
    .Y(net325));
 sky130_fd_sc_hd__nor3_1 _2407_ (.A(_0913_),
    .B(_0448_),
    .C(_0445_),
    .Y(_0576_));
 sky130_fd_sc_hd__a211oi_1 _2408_ (.A1(\input_buffer[1][6] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__o21ai_0 _2409_ (.A1(\input_buffer[2][6] ),
    .A2(_0443_),
    .B1(_0467_),
    .Y(_0578_));
 sky130_fd_sc_hd__a22oi_1 _2410_ (.A1(\input_buffer[4][6] ),
    .A2(_0456_),
    .B1(_0524_),
    .B2(\input_buffer[3][6] ),
    .Y(_0579_));
 sky130_fd_sc_hd__o21ai_0 _2411_ (.A1(_0577_),
    .A2(_0578_),
    .B1(_0579_),
    .Y(net326));
 sky130_fd_sc_hd__nor3_1 _2412_ (.A(_0919_),
    .B(_0448_),
    .C(_0445_),
    .Y(_0580_));
 sky130_fd_sc_hd__a211oi_1 _2413_ (.A1(\input_buffer[1][7] ),
    .A2(_0518_),
    .B1(_0519_),
    .C1(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__o21ai_0 _2414_ (.A1(\input_buffer[2][7] ),
    .A2(_0443_),
    .B1(_0467_),
    .Y(_0582_));
 sky130_fd_sc_hd__a22oi_1 _2415_ (.A1(\input_buffer[4][7] ),
    .A2(_0456_),
    .B1(_0470_),
    .B2(\input_buffer[3][7] ),
    .Y(_0583_));
 sky130_fd_sc_hd__o21ai_1 _2416_ (.A1(_0581_),
    .A2(_0582_),
    .B1(_0583_),
    .Y(net327));
 sky130_fd_sc_hd__nor3_1 _2417_ (.A(_0925_),
    .B(_0448_),
    .C(_0445_),
    .Y(_0584_));
 sky130_fd_sc_hd__a211oi_1 _2418_ (.A1(\input_buffer[1][8] ),
    .A2(_0450_),
    .B1(_0446_),
    .C1(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__o21ai_0 _2419_ (.A1(\input_buffer[2][8] ),
    .A2(_0443_),
    .B1(_0467_),
    .Y(_0586_));
 sky130_fd_sc_hd__a22oi_1 _2420_ (.A1(\input_buffer[4][8] ),
    .A2(_0456_),
    .B1(_0470_),
    .B2(\input_buffer[3][8] ),
    .Y(_0587_));
 sky130_fd_sc_hd__o21ai_1 _2421_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0587_),
    .Y(net328));
 sky130_fd_sc_hd__nor3_1 _2422_ (.A(_0931_),
    .B(_0448_),
    .C(_0445_),
    .Y(_0588_));
 sky130_fd_sc_hd__a211oi_1 _2423_ (.A1(\input_buffer[1][9] ),
    .A2(_0450_),
    .B1(_0446_),
    .C1(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__o21ai_0 _2424_ (.A1(\input_buffer[2][9] ),
    .A2(_0443_),
    .B1(_0467_),
    .Y(_0590_));
 sky130_fd_sc_hd__a22oi_1 _2425_ (.A1(\input_buffer[4][9] ),
    .A2(_0456_),
    .B1(_0470_),
    .B2(\input_buffer[3][9] ),
    .Y(_0591_));
 sky130_fd_sc_hd__o21ai_1 _2426_ (.A1(_0589_),
    .A2(_0590_),
    .B1(_0591_),
    .Y(net329));
 sky130_fd_sc_hd__nand3_1 _2427_ (.A(_0625_),
    .B(_1161_),
    .C(_1155_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand3_1 _2428_ (.A(_0599_),
    .B(_1131_),
    .C(_1125_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand3_1 _2429_ (.A(_0714_),
    .B(_1101_),
    .C(_1092_),
    .Y(_0594_));
 sky130_fd_sc_hd__and3_1 _2430_ (.A(_0602_),
    .B(_1116_),
    .C(_1110_),
    .X(_0595_));
 sky130_fd_sc_hd__a31oi_1 _2431_ (.A1(_0637_),
    .A2(_1146_),
    .A3(_1140_),
    .B1(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand4_1 _2432_ (.A(_0592_),
    .B(_0593_),
    .C(_0594_),
    .D(_0596_),
    .Y(net330));
 sky130_fd_sc_hd__ha_2 _2433_ (.A(_1087_),
    .B(_1088_),
    .COUT(_1089_),
    .SUM(_1090_));
 sky130_fd_sc_hd__ha_4 _2434_ (.A(_1087_),
    .B(_1091_),
    .COUT(_1092_),
    .SUM(_1093_));
 sky130_fd_sc_hd__ha_1 _2435_ (.A(_1094_),
    .B(_1088_),
    .COUT(_1095_),
    .SUM(_1096_));
 sky130_fd_sc_hd__ha_2 _2436_ (.A(_1094_),
    .B(_1091_),
    .COUT(_1097_),
    .SUM(_1098_));
 sky130_fd_sc_hd__ha_1 _2437_ (.A(_1095_),
    .B(_1099_),
    .COUT(_1100_),
    .SUM(_1101_));
 sky130_fd_sc_hd__ha_2 _2438_ (.A(_1102_),
    .B(_1103_),
    .COUT(_1104_),
    .SUM(_1105_));
 sky130_fd_sc_hd__ha_1 _2439_ (.A(_1102_),
    .B(_1106_),
    .COUT(_1107_),
    .SUM(_1108_));
 sky130_fd_sc_hd__ha_4 _2440_ (.A(_1109_),
    .B(_1103_),
    .COUT(_1110_),
    .SUM(_1111_));
 sky130_fd_sc_hd__ha_2 _2441_ (.A(_1109_),
    .B(_1106_),
    .COUT(_1112_),
    .SUM(_1113_));
 sky130_fd_sc_hd__ha_1 _2442_ (.A(_1107_),
    .B(_1114_),
    .COUT(_1115_),
    .SUM(_1116_));
 sky130_fd_sc_hd__ha_1 _2443_ (.A(_1117_),
    .B(_1118_),
    .COUT(_1119_),
    .SUM(_1120_));
 sky130_fd_sc_hd__ha_1 _2444_ (.A(_1117_),
    .B(_1121_),
    .COUT(_1122_),
    .SUM(_1123_));
 sky130_fd_sc_hd__ha_1 _2445_ (.A(_1124_),
    .B(_1118_),
    .COUT(_1125_),
    .SUM(_1126_));
 sky130_fd_sc_hd__ha_1 _2446_ (.A(_1124_),
    .B(_1121_),
    .COUT(_1127_),
    .SUM(_1128_));
 sky130_fd_sc_hd__ha_2 _2447_ (.A(_1122_),
    .B(_1129_),
    .COUT(_1130_),
    .SUM(_1131_));
 sky130_fd_sc_hd__ha_1 _2448_ (.A(_1132_),
    .B(_1133_),
    .COUT(_1134_),
    .SUM(_1135_));
 sky130_fd_sc_hd__ha_1 _2449_ (.A(_1132_),
    .B(_1136_),
    .COUT(_1137_),
    .SUM(_1138_));
 sky130_fd_sc_hd__ha_2 _2450_ (.A(_1139_),
    .B(_1133_),
    .COUT(_1140_),
    .SUM(_1141_));
 sky130_fd_sc_hd__ha_1 _2451_ (.A(_1139_),
    .B(_1136_),
    .COUT(_1142_),
    .SUM(_1143_));
 sky130_fd_sc_hd__ha_1 _2452_ (.A(_1137_),
    .B(_1144_),
    .COUT(_1145_),
    .SUM(_1146_));
 sky130_fd_sc_hd__ha_1 _2453_ (.A(_1147_),
    .B(_1148_),
    .COUT(_1149_),
    .SUM(_1150_));
 sky130_fd_sc_hd__ha_1 _2454_ (.A(_1147_),
    .B(_1151_),
    .COUT(_1152_),
    .SUM(_1153_));
 sky130_fd_sc_hd__ha_1 _2455_ (.A(_1154_),
    .B(_1148_),
    .COUT(_1155_),
    .SUM(_1156_));
 sky130_fd_sc_hd__ha_1 _2456_ (.A(_1154_),
    .B(_1151_),
    .COUT(_1157_),
    .SUM(_1158_));
 sky130_fd_sc_hd__ha_1 _2457_ (.A(_1152_),
    .B(_1159_),
    .COUT(_1160_),
    .SUM(_1161_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_4 _2459_ (.A(net331),
    .X(east_out_data[28]));
 sky130_fd_sc_hd__buf_4 _2460_ (.A(net332),
    .X(east_out_data[29]));
 sky130_fd_sc_hd__buf_4 _2461_ (.A(net333),
    .X(east_out_data[30]));
 sky130_fd_sc_hd__buf_4 _2462_ (.A(net334),
    .X(east_out_data[31]));
 sky130_fd_sc_hd__buf_4 _2463_ (.A(net335),
    .X(south_out_data[28]));
 sky130_fd_sc_hd__buf_4 _2464_ (.A(net336),
    .X(south_out_data[29]));
 sky130_fd_sc_hd__buf_4 _2465_ (.A(net337),
    .X(south_out_data[30]));
 sky130_fd_sc_hd__buf_4 _2466_ (.A(net338),
    .X(south_out_data[31]));
 sky130_fd_sc_hd__buf_4 _2467_ (.A(net339),
    .X(west_out_data[28]));
 sky130_fd_sc_hd__buf_4 _2468_ (.A(net340),
    .X(west_out_data[29]));
 sky130_fd_sc_hd__buf_4 _2469_ (.A(net341),
    .X(west_out_data[30]));
 sky130_fd_sc_hd__buf_4 _2470_ (.A(net342),
    .X(west_out_data[31]));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][0]$_DFFE_PP_  (.D(net70),
    .DE(_0009_),
    .Q(\input_buffer[0][0] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][10]$_DFFE_PP_  (.D(net71),
    .DE(_0009_),
    .Q(\input_buffer[0][10] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][11]$_DFFE_PP_  (.D(net72),
    .DE(_0009_),
    .Q(\input_buffer[0][11] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][12]$_DFFE_PP_  (.D(net73),
    .DE(_0009_),
    .Q(\input_buffer[0][12] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][13]$_DFFE_PP_  (.D(net74),
    .DE(_0009_),
    .Q(\input_buffer[0][13] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][14]$_DFFE_PP_  (.D(net75),
    .DE(_0009_),
    .Q(\input_buffer[0][14] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][15]$_DFFE_PP_  (.D(net76),
    .DE(_0009_),
    .Q(\input_buffer[0][15] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][16]$_DFFE_PP_  (.D(net77),
    .DE(_0009_),
    .Q(\input_buffer[0][16] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][17]$_DFFE_PP_  (.D(net78),
    .DE(_0009_),
    .Q(\input_buffer[0][17] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][18]$_DFFE_PP_  (.D(net79),
    .DE(_0009_),
    .Q(\input_buffer[0][18] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][19]$_DFFE_PP_  (.D(net80),
    .DE(_0009_),
    .Q(\input_buffer[0][19] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][1]$_DFFE_PP_  (.D(net81),
    .DE(_0009_),
    .Q(\input_buffer[0][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][20]$_DFFE_PP_  (.D(net82),
    .DE(_0009_),
    .Q(\input_buffer[0][20] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][21]$_DFFE_PP_  (.D(net83),
    .DE(_0009_),
    .Q(\input_buffer[0][21] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][22]$_DFFE_PP_  (.D(net84),
    .DE(_0009_),
    .Q(\input_buffer[0][22] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][23]$_DFFE_PP_  (.D(net85),
    .DE(_0009_),
    .Q(\input_buffer[0][23] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][24]$_DFFE_PP_  (.D(net86),
    .DE(_0009_),
    .Q(\dest_id[0][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][25]$_DFFE_PP_  (.D(net87),
    .DE(_0009_),
    .Q(\dest_id[0][1] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][26]$_DFFE_PP_  (.D(net88),
    .DE(_0009_),
    .Q(\dest_id[0][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][27]$_DFFE_PP_  (.D(net89),
    .DE(_0009_),
    .Q(\dest_id[0][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][28]$_DFFE_PP_  (.D(net90),
    .DE(_0009_),
    .Q(\dest_id[0][4] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][29]$_DFFE_PP_  (.D(net91),
    .DE(_0009_),
    .Q(\dest_id[0][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][2]$_DFFE_PP_  (.D(net92),
    .DE(_0009_),
    .Q(\input_buffer[0][2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][30]$_DFFE_PP_  (.D(net93),
    .DE(_0009_),
    .Q(\dest_id[0][6] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][31]$_DFFE_PP_  (.D(net94),
    .DE(_0009_),
    .Q(\dest_id[0][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][3]$_DFFE_PP_  (.D(net95),
    .DE(_0009_),
    .Q(\input_buffer[0][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][4]$_DFFE_PP_  (.D(net96),
    .DE(_0009_),
    .Q(\input_buffer[0][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][5]$_DFFE_PP_  (.D(net97),
    .DE(_0009_),
    .Q(\input_buffer[0][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][6]$_DFFE_PP_  (.D(net98),
    .DE(_0009_),
    .Q(\input_buffer[0][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][7]$_DFFE_PP_  (.D(net99),
    .DE(_0009_),
    .Q(\input_buffer[0][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][8]$_DFFE_PP_  (.D(net100),
    .DE(_0009_),
    .Q(\input_buffer[0][8] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[0][9]$_DFFE_PP_  (.D(net101),
    .DE(_0009_),
    .Q(\input_buffer[0][9] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][0]$_DFFE_PP_  (.D(net2),
    .DE(_0008_),
    .Q(\input_buffer[1][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][10]$_DFFE_PP_  (.D(net3),
    .DE(_0008_),
    .Q(\input_buffer[1][10] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][11]$_DFFE_PP_  (.D(net4),
    .DE(_0008_),
    .Q(\input_buffer[1][11] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][12]$_DFFE_PP_  (.D(net5),
    .DE(_0008_),
    .Q(\input_buffer[1][12] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][13]$_DFFE_PP_  (.D(net6),
    .DE(_0008_),
    .Q(\input_buffer[1][13] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][14]$_DFFE_PP_  (.D(net7),
    .DE(_0008_),
    .Q(\input_buffer[1][14] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][15]$_DFFE_PP_  (.D(net8),
    .DE(_0008_),
    .Q(\input_buffer[1][15] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][16]$_DFFE_PP_  (.D(net9),
    .DE(_0008_),
    .Q(\input_buffer[1][16] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][17]$_DFFE_PP_  (.D(net10),
    .DE(_0008_),
    .Q(\input_buffer[1][17] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][18]$_DFFE_PP_  (.D(net11),
    .DE(_0008_),
    .Q(\input_buffer[1][18] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][19]$_DFFE_PP_  (.D(net12),
    .DE(_0008_),
    .Q(\input_buffer[1][19] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][1]$_DFFE_PP_  (.D(net13),
    .DE(_0008_),
    .Q(\input_buffer[1][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][20]$_DFFE_PP_  (.D(net14),
    .DE(_0008_),
    .Q(\input_buffer[1][20] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][21]$_DFFE_PP_  (.D(net15),
    .DE(_0008_),
    .Q(\input_buffer[1][21] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][22]$_DFFE_PP_  (.D(net16),
    .DE(_0008_),
    .Q(\input_buffer[1][22] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][23]$_DFFE_PP_  (.D(net17),
    .DE(_0008_),
    .Q(\input_buffer[1][23] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][24]$_DFFE_PP_  (.D(net18),
    .DE(_0008_),
    .Q(\dest_id[1][0] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][25]$_DFFE_PP_  (.D(net19),
    .DE(_0008_),
    .Q(\dest_id[1][1] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][26]$_DFFE_PP_  (.D(net20),
    .DE(_0008_),
    .Q(\dest_id[1][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][27]$_DFFE_PP_  (.D(net21),
    .DE(_0008_),
    .Q(\dest_id[1][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][28]$_DFFE_PP_  (.D(net22),
    .DE(_0008_),
    .Q(\dest_id[1][4] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][29]$_DFFE_PP_  (.D(net23),
    .DE(_0008_),
    .Q(\dest_id[1][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][2]$_DFFE_PP_  (.D(net24),
    .DE(_0008_),
    .Q(\input_buffer[1][2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][30]$_DFFE_PP_  (.D(net25),
    .DE(_0008_),
    .Q(\dest_id[1][6] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][31]$_DFFE_PP_  (.D(net26),
    .DE(_0008_),
    .Q(\dest_id[1][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][3]$_DFFE_PP_  (.D(net27),
    .DE(_0008_),
    .Q(\input_buffer[1][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][4]$_DFFE_PP_  (.D(net28),
    .DE(_0008_),
    .Q(\input_buffer[1][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][5]$_DFFE_PP_  (.D(net29),
    .DE(_0008_),
    .Q(\input_buffer[1][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][6]$_DFFE_PP_  (.D(net30),
    .DE(_0008_),
    .Q(\input_buffer[1][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][7]$_DFFE_PP_  (.D(net31),
    .DE(_0008_),
    .Q(\input_buffer[1][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][8]$_DFFE_PP_  (.D(net32),
    .DE(_0008_),
    .Q(\input_buffer[1][8] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[1][9]$_DFFE_PP_  (.D(net33),
    .DE(_0008_),
    .Q(\input_buffer[1][9] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][0]$_DFFE_PP_  (.D(net105),
    .DE(_0007_),
    .Q(\input_buffer[2][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][10]$_DFFE_PP_  (.D(net106),
    .DE(_0007_),
    .Q(\input_buffer[2][10] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][11]$_DFFE_PP_  (.D(net107),
    .DE(_0007_),
    .Q(\input_buffer[2][11] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][12]$_DFFE_PP_  (.D(net108),
    .DE(_0007_),
    .Q(\input_buffer[2][12] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][13]$_DFFE_PP_  (.D(net109),
    .DE(_0007_),
    .Q(\input_buffer[2][13] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][14]$_DFFE_PP_  (.D(net110),
    .DE(_0007_),
    .Q(\input_buffer[2][14] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][15]$_DFFE_PP_  (.D(net111),
    .DE(_0007_),
    .Q(\input_buffer[2][15] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][16]$_DFFE_PP_  (.D(net112),
    .DE(_0007_),
    .Q(\input_buffer[2][16] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][17]$_DFFE_PP_  (.D(net113),
    .DE(_0007_),
    .Q(\input_buffer[2][17] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][18]$_DFFE_PP_  (.D(net114),
    .DE(_0007_),
    .Q(\input_buffer[2][18] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][19]$_DFFE_PP_  (.D(net115),
    .DE(_0007_),
    .Q(\input_buffer[2][19] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][1]$_DFFE_PP_  (.D(net116),
    .DE(_0007_),
    .Q(\input_buffer[2][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][20]$_DFFE_PP_  (.D(net117),
    .DE(_0007_),
    .Q(\input_buffer[2][20] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][21]$_DFFE_PP_  (.D(net118),
    .DE(_0007_),
    .Q(\input_buffer[2][21] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][22]$_DFFE_PP_  (.D(net119),
    .DE(_0007_),
    .Q(\input_buffer[2][22] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][23]$_DFFE_PP_  (.D(net120),
    .DE(_0007_),
    .Q(\input_buffer[2][23] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][24]$_DFFE_PP_  (.D(net121),
    .DE(_0007_),
    .Q(\dest_id[2][0] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][25]$_DFFE_PP_  (.D(net122),
    .DE(_0007_),
    .Q(\dest_id[2][1] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][26]$_DFFE_PP_  (.D(net123),
    .DE(_0007_),
    .Q(\dest_id[2][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][27]$_DFFE_PP_  (.D(net124),
    .DE(_0007_),
    .Q(\dest_id[2][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][28]$_DFFE_PP_  (.D(net125),
    .DE(_0007_),
    .Q(\dest_id[2][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][29]$_DFFE_PP_  (.D(net126),
    .DE(_0007_),
    .Q(\dest_id[2][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][2]$_DFFE_PP_  (.D(net127),
    .DE(_0007_),
    .Q(\input_buffer[2][2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][30]$_DFFE_PP_  (.D(net128),
    .DE(_0007_),
    .Q(\dest_id[2][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][31]$_DFFE_PP_  (.D(net129),
    .DE(_0007_),
    .Q(\dest_id[2][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][3]$_DFFE_PP_  (.D(net130),
    .DE(_0007_),
    .Q(\input_buffer[2][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][4]$_DFFE_PP_  (.D(net131),
    .DE(_0007_),
    .Q(\input_buffer[2][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][5]$_DFFE_PP_  (.D(net132),
    .DE(_0007_),
    .Q(\input_buffer[2][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][6]$_DFFE_PP_  (.D(net133),
    .DE(_0007_),
    .Q(\input_buffer[2][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][7]$_DFFE_PP_  (.D(net134),
    .DE(_0007_),
    .Q(\input_buffer[2][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][8]$_DFFE_PP_  (.D(net135),
    .DE(_0007_),
    .Q(\input_buffer[2][8] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[2][9]$_DFFE_PP_  (.D(net136),
    .DE(_0007_),
    .Q(\input_buffer[2][9] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][0]$_DFFE_PP_  (.D(net139),
    .DE(_0006_),
    .Q(\input_buffer[3][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][10]$_DFFE_PP_  (.D(net140),
    .DE(_0006_),
    .Q(\input_buffer[3][10] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][11]$_DFFE_PP_  (.D(net141),
    .DE(_0006_),
    .Q(\input_buffer[3][11] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][12]$_DFFE_PP_  (.D(net142),
    .DE(_0006_),
    .Q(\input_buffer[3][12] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][13]$_DFFE_PP_  (.D(net143),
    .DE(_0006_),
    .Q(\input_buffer[3][13] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][14]$_DFFE_PP_  (.D(net144),
    .DE(_0006_),
    .Q(\input_buffer[3][14] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][15]$_DFFE_PP_  (.D(net145),
    .DE(_0006_),
    .Q(\input_buffer[3][15] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][16]$_DFFE_PP_  (.D(net146),
    .DE(_0006_),
    .Q(\input_buffer[3][16] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][17]$_DFFE_PP_  (.D(net147),
    .DE(_0006_),
    .Q(\input_buffer[3][17] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][18]$_DFFE_PP_  (.D(net148),
    .DE(_0006_),
    .Q(\input_buffer[3][18] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][19]$_DFFE_PP_  (.D(net149),
    .DE(_0006_),
    .Q(\input_buffer[3][19] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][1]$_DFFE_PP_  (.D(net150),
    .DE(_0006_),
    .Q(\input_buffer[3][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][20]$_DFFE_PP_  (.D(net151),
    .DE(_0006_),
    .Q(\input_buffer[3][20] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][21]$_DFFE_PP_  (.D(net152),
    .DE(_0006_),
    .Q(\input_buffer[3][21] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][22]$_DFFE_PP_  (.D(net153),
    .DE(_0006_),
    .Q(\input_buffer[3][22] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][23]$_DFFE_PP_  (.D(net154),
    .DE(_0006_),
    .Q(\input_buffer[3][23] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][24]$_DFFE_PP_  (.D(net155),
    .DE(_0006_),
    .Q(\dest_id[3][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][25]$_DFFE_PP_  (.D(net156),
    .DE(_0006_),
    .Q(\dest_id[3][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][26]$_DFFE_PP_  (.D(net157),
    .DE(_0006_),
    .Q(\dest_id[3][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][27]$_DFFE_PP_  (.D(net158),
    .DE(_0006_),
    .Q(\dest_id[3][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][28]$_DFFE_PP_  (.D(net159),
    .DE(_0006_),
    .Q(\dest_id[3][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][29]$_DFFE_PP_  (.D(net160),
    .DE(_0006_),
    .Q(\dest_id[3][5] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][2]$_DFFE_PP_  (.D(net161),
    .DE(_0006_),
    .Q(\input_buffer[3][2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][30]$_DFFE_PP_  (.D(net162),
    .DE(_0006_),
    .Q(\dest_id[3][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][31]$_DFFE_PP_  (.D(net163),
    .DE(_0006_),
    .Q(\dest_id[3][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][3]$_DFFE_PP_  (.D(net164),
    .DE(_0006_),
    .Q(\input_buffer[3][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][4]$_DFFE_PP_  (.D(net165),
    .DE(_0006_),
    .Q(\input_buffer[3][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][5]$_DFFE_PP_  (.D(net166),
    .DE(_0006_),
    .Q(\input_buffer[3][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][6]$_DFFE_PP_  (.D(net167),
    .DE(_0006_),
    .Q(\input_buffer[3][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][7]$_DFFE_PP_  (.D(net168),
    .DE(_0006_),
    .Q(\input_buffer[3][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][8]$_DFFE_PP_  (.D(net169),
    .DE(_0006_),
    .Q(\input_buffer[3][8] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[3][9]$_DFFE_PP_  (.D(net170),
    .DE(_0006_),
    .Q(\input_buffer[3][9] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][0]$_DFFE_PP_  (.D(net36),
    .DE(_0005_),
    .Q(\input_buffer[4][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][10]$_DFFE_PP_  (.D(net37),
    .DE(_0005_),
    .Q(\input_buffer[4][10] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][11]$_DFFE_PP_  (.D(net38),
    .DE(_0005_),
    .Q(\input_buffer[4][11] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][12]$_DFFE_PP_  (.D(net39),
    .DE(_0005_),
    .Q(\input_buffer[4][12] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][13]$_DFFE_PP_  (.D(net40),
    .DE(_0005_),
    .Q(\input_buffer[4][13] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][14]$_DFFE_PP_  (.D(net41),
    .DE(_0005_),
    .Q(\input_buffer[4][14] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][15]$_DFFE_PP_  (.D(net42),
    .DE(_0005_),
    .Q(\input_buffer[4][15] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][16]$_DFFE_PP_  (.D(net43),
    .DE(_0005_),
    .Q(\input_buffer[4][16] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][17]$_DFFE_PP_  (.D(net44),
    .DE(_0005_),
    .Q(\input_buffer[4][17] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][18]$_DFFE_PP_  (.D(net45),
    .DE(_0005_),
    .Q(\input_buffer[4][18] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][19]$_DFFE_PP_  (.D(net46),
    .DE(_0005_),
    .Q(\input_buffer[4][19] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][1]$_DFFE_PP_  (.D(net47),
    .DE(_0005_),
    .Q(\input_buffer[4][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][20]$_DFFE_PP_  (.D(net48),
    .DE(_0005_),
    .Q(\input_buffer[4][20] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][21]$_DFFE_PP_  (.D(net49),
    .DE(_0005_),
    .Q(\input_buffer[4][21] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][22]$_DFFE_PP_  (.D(net50),
    .DE(_0005_),
    .Q(\input_buffer[4][22] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][23]$_DFFE_PP_  (.D(net51),
    .DE(_0005_),
    .Q(\input_buffer[4][23] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][24]$_DFFE_PP_  (.D(net52),
    .DE(_0005_),
    .Q(\dest_id[4][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][25]$_DFFE_PP_  (.D(net53),
    .DE(_0005_),
    .Q(\dest_id[4][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][26]$_DFFE_PP_  (.D(net54),
    .DE(_0005_),
    .Q(\dest_id[4][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][27]$_DFFE_PP_  (.D(net55),
    .DE(_0005_),
    .Q(\dest_id[4][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][28]$_DFFE_PP_  (.D(net56),
    .DE(_0005_),
    .Q(\dest_id[4][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][29]$_DFFE_PP_  (.D(net57),
    .DE(_0005_),
    .Q(\dest_id[4][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][2]$_DFFE_PP_  (.D(net58),
    .DE(_0005_),
    .Q(\input_buffer[4][2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][30]$_DFFE_PP_  (.D(net59),
    .DE(_0005_),
    .Q(\dest_id[4][6] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][31]$_DFFE_PP_  (.D(net60),
    .DE(_0005_),
    .Q(\dest_id[4][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][3]$_DFFE_PP_  (.D(net61),
    .DE(_0005_),
    .Q(\input_buffer[4][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][4]$_DFFE_PP_  (.D(net62),
    .DE(_0005_),
    .Q(\input_buffer[4][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][5]$_DFFE_PP_  (.D(net63),
    .DE(_0005_),
    .Q(\input_buffer[4][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][6]$_DFFE_PP_  (.D(net64),
    .DE(_0005_),
    .Q(\input_buffer[4][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][7]$_DFFE_PP_  (.D(net65),
    .DE(_0005_),
    .Q(\input_buffer[4][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][8]$_DFFE_PP_  (.D(net66),
    .DE(_0005_),
    .Q(\input_buffer[4][8] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \input_buffer[4][9]$_DFFE_PP_  (.D(net67),
    .DE(_0005_),
    .Q(\input_buffer[4][9] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \input_buffer_valid[0]$_DFF_PN0_  (.D(_0000_),
    .Q(\input_buffer_valid[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \input_buffer_valid[1]$_DFF_PN0_  (.D(_0001_),
    .Q(\input_buffer_valid[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \input_buffer_valid[2]$_DFF_PN0_  (.D(_0002_),
    .Q(\input_buffer_valid[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \input_buffer_valid[3]$_DFF_PN0_  (.D(_0003_),
    .Q(\input_buffer_valid[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \input_buffer_valid[4]$_DFF_PN0_  (.D(_0004_),
    .Q(\input_buffer_valid[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_2 hold1 (.A(net104),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_312 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(net498),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net447),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net436),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net480),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net457),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net390),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net460),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net452),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net499),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net411),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net376),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(net364),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net348),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(net362),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(net379),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net425),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(net495),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(net409),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(net492),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(net497),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(net488),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(net465),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net408),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(net469),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(net477),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(net496),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net357),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(net372),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(net352),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net360),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(net481),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(net471),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(east_in_valid),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(east_out_ready),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(net484),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(net433),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(net479),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(net444),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(net458),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(net467),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(net403),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(net478),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net427),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(net483),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net374),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(net472),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net356),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(net387),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(net449),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(net487),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(net416),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(net437),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(net490),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net442),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(net422),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(net429),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(net424),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(net365),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(net464),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(local_in_data[3]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(net371),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(net383),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(net388),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net386),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(local_in_data[8]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(local_in_data[9]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(local_in_valid),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input68 (.A(local_out_ready),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(net414),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(net399),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(net441),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(net406),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(net400),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(net396),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(net382),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(net404),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(net373),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(net369),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(net451),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(net461),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(net401),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(net491),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(net349),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(net350),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(net381),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(net454),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(net380),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(net430),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(net459),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(net440),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(net468),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(net466),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(net412),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(net358),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(net361),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(net410),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(net394),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(net476),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(net415),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(net393),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(north_in_valid),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(north_out_ready),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input103 (.A(net343),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(south_in_data[0]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(net475),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(net405),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(net485),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(net482),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(net426),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(net368),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(net397),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(net474),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(net423),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(net377),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(net363),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(net351),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(net417),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(net398),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(net392),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(net413),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(net494),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(net431),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(net375),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(net378),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(net402),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(net391),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(net446),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(net455),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(net359),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(net346),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(net347),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(net367),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(net443),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(net407),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(net420),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(south_in_valid),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(south_out_ready),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(net470),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(net428),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(net370),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(net453),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(net456),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(net463),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(net438),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(net473),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(net462),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(net486),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(net366),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(net448),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(net353),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(net344),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(net345),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(net432),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(net489),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(net419),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(net439),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(net435),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(net395),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(net450),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(net389),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(net418),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(net421),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(net385),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(net384),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(net354),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(net434),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(net355),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(net445),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(net493),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(west_in_valid),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input171 (.A(west_out_ready),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net173),
    .X(east_in_ready));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net174),
    .X(east_out_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net175),
    .X(east_out_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net176),
    .X(east_out_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net177),
    .X(east_out_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net178),
    .X(east_out_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net179),
    .X(east_out_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net180),
    .X(east_out_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net181),
    .X(east_out_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net182),
    .X(east_out_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net183),
    .X(east_out_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net184),
    .X(east_out_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net185),
    .X(east_out_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net186),
    .X(east_out_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net187),
    .X(east_out_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net188),
    .X(east_out_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net189),
    .X(east_out_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net190),
    .X(east_out_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net191),
    .X(east_out_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net192),
    .X(east_out_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net193),
    .X(east_out_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net194),
    .X(east_out_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net195),
    .X(east_out_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net196),
    .X(east_out_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net197),
    .X(east_out_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net198),
    .X(east_out_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net199),
    .X(east_out_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net200),
    .X(east_out_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net201),
    .X(east_out_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net202),
    .X(east_out_valid));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net203),
    .X(local_in_ready));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net204),
    .X(local_out_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net205),
    .X(local_out_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net206),
    .X(local_out_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net207),
    .X(local_out_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net208),
    .X(local_out_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net209),
    .X(local_out_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net210),
    .X(local_out_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net211),
    .X(local_out_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net212),
    .X(local_out_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net213),
    .X(local_out_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net214),
    .X(local_out_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net215),
    .X(local_out_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net216),
    .X(local_out_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net217),
    .X(local_out_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net218),
    .X(local_out_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net219),
    .X(local_out_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net220),
    .X(local_out_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output220 (.A(net221),
    .X(local_out_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net222),
    .X(local_out_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net223),
    .X(local_out_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output223 (.A(net224),
    .X(local_out_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net225),
    .X(local_out_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output225 (.A(net226),
    .X(local_out_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net227),
    .X(local_out_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output227 (.A(net228),
    .X(local_out_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output228 (.A(net229),
    .X(local_out_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net230),
    .X(local_out_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net231),
    .X(local_out_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output231 (.A(net232),
    .X(local_out_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output232 (.A(net233),
    .X(local_out_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net234),
    .X(local_out_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output234 (.A(net235),
    .X(local_out_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(net236),
    .X(local_out_valid));
 sky130_fd_sc_hd__clkbuf_1 output236 (.A(net237),
    .X(north_in_ready));
 sky130_fd_sc_hd__clkbuf_1 output237 (.A(net238),
    .X(north_out_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net239),
    .X(north_out_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output239 (.A(net240),
    .X(north_out_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output240 (.A(net241),
    .X(north_out_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net242),
    .X(north_out_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net243),
    .X(north_out_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output243 (.A(net244),
    .X(north_out_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output244 (.A(net245),
    .X(north_out_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net246),
    .X(north_out_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output246 (.A(net247),
    .X(north_out_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net248),
    .X(north_out_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output248 (.A(net249),
    .X(north_out_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output249 (.A(net250),
    .X(north_out_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output250 (.A(net251),
    .X(north_out_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output251 (.A(net252),
    .X(north_out_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output252 (.A(net253),
    .X(north_out_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output253 (.A(net254),
    .X(north_out_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output254 (.A(net255),
    .X(north_out_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output255 (.A(net256),
    .X(north_out_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output256 (.A(net257),
    .X(north_out_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output257 (.A(net258),
    .X(north_out_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output258 (.A(net259),
    .X(north_out_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output259 (.A(net260),
    .X(north_out_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output260 (.A(net261),
    .X(north_out_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output261 (.A(net262),
    .X(north_out_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output262 (.A(net263),
    .X(north_out_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output263 (.A(net264),
    .X(north_out_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output264 (.A(net265),
    .X(north_out_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output265 (.A(net266),
    .X(north_out_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output266 (.A(net267),
    .X(north_out_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output267 (.A(net268),
    .X(north_out_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output268 (.A(net269),
    .X(north_out_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output269 (.A(net270),
    .X(north_out_valid));
 sky130_fd_sc_hd__clkbuf_1 output270 (.A(net271),
    .X(south_in_ready));
 sky130_fd_sc_hd__clkbuf_1 output271 (.A(net272),
    .X(south_out_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output272 (.A(net273),
    .X(south_out_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output273 (.A(net274),
    .X(south_out_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output274 (.A(net275),
    .X(south_out_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output275 (.A(net276),
    .X(south_out_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output276 (.A(net277),
    .X(south_out_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output277 (.A(net278),
    .X(south_out_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output278 (.A(net279),
    .X(south_out_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output279 (.A(net280),
    .X(south_out_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output280 (.A(net281),
    .X(south_out_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output281 (.A(net282),
    .X(south_out_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output282 (.A(net283),
    .X(south_out_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output283 (.A(net284),
    .X(south_out_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output284 (.A(net285),
    .X(south_out_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output285 (.A(net286),
    .X(south_out_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output286 (.A(net287),
    .X(south_out_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output287 (.A(net288),
    .X(south_out_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output288 (.A(net289),
    .X(south_out_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output289 (.A(net290),
    .X(south_out_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output290 (.A(net291),
    .X(south_out_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output291 (.A(net292),
    .X(south_out_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output292 (.A(net293),
    .X(south_out_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output293 (.A(net294),
    .X(south_out_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output294 (.A(net295),
    .X(south_out_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output295 (.A(net296),
    .X(south_out_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output296 (.A(net297),
    .X(south_out_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output297 (.A(net298),
    .X(south_out_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output298 (.A(net299),
    .X(south_out_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output299 (.A(net300),
    .X(south_out_valid));
 sky130_fd_sc_hd__clkbuf_1 output300 (.A(net301),
    .X(west_in_ready));
 sky130_fd_sc_hd__clkbuf_1 output301 (.A(net302),
    .X(west_out_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output302 (.A(net303),
    .X(west_out_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output303 (.A(net304),
    .X(west_out_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output304 (.A(net305),
    .X(west_out_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output305 (.A(net306),
    .X(west_out_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output306 (.A(net307),
    .X(west_out_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output307 (.A(net308),
    .X(west_out_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output308 (.A(net309),
    .X(west_out_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output309 (.A(net310),
    .X(west_out_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output310 (.A(net311),
    .X(west_out_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output311 (.A(net312),
    .X(west_out_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output312 (.A(net313),
    .X(west_out_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output313 (.A(net314),
    .X(west_out_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output314 (.A(net315),
    .X(west_out_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output315 (.A(net316),
    .X(west_out_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output316 (.A(net317),
    .X(west_out_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output317 (.A(net318),
    .X(west_out_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output318 (.A(net319),
    .X(west_out_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output319 (.A(net320),
    .X(west_out_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output320 (.A(net321),
    .X(west_out_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output321 (.A(net322),
    .X(west_out_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output322 (.A(net323),
    .X(west_out_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output323 (.A(net324),
    .X(west_out_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output324 (.A(net325),
    .X(west_out_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output325 (.A(net326),
    .X(west_out_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output326 (.A(net327),
    .X(west_out_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output327 (.A(net328),
    .X(west_out_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output328 (.A(net329),
    .X(west_out_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output329 (.A(net330),
    .X(west_out_valid));
 sky130_fd_sc_hd__conb_1 _2459__330 (.LO(net331));
 sky130_fd_sc_hd__conb_1 _2460__331 (.LO(net332));
 sky130_fd_sc_hd__conb_1 _2461__332 (.LO(net333));
 sky130_fd_sc_hd__conb_1 _2462__333 (.LO(net334));
 sky130_fd_sc_hd__conb_1 _2463__334 (.LO(net335));
 sky130_fd_sc_hd__conb_1 _2464__335 (.LO(net336));
 sky130_fd_sc_hd__conb_1 _2465__336 (.LO(net337));
 sky130_fd_sc_hd__conb_1 _2466__337 (.LO(net338));
 sky130_fd_sc_hd__conb_1 _2467__338 (.LO(net339));
 sky130_fd_sc_hd__conb_1 _2468__339 (.LO(net340));
 sky130_fd_sc_hd__conb_1 _2469__340 (.LO(net341));
 sky130_fd_sc_hd__conb_1 _2470__341 (.LO(net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_8 clkload1 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload6 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload7 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload8 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload10 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_8 clkload12 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload13 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(west_in_data[21]),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(west_in_data[22]),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(south_in_data[4]),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(south_in_data[5]),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(east_in_data[20]),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(north_in_data[22]),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(north_in_data[23]),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(south_in_data[20]),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(east_in_data[6]),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(west_in_data[20]),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(west_in_data[5]),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(west_in_data[7]),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(local_in_data[20]),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(east_in_data[4]),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(north_in_data[3]),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(south_in_data[3]),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(east_in_data[7]),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(north_in_data[4]),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(east_in_data[21]),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(south_in_data[1]),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(east_in_data[1]),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(local_in_data[30]),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(west_in_data[19]),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(south_in_data[6]),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(south_in_data[15]),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(north_in_data[18]),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(west_in_data[11]),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(local_in_data[4]),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(east_in_data[5]),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(north_in_data[17]),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(local_in_data[19]),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(south_in_data[27]),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(east_in_data[19]),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(south_in_data[19]),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(south_in_data[28]),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(east_in_data[22]),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(north_in_data[26]),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(north_in_data[24]),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(north_in_data[15]),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(local_in_data[5]),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(west_in_data[4]),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(west_in_data[3]),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(local_in_data[7]),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(local_in_data[21]),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(local_in_data[6]),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(west_in_data[2]),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(east_in_data[14]),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(south_in_data[2]),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(south_in_data[23]),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(north_in_data[9]),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(north_in_data[6]),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(west_in_data[28]),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(north_in_data[14]),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(south_in_data[16]),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(south_in_data[22]),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(north_in_data[10]),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(north_in_data[13]),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(north_in_data[20]),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(south_in_data[29]),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(local_in_data[15]),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(north_in_data[16]),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(south_in_data[11]),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(north_in_data[12]),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(south_in_data[8]),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(east_in_data[2]),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(east_in_data[25]),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(north_in_data[5]),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(east_in_data[18]),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(north_in_data[31]),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(south_in_data[24]),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(north_in_data[0]),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(north_in_data[8]),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(local_in_data[24]),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(south_in_data[21]),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(west_in_data[30]),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(west_in_data[25]),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(south_in_data[9]),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(west_in_data[31]),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(local_in_data[28]),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(south_in_data[18]),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(local_in_data[2]),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(east_in_data[23]),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(south_in_data[14]),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(local_in_data[17]),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(west_in_data[10]),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(local_in_data[29]),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(north_in_data[27]),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(south_in_data[26]),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(west_in_data[23]),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(local_in_data[10]),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(west_in_data[6]),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(west_in_data[27]),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(east_in_data[11]),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(local_in_data[25]),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(west_in_data[15]),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(west_in_data[26]),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(north_in_data[29]),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(north_in_data[11]),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(local_in_data[27]),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(south_in_data[7]),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(local_in_data[12]),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(west_in_data[8]),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(south_in_data[30]),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(east_in_data[10]),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(west_in_data[1]),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(local_in_data[22]),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(west_in_data[29]),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(north_in_data[19]),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(east_in_data[16]),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(west_in_data[12]),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(north_in_data[25]),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(south_in_data[31]),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(west_in_data[13]),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(east_in_data[13]),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(local_in_data[13]),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(north_in_data[28]),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(east_in_data[15]),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(north_in_data[1]),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(west_in_data[17]),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(west_in_data[14]),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(local_in_data[31]),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(east_in_data[29]),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(north_in_data[30]),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(local_in_data[14]),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(north_in_data[2]),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(east_in_data[30]),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(west_in_data[0]),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(east_in_data[9]),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(local_in_data[1]),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(west_in_data[16]),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(south_in_data[17]),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(south_in_data[10]),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(north_in_data[7]),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(east_in_data[31]),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(local_in_data[16]),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(local_in_data[11]),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(east_in_data[12]),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(east_in_data[8]),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(south_in_data[13]),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(local_in_data[18]),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(local_in_data[0]),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(south_in_data[12]),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(west_in_data[18]),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(local_in_data[23]),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(east_in_data[28]),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(west_in_data[24]),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(local_in_data[26]),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(north_in_data[21]),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(east_in_data[26]),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(west_in_data[9]),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(south_in_data[25]),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(east_in_data[24]),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(east_in_data[3]),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(east_in_data[27]),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(east_in_data[0]),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(east_in_data[17]),
    .X(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0344_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_328 ();
endmodule
