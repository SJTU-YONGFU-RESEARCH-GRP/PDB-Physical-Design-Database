module jtag_controller (clk,
    dr_shift_en,
    rst_n,
    tck,
    tdi,
    tdo,
    tms,
    trst_n,
    update_dr,
    dr_in,
    dr_out,
    instruction);
 input clk;
 output dr_shift_en;
 input rst_n;
 input tck;
 input tdi;
 output tdo;
 input tms;
 input trst_n;
 output update_dr;
 input [31:0] dr_in;
 output [31:0] dr_out;
 output [4:0] instruction;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire \dr_shift_reg[0] ;
 wire \dr_shift_reg[10] ;
 wire \dr_shift_reg[11] ;
 wire \dr_shift_reg[12] ;
 wire \dr_shift_reg[13] ;
 wire \dr_shift_reg[14] ;
 wire \dr_shift_reg[15] ;
 wire \dr_shift_reg[16] ;
 wire \dr_shift_reg[17] ;
 wire \dr_shift_reg[18] ;
 wire \dr_shift_reg[19] ;
 wire \dr_shift_reg[1] ;
 wire \dr_shift_reg[20] ;
 wire \dr_shift_reg[21] ;
 wire \dr_shift_reg[22] ;
 wire \dr_shift_reg[23] ;
 wire \dr_shift_reg[24] ;
 wire \dr_shift_reg[25] ;
 wire \dr_shift_reg[26] ;
 wire \dr_shift_reg[27] ;
 wire \dr_shift_reg[28] ;
 wire \dr_shift_reg[29] ;
 wire \dr_shift_reg[2] ;
 wire \dr_shift_reg[30] ;
 wire \dr_shift_reg[31] ;
 wire \dr_shift_reg[3] ;
 wire \dr_shift_reg[4] ;
 wire \dr_shift_reg[5] ;
 wire \dr_shift_reg[6] ;
 wire \dr_shift_reg[7] ;
 wire \dr_shift_reg[8] ;
 wire \dr_shift_reg[9] ;
 wire \ir_shift_reg[0] ;
 wire \ir_shift_reg[1] ;
 wire \ir_shift_reg[2] ;
 wire \ir_shift_reg[3] ;
 wire \ir_shift_reg[4] ;
 wire \next_tap_state[0] ;
 wire \next_tap_state[1] ;
 wire \next_tap_state[2] ;
 wire \next_tap_state[3] ;
 wire \tap_state[0] ;
 wire \tap_state[1] ;
 wire \tap_state[2] ;
 wire \tap_state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;

 BUF_X4 _247_ (.A(\tap_state[3] ),
    .Z(_076_));
 INV_X2 _248_ (.A(_076_),
    .ZN(_077_));
 BUF_X4 _249_ (.A(\tap_state[0] ),
    .Z(_078_));
 NOR2_X2 _250_ (.A1(\tap_state[1] ),
    .A2(_078_),
    .ZN(_079_));
 NAND3_X2 _251_ (.A1(_077_),
    .A2(\tap_state[2] ),
    .A3(_079_),
    .ZN(_080_));
 INV_X2 _252_ (.A(_080_),
    .ZN(net68));
 INV_X1 _253_ (.A(\dr_shift_reg[0] ),
    .ZN(_081_));
 BUF_X4 _254_ (.A(\tap_state[1] ),
    .Z(_082_));
 NAND2_X1 _255_ (.A1(_082_),
    .A2(_078_),
    .ZN(_083_));
 BUF_X4 _256_ (.A(\tap_state[2] ),
    .Z(_084_));
 NOR2_X2 _257_ (.A1(_077_),
    .A2(_084_),
    .ZN(_085_));
 NAND2_X1 _258_ (.A1(\ir_shift_reg[0] ),
    .A2(_085_),
    .ZN(_086_));
 OAI22_X1 _259_ (.A1(_081_),
    .A2(_080_),
    .B1(_083_),
    .B2(_086_),
    .ZN(_000_));
 NAND2_X4 _260_ (.A1(_079_),
    .A2(_085_),
    .ZN(_087_));
 BUF_X4 _261_ (.A(_087_),
    .Z(_088_));
 INV_X1 _262_ (.A(_088_),
    .ZN(net75));
 INV_X8 _263_ (.A(net33),
    .ZN(_001_));
 MUX2_X1 _264_ (.A(\dr_shift_reg[17] ),
    .B(net44),
    .S(_088_),
    .Z(_002_));
 MUX2_X1 _265_ (.A(\dr_shift_reg[18] ),
    .B(net45),
    .S(_088_),
    .Z(_003_));
 MUX2_X1 _266_ (.A(\dr_shift_reg[19] ),
    .B(net46),
    .S(_088_),
    .Z(_004_));
 MUX2_X1 _267_ (.A(\dr_shift_reg[1] ),
    .B(net47),
    .S(_088_),
    .Z(_005_));
 MUX2_X1 _268_ (.A(\dr_shift_reg[20] ),
    .B(net48),
    .S(_088_),
    .Z(_006_));
 MUX2_X1 _269_ (.A(\dr_shift_reg[21] ),
    .B(net49),
    .S(_088_),
    .Z(_007_));
 MUX2_X1 _270_ (.A(\dr_shift_reg[22] ),
    .B(net50),
    .S(_088_),
    .Z(_008_));
 MUX2_X1 _271_ (.A(\dr_shift_reg[23] ),
    .B(net51),
    .S(_088_),
    .Z(_009_));
 MUX2_X1 _272_ (.A(\dr_shift_reg[24] ),
    .B(net52),
    .S(_088_),
    .Z(_010_));
 BUF_X4 _273_ (.A(_087_),
    .Z(_089_));
 MUX2_X1 _274_ (.A(\dr_shift_reg[25] ),
    .B(net53),
    .S(_089_),
    .Z(_011_));
 MUX2_X1 _275_ (.A(\dr_shift_reg[26] ),
    .B(net54),
    .S(_089_),
    .Z(_012_));
 MUX2_X1 _276_ (.A(\dr_shift_reg[27] ),
    .B(net55),
    .S(_089_),
    .Z(_013_));
 MUX2_X1 _277_ (.A(\dr_shift_reg[28] ),
    .B(net56),
    .S(_089_),
    .Z(_014_));
 MUX2_X1 _278_ (.A(\dr_shift_reg[29] ),
    .B(net57),
    .S(_089_),
    .Z(_015_));
 MUX2_X1 _279_ (.A(\dr_shift_reg[2] ),
    .B(net58),
    .S(_089_),
    .Z(_016_));
 MUX2_X1 _280_ (.A(\dr_shift_reg[30] ),
    .B(net59),
    .S(_089_),
    .Z(_017_));
 MUX2_X1 _281_ (.A(\dr_shift_reg[31] ),
    .B(net60),
    .S(_089_),
    .Z(_018_));
 MUX2_X1 _282_ (.A(\dr_shift_reg[3] ),
    .B(net61),
    .S(_089_),
    .Z(_019_));
 MUX2_X1 _283_ (.A(\dr_shift_reg[4] ),
    .B(net62),
    .S(_089_),
    .Z(_020_));
 BUF_X4 _284_ (.A(_087_),
    .Z(_090_));
 MUX2_X1 _285_ (.A(\dr_shift_reg[5] ),
    .B(net63),
    .S(_090_),
    .Z(_021_));
 MUX2_X1 _286_ (.A(\dr_shift_reg[6] ),
    .B(net64),
    .S(_090_),
    .Z(_022_));
 MUX2_X1 _287_ (.A(\dr_shift_reg[7] ),
    .B(net65),
    .S(_090_),
    .Z(_023_));
 MUX2_X1 _288_ (.A(\dr_shift_reg[8] ),
    .B(net66),
    .S(_090_),
    .Z(_024_));
 MUX2_X1 _289_ (.A(\dr_shift_reg[9] ),
    .B(net67),
    .S(_090_),
    .Z(_025_));
 NAND2_X1 _290_ (.A1(\dr_shift_reg[1] ),
    .A2(net68),
    .ZN(_091_));
 NOR2_X2 _291_ (.A1(_076_),
    .A2(\tap_state[2] ),
    .ZN(_092_));
 NAND3_X4 _292_ (.A1(_082_),
    .A2(_078_),
    .A3(_092_),
    .ZN(_093_));
 NAND2_X4 _293_ (.A1(_080_),
    .A2(_093_),
    .ZN(_094_));
 BUF_X8 _294_ (.A(_094_),
    .Z(_095_));
 INV_X1 _295_ (.A(net1),
    .ZN(_096_));
 BUF_X4 _296_ (.A(_093_),
    .Z(_097_));
 OAI221_X1 _297_ (.A(_091_),
    .B1(_095_),
    .B2(_081_),
    .C1(_096_),
    .C2(_097_),
    .ZN(_026_));
 NAND2_X1 _298_ (.A1(\dr_shift_reg[11] ),
    .A2(net68),
    .ZN(_098_));
 INV_X1 _299_ (.A(net2),
    .ZN(_099_));
 INV_X1 _300_ (.A(\dr_shift_reg[10] ),
    .ZN(_100_));
 OAI221_X1 _301_ (.A(_098_),
    .B1(_097_),
    .B2(_099_),
    .C1(_100_),
    .C2(_095_),
    .ZN(_027_));
 MUX2_X1 _302_ (.A(net3),
    .B(\dr_shift_reg[12] ),
    .S(_097_),
    .Z(_101_));
 MUX2_X1 _303_ (.A(\dr_shift_reg[11] ),
    .B(_101_),
    .S(_095_),
    .Z(_028_));
 MUX2_X1 _304_ (.A(net4),
    .B(\dr_shift_reg[13] ),
    .S(_097_),
    .Z(_102_));
 MUX2_X1 _305_ (.A(\dr_shift_reg[12] ),
    .B(_102_),
    .S(_095_),
    .Z(_029_));
 MUX2_X1 _306_ (.A(net5),
    .B(\dr_shift_reg[14] ),
    .S(_097_),
    .Z(_103_));
 MUX2_X1 _307_ (.A(\dr_shift_reg[13] ),
    .B(_103_),
    .S(_095_),
    .Z(_030_));
 MUX2_X1 _308_ (.A(\dr_shift_reg[14] ),
    .B(\dr_shift_reg[15] ),
    .S(net68),
    .Z(_104_));
 MUX2_X1 _309_ (.A(net6),
    .B(_104_),
    .S(_097_),
    .Z(_031_));
 MUX2_X1 _310_ (.A(net7),
    .B(\dr_shift_reg[16] ),
    .S(_097_),
    .Z(_105_));
 MUX2_X1 _311_ (.A(\dr_shift_reg[15] ),
    .B(_105_),
    .S(_095_),
    .Z(_032_));
 MUX2_X1 _312_ (.A(net8),
    .B(\dr_shift_reg[17] ),
    .S(_097_),
    .Z(_106_));
 MUX2_X1 _313_ (.A(\dr_shift_reg[16] ),
    .B(_106_),
    .S(_095_),
    .Z(_033_));
 MUX2_X1 _314_ (.A(net9),
    .B(\dr_shift_reg[18] ),
    .S(_097_),
    .Z(_107_));
 MUX2_X1 _315_ (.A(\dr_shift_reg[17] ),
    .B(_107_),
    .S(_095_),
    .Z(_034_));
 BUF_X8 _316_ (.A(_093_),
    .Z(_108_));
 MUX2_X1 _317_ (.A(net10),
    .B(\dr_shift_reg[19] ),
    .S(_108_),
    .Z(_109_));
 MUX2_X1 _318_ (.A(\dr_shift_reg[18] ),
    .B(_109_),
    .S(_095_),
    .Z(_035_));
 MUX2_X1 _319_ (.A(net11),
    .B(\dr_shift_reg[20] ),
    .S(_108_),
    .Z(_110_));
 MUX2_X1 _320_ (.A(\dr_shift_reg[19] ),
    .B(_110_),
    .S(_095_),
    .Z(_036_));
 MUX2_X1 _321_ (.A(net12),
    .B(\dr_shift_reg[2] ),
    .S(_108_),
    .Z(_111_));
 BUF_X8 _322_ (.A(_094_),
    .Z(_112_));
 MUX2_X1 _323_ (.A(\dr_shift_reg[1] ),
    .B(_111_),
    .S(_112_),
    .Z(_037_));
 MUX2_X1 _324_ (.A(net13),
    .B(\dr_shift_reg[21] ),
    .S(_108_),
    .Z(_113_));
 MUX2_X1 _325_ (.A(\dr_shift_reg[20] ),
    .B(_113_),
    .S(_112_),
    .Z(_038_));
 MUX2_X1 _326_ (.A(net14),
    .B(\dr_shift_reg[22] ),
    .S(_108_),
    .Z(_114_));
 MUX2_X1 _327_ (.A(\dr_shift_reg[21] ),
    .B(_114_),
    .S(_112_),
    .Z(_039_));
 MUX2_X1 _328_ (.A(net15),
    .B(\dr_shift_reg[23] ),
    .S(_108_),
    .Z(_115_));
 MUX2_X1 _329_ (.A(\dr_shift_reg[22] ),
    .B(_115_),
    .S(_112_),
    .Z(_040_));
 MUX2_X1 _330_ (.A(net16),
    .B(\dr_shift_reg[24] ),
    .S(_108_),
    .Z(_116_));
 MUX2_X1 _331_ (.A(\dr_shift_reg[23] ),
    .B(_116_),
    .S(_112_),
    .Z(_041_));
 MUX2_X1 _332_ (.A(net17),
    .B(\dr_shift_reg[25] ),
    .S(_108_),
    .Z(_117_));
 MUX2_X1 _333_ (.A(\dr_shift_reg[24] ),
    .B(_117_),
    .S(_112_),
    .Z(_042_));
 MUX2_X1 _334_ (.A(net18),
    .B(\dr_shift_reg[26] ),
    .S(_108_),
    .Z(_118_));
 MUX2_X1 _335_ (.A(\dr_shift_reg[25] ),
    .B(_118_),
    .S(_112_),
    .Z(_043_));
 MUX2_X1 _336_ (.A(net19),
    .B(\dr_shift_reg[27] ),
    .S(_108_),
    .Z(_119_));
 MUX2_X1 _337_ (.A(\dr_shift_reg[26] ),
    .B(_119_),
    .S(_112_),
    .Z(_044_));
 BUF_X4 _338_ (.A(_093_),
    .Z(_120_));
 MUX2_X1 _339_ (.A(net20),
    .B(\dr_shift_reg[28] ),
    .S(_120_),
    .Z(_121_));
 MUX2_X1 _340_ (.A(\dr_shift_reg[27] ),
    .B(_121_),
    .S(_112_),
    .Z(_045_));
 MUX2_X1 _341_ (.A(net21),
    .B(\dr_shift_reg[29] ),
    .S(_120_),
    .Z(_122_));
 MUX2_X1 _342_ (.A(\dr_shift_reg[28] ),
    .B(_122_),
    .S(_112_),
    .Z(_046_));
 MUX2_X1 _343_ (.A(net22),
    .B(\dr_shift_reg[30] ),
    .S(_120_),
    .Z(_123_));
 BUF_X8 _344_ (.A(_094_),
    .Z(_124_));
 MUX2_X1 _345_ (.A(\dr_shift_reg[29] ),
    .B(_123_),
    .S(_124_),
    .Z(_047_));
 MUX2_X1 _346_ (.A(net23),
    .B(\dr_shift_reg[3] ),
    .S(_120_),
    .Z(_125_));
 MUX2_X1 _347_ (.A(\dr_shift_reg[2] ),
    .B(_125_),
    .S(_124_),
    .Z(_048_));
 MUX2_X1 _348_ (.A(\dr_shift_reg[30] ),
    .B(\dr_shift_reg[31] ),
    .S(net68),
    .Z(_126_));
 MUX2_X1 _349_ (.A(net24),
    .B(_126_),
    .S(_097_),
    .Z(_049_));
 MUX2_X1 _350_ (.A(net25),
    .B(net34),
    .S(_120_),
    .Z(_127_));
 MUX2_X1 _351_ (.A(\dr_shift_reg[31] ),
    .B(_127_),
    .S(_124_),
    .Z(_050_));
 MUX2_X1 _352_ (.A(net26),
    .B(\dr_shift_reg[4] ),
    .S(_120_),
    .Z(_128_));
 MUX2_X1 _353_ (.A(\dr_shift_reg[3] ),
    .B(_128_),
    .S(_124_),
    .Z(_051_));
 MUX2_X1 _354_ (.A(net27),
    .B(\dr_shift_reg[5] ),
    .S(_120_),
    .Z(_129_));
 MUX2_X1 _355_ (.A(\dr_shift_reg[4] ),
    .B(_129_),
    .S(_124_),
    .Z(_052_));
 MUX2_X1 _356_ (.A(net28),
    .B(\dr_shift_reg[6] ),
    .S(_120_),
    .Z(_130_));
 MUX2_X1 _357_ (.A(\dr_shift_reg[5] ),
    .B(_130_),
    .S(_124_),
    .Z(_053_));
 MUX2_X1 _358_ (.A(net29),
    .B(\dr_shift_reg[7] ),
    .S(_120_),
    .Z(_131_));
 MUX2_X1 _359_ (.A(\dr_shift_reg[6] ),
    .B(_131_),
    .S(_124_),
    .Z(_054_));
 MUX2_X1 _360_ (.A(net30),
    .B(\dr_shift_reg[8] ),
    .S(_120_),
    .Z(_132_));
 MUX2_X1 _361_ (.A(\dr_shift_reg[7] ),
    .B(_132_),
    .S(_124_),
    .Z(_055_));
 MUX2_X1 _362_ (.A(net31),
    .B(\dr_shift_reg[9] ),
    .S(_093_),
    .Z(_133_));
 MUX2_X1 _363_ (.A(\dr_shift_reg[8] ),
    .B(_133_),
    .S(_124_),
    .Z(_056_));
 MUX2_X1 _364_ (.A(net32),
    .B(\dr_shift_reg[10] ),
    .S(_093_),
    .Z(_134_));
 MUX2_X1 _365_ (.A(\dr_shift_reg[9] ),
    .B(_134_),
    .S(_124_),
    .Z(_057_));
 INV_X2 _366_ (.A(_078_),
    .ZN(_135_));
 OR2_X1 _367_ (.A1(_135_),
    .A2(\ir_shift_reg[1] ),
    .ZN(_136_));
 NAND2_X2 _368_ (.A1(_082_),
    .A2(_085_),
    .ZN(_137_));
 MUX2_X1 _369_ (.A(_136_),
    .B(\ir_shift_reg[0] ),
    .S(_137_),
    .Z(_063_));
 OR2_X1 _370_ (.A1(_135_),
    .A2(\ir_shift_reg[2] ),
    .ZN(_138_));
 MUX2_X1 _371_ (.A(_138_),
    .B(\ir_shift_reg[1] ),
    .S(_137_),
    .Z(_064_));
 OR2_X1 _372_ (.A1(_135_),
    .A2(\ir_shift_reg[3] ),
    .ZN(_139_));
 MUX2_X1 _373_ (.A(_139_),
    .B(\ir_shift_reg[2] ),
    .S(_137_),
    .Z(_065_));
 OR2_X1 _374_ (.A1(_135_),
    .A2(\ir_shift_reg[4] ),
    .ZN(_140_));
 MUX2_X1 _375_ (.A(_140_),
    .B(\ir_shift_reg[3] ),
    .S(_137_),
    .Z(_066_));
 AND2_X1 _376_ (.A1(_078_),
    .A2(net34),
    .ZN(_141_));
 MUX2_X1 _377_ (.A(_141_),
    .B(\ir_shift_reg[4] ),
    .S(_137_),
    .Z(_067_));
 MUX2_X1 _378_ (.A(\dr_shift_reg[0] ),
    .B(net36),
    .S(_090_),
    .Z(_068_));
 MUX2_X1 _379_ (.A(\dr_shift_reg[10] ),
    .B(net37),
    .S(_090_),
    .Z(_069_));
 MUX2_X1 _380_ (.A(\dr_shift_reg[11] ),
    .B(net38),
    .S(_090_),
    .Z(_070_));
 MUX2_X1 _381_ (.A(\dr_shift_reg[12] ),
    .B(net39),
    .S(_090_),
    .Z(_071_));
 MUX2_X1 _382_ (.A(\dr_shift_reg[13] ),
    .B(net40),
    .S(_090_),
    .Z(_072_));
 MUX2_X1 _383_ (.A(\dr_shift_reg[14] ),
    .B(net41),
    .S(_087_),
    .Z(_073_));
 MUX2_X1 _384_ (.A(\dr_shift_reg[15] ),
    .B(net42),
    .S(_087_),
    .Z(_074_));
 MUX2_X1 _385_ (.A(\dr_shift_reg[16] ),
    .B(net43),
    .S(_087_),
    .Z(_075_));
 NAND2_X1 _386_ (.A1(_076_),
    .A2(_084_),
    .ZN(_142_));
 OR2_X2 _387_ (.A1(_083_),
    .A2(_142_),
    .ZN(_143_));
 MUX2_X1 _388_ (.A(\ir_shift_reg[0] ),
    .B(net69),
    .S(_143_),
    .Z(_058_));
 MUX2_X1 _389_ (.A(\ir_shift_reg[1] ),
    .B(net70),
    .S(_143_),
    .Z(_059_));
 MUX2_X1 _390_ (.A(\ir_shift_reg[2] ),
    .B(net71),
    .S(_143_),
    .Z(_060_));
 MUX2_X1 _391_ (.A(\ir_shift_reg[3] ),
    .B(net72),
    .S(_143_),
    .Z(_061_));
 MUX2_X1 _392_ (.A(\ir_shift_reg[4] ),
    .B(net73),
    .S(_143_),
    .Z(_062_));
 INV_X1 _393_ (.A(_084_),
    .ZN(_144_));
 BUF_X2 _394_ (.A(tms),
    .Z(_145_));
 INV_X1 _395_ (.A(_145_),
    .ZN(_146_));
 AOI21_X1 _396_ (.A(_084_),
    .B1(_146_),
    .B2(_082_),
    .ZN(_147_));
 OAI22_X1 _397_ (.A1(_144_),
    .A2(_145_),
    .B1(_147_),
    .B2(_135_),
    .ZN(_148_));
 NAND2_X1 _398_ (.A1(_076_),
    .A2(_145_),
    .ZN(_149_));
 AOI21_X1 _399_ (.A(_145_),
    .B1(_076_),
    .B2(_078_),
    .ZN(_150_));
 OAI21_X1 _400_ (.A(_149_),
    .B1(_150_),
    .B2(_082_),
    .ZN(_151_));
 OAI21_X1 _401_ (.A(_084_),
    .B1(_149_),
    .B2(_135_),
    .ZN(_152_));
 AOI22_X1 _402_ (.A1(_077_),
    .A2(_148_),
    .B1(_151_),
    .B2(_152_),
    .ZN(\next_tap_state[0] ));
 XNOR2_X1 _403_ (.A(_084_),
    .B(_145_),
    .ZN(_153_));
 NOR3_X1 _404_ (.A1(_082_),
    .A2(_076_),
    .A3(_153_),
    .ZN(_154_));
 NOR3_X1 _405_ (.A1(_077_),
    .A2(_084_),
    .A3(_145_),
    .ZN(_155_));
 OAI21_X1 _406_ (.A(_078_),
    .B1(_154_),
    .B2(_155_),
    .ZN(_156_));
 NOR2_X1 _407_ (.A1(_084_),
    .A2(_146_),
    .ZN(_157_));
 MUX2_X1 _408_ (.A(_149_),
    .B(_157_),
    .S(_082_),
    .Z(_158_));
 OAI221_X1 _409_ (.A(_156_),
    .B1(_142_),
    .B2(_146_),
    .C1(_078_),
    .C2(_158_),
    .ZN(\next_tap_state[1] ));
 AND2_X1 _410_ (.A1(_078_),
    .A2(_145_),
    .ZN(_159_));
 AOI21_X1 _411_ (.A(_144_),
    .B1(_159_),
    .B2(_077_),
    .ZN(_160_));
 NOR2_X1 _412_ (.A1(_082_),
    .A2(_160_),
    .ZN(_161_));
 NAND2_X1 _413_ (.A1(_084_),
    .A2(_159_),
    .ZN(_162_));
 OAI21_X1 _414_ (.A(_162_),
    .B1(_145_),
    .B2(_077_),
    .ZN(_163_));
 AOI221_X1 _415_ (.A(_161_),
    .B1(_092_),
    .B2(_135_),
    .C1(_082_),
    .C2(_163_),
    .ZN(\next_tap_state[2] ));
 AOI21_X1 _416_ (.A(_146_),
    .B1(_084_),
    .B2(_135_),
    .ZN(_164_));
 OAI21_X1 _417_ (.A(_143_),
    .B1(_164_),
    .B2(_076_),
    .ZN(_165_));
 NOR2_X1 _418_ (.A1(_135_),
    .A2(_145_),
    .ZN(_166_));
 OAI22_X1 _419_ (.A1(_135_),
    .A2(_076_),
    .B1(_166_),
    .B2(_082_),
    .ZN(_167_));
 AOI21_X1 _420_ (.A(_165_),
    .B1(_167_),
    .B2(_144_),
    .ZN(\next_tap_state[3] ));
 DFFR_X1 \dr_reg[0]$_DFFE_NN0P_  (.D(_068_),
    .RN(net35),
    .CK(_001_),
    .Q(net36),
    .QN(_242_));
 DFFR_X1 \dr_reg[10]$_DFFE_NN0P_  (.D(_069_),
    .RN(net35),
    .CK(_001_),
    .Q(net37),
    .QN(_241_));
 DFFR_X1 \dr_reg[11]$_DFFE_NN0P_  (.D(_070_),
    .RN(net35),
    .CK(_001_),
    .Q(net38),
    .QN(_240_));
 DFFR_X1 \dr_reg[12]$_DFFE_NN0P_  (.D(_071_),
    .RN(net35),
    .CK(_001_),
    .Q(net39),
    .QN(_239_));
 DFFR_X1 \dr_reg[13]$_DFFE_NN0P_  (.D(_072_),
    .RN(net35),
    .CK(_001_),
    .Q(net40),
    .QN(_238_));
 DFFR_X1 \dr_reg[14]$_DFFE_NN0P_  (.D(_073_),
    .RN(net35),
    .CK(_001_),
    .Q(net41),
    .QN(_237_));
 DFFR_X1 \dr_reg[15]$_DFFE_NN0P_  (.D(_074_),
    .RN(net35),
    .CK(_001_),
    .Q(net42),
    .QN(_236_));
 DFFR_X1 \dr_reg[16]$_DFFE_NN0P_  (.D(_075_),
    .RN(net35),
    .CK(_001_),
    .Q(net43),
    .QN(_235_));
 DFFR_X1 \dr_reg[17]$_DFFE_NN0P_  (.D(_002_),
    .RN(net35),
    .CK(_001_),
    .Q(net44),
    .QN(_234_));
 DFFR_X1 \dr_reg[18]$_DFFE_NN0P_  (.D(_003_),
    .RN(net35),
    .CK(_001_),
    .Q(net45),
    .QN(_233_));
 DFFR_X1 \dr_reg[19]$_DFFE_NN0P_  (.D(_004_),
    .RN(net35),
    .CK(_001_),
    .Q(net46),
    .QN(_232_));
 DFFR_X1 \dr_reg[1]$_DFFE_NN0P_  (.D(_005_),
    .RN(net35),
    .CK(_001_),
    .Q(net47),
    .QN(_231_));
 DFFR_X1 \dr_reg[20]$_DFFE_NN0P_  (.D(_006_),
    .RN(net35),
    .CK(_001_),
    .Q(net48),
    .QN(_230_));
 DFFR_X1 \dr_reg[21]$_DFFE_NN0P_  (.D(_007_),
    .RN(net35),
    .CK(_001_),
    .Q(net49),
    .QN(_229_));
 DFFR_X1 \dr_reg[22]$_DFFE_NN0P_  (.D(_008_),
    .RN(net35),
    .CK(_001_),
    .Q(net50),
    .QN(_228_));
 DFFR_X1 \dr_reg[23]$_DFFE_NN0P_  (.D(_009_),
    .RN(net35),
    .CK(_001_),
    .Q(net51),
    .QN(_227_));
 DFFR_X1 \dr_reg[24]$_DFFE_NN0P_  (.D(_010_),
    .RN(net35),
    .CK(_001_),
    .Q(net52),
    .QN(_226_));
 DFFR_X1 \dr_reg[25]$_DFFE_NN0P_  (.D(_011_),
    .RN(net35),
    .CK(_001_),
    .Q(net53),
    .QN(_225_));
 DFFR_X1 \dr_reg[26]$_DFFE_NN0P_  (.D(_012_),
    .RN(net35),
    .CK(_001_),
    .Q(net54),
    .QN(_224_));
 DFFR_X1 \dr_reg[27]$_DFFE_NN0P_  (.D(_013_),
    .RN(net35),
    .CK(_001_),
    .Q(net55),
    .QN(_223_));
 DFFR_X1 \dr_reg[28]$_DFFE_NN0P_  (.D(_014_),
    .RN(net35),
    .CK(_001_),
    .Q(net56),
    .QN(_222_));
 DFFR_X1 \dr_reg[29]$_DFFE_NN0P_  (.D(_015_),
    .RN(net35),
    .CK(_001_),
    .Q(net57),
    .QN(_221_));
 DFFR_X1 \dr_reg[2]$_DFFE_NN0P_  (.D(_016_),
    .RN(net35),
    .CK(_001_),
    .Q(net58),
    .QN(_220_));
 DFFR_X1 \dr_reg[30]$_DFFE_NN0P_  (.D(_017_),
    .RN(net35),
    .CK(_001_),
    .Q(net59),
    .QN(_219_));
 DFFR_X1 \dr_reg[31]$_DFFE_NN0P_  (.D(_018_),
    .RN(net35),
    .CK(_001_),
    .Q(net60),
    .QN(_218_));
 DFFR_X1 \dr_reg[3]$_DFFE_NN0P_  (.D(_019_),
    .RN(net35),
    .CK(_001_),
    .Q(net61),
    .QN(_217_));
 DFFR_X1 \dr_reg[4]$_DFFE_NN0P_  (.D(_020_),
    .RN(net35),
    .CK(_001_),
    .Q(net62),
    .QN(_216_));
 DFFR_X1 \dr_reg[5]$_DFFE_NN0P_  (.D(_021_),
    .RN(net35),
    .CK(_001_),
    .Q(net63),
    .QN(_215_));
 DFFR_X1 \dr_reg[6]$_DFFE_NN0P_  (.D(_022_),
    .RN(net35),
    .CK(_001_),
    .Q(net64),
    .QN(_214_));
 DFFR_X1 \dr_reg[7]$_DFFE_NN0P_  (.D(_023_),
    .RN(net35),
    .CK(_001_),
    .Q(net65),
    .QN(_213_));
 DFFR_X1 \dr_reg[8]$_DFFE_NN0P_  (.D(_024_),
    .RN(net35),
    .CK(_001_),
    .Q(net66),
    .QN(_212_));
 DFFR_X1 \dr_reg[9]$_DFFE_NN0P_  (.D(_025_),
    .RN(net35),
    .CK(_001_),
    .Q(net67),
    .QN(_211_));
 DFFR_X1 \dr_shift_reg[0]$_DFFE_PN0P_  (.D(_026_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[0] ),
    .QN(_210_));
 DFFR_X1 \dr_shift_reg[10]$_DFFE_PN0P_  (.D(_027_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[10] ),
    .QN(_209_));
 DFFR_X1 \dr_shift_reg[11]$_DFFE_PN0P_  (.D(_028_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[11] ),
    .QN(_208_));
 DFFR_X1 \dr_shift_reg[12]$_DFFE_PN0P_  (.D(_029_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[12] ),
    .QN(_207_));
 DFFR_X1 \dr_shift_reg[13]$_DFFE_PN0P_  (.D(_030_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[13] ),
    .QN(_206_));
 DFFR_X1 \dr_shift_reg[14]$_DFFE_PN0P_  (.D(_031_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[14] ),
    .QN(_205_));
 DFFR_X1 \dr_shift_reg[15]$_DFFE_PN0P_  (.D(_032_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[15] ),
    .QN(_204_));
 DFFR_X1 \dr_shift_reg[16]$_DFFE_PN0P_  (.D(_033_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[16] ),
    .QN(_203_));
 DFFR_X1 \dr_shift_reg[17]$_DFFE_PN0P_  (.D(_034_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[17] ),
    .QN(_202_));
 DFFR_X1 \dr_shift_reg[18]$_DFFE_PN0P_  (.D(_035_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[18] ),
    .QN(_201_));
 DFFR_X1 \dr_shift_reg[19]$_DFFE_PN0P_  (.D(_036_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[19] ),
    .QN(_200_));
 DFFR_X1 \dr_shift_reg[1]$_DFFE_PN0P_  (.D(_037_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[1] ),
    .QN(_199_));
 DFFR_X1 \dr_shift_reg[20]$_DFFE_PN0P_  (.D(_038_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[20] ),
    .QN(_198_));
 DFFR_X1 \dr_shift_reg[21]$_DFFE_PN0P_  (.D(_039_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[21] ),
    .QN(_197_));
 DFFR_X1 \dr_shift_reg[22]$_DFFE_PN0P_  (.D(_040_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[22] ),
    .QN(_196_));
 DFFR_X1 \dr_shift_reg[23]$_DFFE_PN0P_  (.D(_041_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[23] ),
    .QN(_195_));
 DFFR_X1 \dr_shift_reg[24]$_DFFE_PN0P_  (.D(_042_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[24] ),
    .QN(_194_));
 DFFR_X1 \dr_shift_reg[25]$_DFFE_PN0P_  (.D(_043_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[25] ),
    .QN(_193_));
 DFFR_X1 \dr_shift_reg[26]$_DFFE_PN0P_  (.D(_044_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[26] ),
    .QN(_192_));
 DFFR_X1 \dr_shift_reg[27]$_DFFE_PN0P_  (.D(_045_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[27] ),
    .QN(_191_));
 DFFR_X1 \dr_shift_reg[28]$_DFFE_PN0P_  (.D(_046_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[28] ),
    .QN(_190_));
 DFFR_X1 \dr_shift_reg[29]$_DFFE_PN0P_  (.D(_047_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[29] ),
    .QN(_189_));
 DFFR_X1 \dr_shift_reg[2]$_DFFE_PN0P_  (.D(_048_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[2] ),
    .QN(_188_));
 DFFR_X1 \dr_shift_reg[30]$_DFFE_PN0P_  (.D(_049_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[30] ),
    .QN(_187_));
 DFFR_X1 \dr_shift_reg[31]$_DFFE_PN0P_  (.D(_050_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[31] ),
    .QN(_186_));
 DFFR_X1 \dr_shift_reg[3]$_DFFE_PN0P_  (.D(_051_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[3] ),
    .QN(_185_));
 DFFR_X1 \dr_shift_reg[4]$_DFFE_PN0P_  (.D(_052_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[4] ),
    .QN(_184_));
 DFFR_X1 \dr_shift_reg[5]$_DFFE_PN0P_  (.D(_053_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[5] ),
    .QN(_183_));
 DFFR_X1 \dr_shift_reg[6]$_DFFE_PN0P_  (.D(_054_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[6] ),
    .QN(_182_));
 DFFR_X1 \dr_shift_reg[7]$_DFFE_PN0P_  (.D(_055_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[7] ),
    .QN(_181_));
 DFFR_X1 \dr_shift_reg[8]$_DFFE_PN0P_  (.D(_056_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[8] ),
    .QN(_180_));
 DFFR_X1 \dr_shift_reg[9]$_DFFE_PN0P_  (.D(_057_),
    .RN(net35),
    .CK(net33),
    .Q(\dr_shift_reg[9] ),
    .QN(_179_));
 DFFS_X1 \ir_reg[0]$_DFFE_NN1N_  (.D(_058_),
    .SN(net35),
    .CK(_001_),
    .Q(net69),
    .QN(_178_));
 DFFR_X1 \ir_reg[1]$_DFFE_NN0N_  (.D(_059_),
    .RN(net35),
    .CK(_001_),
    .Q(net70),
    .QN(_177_));
 DFFR_X1 \ir_reg[2]$_DFFE_NN0N_  (.D(_060_),
    .RN(net35),
    .CK(_001_),
    .Q(net71),
    .QN(_176_));
 DFFR_X1 \ir_reg[3]$_DFFE_NN0N_  (.D(_061_),
    .RN(net35),
    .CK(_001_),
    .Q(net72),
    .QN(_175_));
 DFFR_X1 \ir_reg[4]$_DFFE_NN0N_  (.D(_062_),
    .RN(net35),
    .CK(_001_),
    .Q(net73),
    .QN(_174_));
 DFFS_X1 \ir_shift_reg[0]$_DFFE_PN1P_  (.D(_063_),
    .SN(net35),
    .CK(net33),
    .Q(\ir_shift_reg[0] ),
    .QN(_173_));
 DFFR_X1 \ir_shift_reg[1]$_DFFE_PN0P_  (.D(_064_),
    .RN(net35),
    .CK(net33),
    .Q(\ir_shift_reg[1] ),
    .QN(_172_));
 DFFR_X1 \ir_shift_reg[2]$_DFFE_PN0P_  (.D(_065_),
    .RN(net35),
    .CK(net33),
    .Q(\ir_shift_reg[2] ),
    .QN(_171_));
 DFFR_X1 \ir_shift_reg[3]$_DFFE_PN0P_  (.D(_066_),
    .RN(net35),
    .CK(net33),
    .Q(\ir_shift_reg[3] ),
    .QN(_170_));
 DFFR_X1 \ir_shift_reg[4]$_DFFE_PN0P_  (.D(_067_),
    .RN(net35),
    .CK(net33),
    .Q(\ir_shift_reg[4] ),
    .QN(_243_));
 DFFR_X1 \tap_state[0]$_DFF_PN0_  (.D(\next_tap_state[0] ),
    .RN(net35),
    .CK(net33),
    .Q(\tap_state[0] ),
    .QN(_244_));
 DFFR_X1 \tap_state[1]$_DFF_PN0_  (.D(\next_tap_state[1] ),
    .RN(net35),
    .CK(net33),
    .Q(\tap_state[1] ),
    .QN(_245_));
 DFFR_X2 \tap_state[2]$_DFF_PN0_  (.D(\next_tap_state[2] ),
    .RN(net35),
    .CK(net33),
    .Q(\tap_state[2] ),
    .QN(_246_));
 DFFR_X1 \tap_state[3]$_DFF_PN0_  (.D(\next_tap_state[3] ),
    .RN(net35),
    .CK(net33),
    .Q(\tap_state[3] ),
    .QN(_169_));
 DFFR_X1 \tdo_mux$_DFF_NN0_  (.D(_000_),
    .RN(net35),
    .CK(_001_),
    .Q(net74),
    .QN(_168_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_51 ();
 BUF_X1 input1 (.A(dr_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(dr_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(dr_in[11]),
    .Z(net3));
 BUF_X1 input4 (.A(dr_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(dr_in[13]),
    .Z(net5));
 BUF_X1 input6 (.A(dr_in[14]),
    .Z(net6));
 BUF_X1 input7 (.A(dr_in[15]),
    .Z(net7));
 BUF_X1 input8 (.A(dr_in[16]),
    .Z(net8));
 BUF_X1 input9 (.A(dr_in[17]),
    .Z(net9));
 BUF_X1 input10 (.A(dr_in[18]),
    .Z(net10));
 BUF_X1 input11 (.A(dr_in[19]),
    .Z(net11));
 BUF_X1 input12 (.A(dr_in[1]),
    .Z(net12));
 BUF_X1 input13 (.A(dr_in[20]),
    .Z(net13));
 BUF_X1 input14 (.A(dr_in[21]),
    .Z(net14));
 BUF_X1 input15 (.A(dr_in[22]),
    .Z(net15));
 BUF_X1 input16 (.A(dr_in[23]),
    .Z(net16));
 BUF_X1 input17 (.A(dr_in[24]),
    .Z(net17));
 BUF_X1 input18 (.A(dr_in[25]),
    .Z(net18));
 BUF_X1 input19 (.A(dr_in[26]),
    .Z(net19));
 BUF_X1 input20 (.A(dr_in[27]),
    .Z(net20));
 BUF_X1 input21 (.A(dr_in[28]),
    .Z(net21));
 BUF_X1 input22 (.A(dr_in[29]),
    .Z(net22));
 BUF_X1 input23 (.A(dr_in[2]),
    .Z(net23));
 BUF_X1 input24 (.A(dr_in[30]),
    .Z(net24));
 BUF_X1 input25 (.A(dr_in[31]),
    .Z(net25));
 BUF_X1 input26 (.A(dr_in[3]),
    .Z(net26));
 BUF_X1 input27 (.A(dr_in[4]),
    .Z(net27));
 BUF_X1 input28 (.A(dr_in[5]),
    .Z(net28));
 BUF_X1 input29 (.A(dr_in[6]),
    .Z(net29));
 BUF_X1 input30 (.A(dr_in[7]),
    .Z(net30));
 BUF_X1 input31 (.A(dr_in[8]),
    .Z(net31));
 BUF_X1 input32 (.A(dr_in[9]),
    .Z(net32));
 BUF_X8 input33 (.A(tck),
    .Z(net33));
 BUF_X1 input34 (.A(tdi),
    .Z(net34));
 BUF_X16 input35 (.A(trst_n),
    .Z(net35));
 BUF_X1 output36 (.A(net36),
    .Z(dr_out[0]));
 BUF_X1 output37 (.A(net37),
    .Z(dr_out[10]));
 BUF_X1 output38 (.A(net38),
    .Z(dr_out[11]));
 BUF_X1 output39 (.A(net39),
    .Z(dr_out[12]));
 BUF_X1 output40 (.A(net40),
    .Z(dr_out[13]));
 BUF_X1 output41 (.A(net41),
    .Z(dr_out[14]));
 BUF_X1 output42 (.A(net42),
    .Z(dr_out[15]));
 BUF_X1 output43 (.A(net43),
    .Z(dr_out[16]));
 BUF_X1 output44 (.A(net44),
    .Z(dr_out[17]));
 BUF_X1 output45 (.A(net45),
    .Z(dr_out[18]));
 BUF_X1 output46 (.A(net46),
    .Z(dr_out[19]));
 BUF_X1 output47 (.A(net47),
    .Z(dr_out[1]));
 BUF_X1 output48 (.A(net48),
    .Z(dr_out[20]));
 BUF_X1 output49 (.A(net49),
    .Z(dr_out[21]));
 BUF_X1 output50 (.A(net50),
    .Z(dr_out[22]));
 BUF_X1 output51 (.A(net51),
    .Z(dr_out[23]));
 BUF_X1 output52 (.A(net52),
    .Z(dr_out[24]));
 BUF_X1 output53 (.A(net53),
    .Z(dr_out[25]));
 BUF_X1 output54 (.A(net54),
    .Z(dr_out[26]));
 BUF_X1 output55 (.A(net55),
    .Z(dr_out[27]));
 BUF_X1 output56 (.A(net56),
    .Z(dr_out[28]));
 BUF_X1 output57 (.A(net57),
    .Z(dr_out[29]));
 BUF_X1 output58 (.A(net58),
    .Z(dr_out[2]));
 BUF_X1 output59 (.A(net59),
    .Z(dr_out[30]));
 BUF_X1 output60 (.A(net60),
    .Z(dr_out[31]));
 BUF_X1 output61 (.A(net61),
    .Z(dr_out[3]));
 BUF_X1 output62 (.A(net62),
    .Z(dr_out[4]));
 BUF_X1 output63 (.A(net63),
    .Z(dr_out[5]));
 BUF_X1 output64 (.A(net64),
    .Z(dr_out[6]));
 BUF_X1 output65 (.A(net65),
    .Z(dr_out[7]));
 BUF_X1 output66 (.A(net66),
    .Z(dr_out[8]));
 BUF_X1 output67 (.A(net67),
    .Z(dr_out[9]));
 BUF_X1 output68 (.A(net68),
    .Z(dr_shift_en));
 BUF_X1 output69 (.A(net69),
    .Z(instruction[0]));
 BUF_X1 output70 (.A(net70),
    .Z(instruction[1]));
 BUF_X1 output71 (.A(net71),
    .Z(instruction[2]));
 BUF_X1 output72 (.A(net72),
    .Z(instruction[3]));
 BUF_X1 output73 (.A(net73),
    .Z(instruction[4]));
 BUF_X1 output74 (.A(net74),
    .Z(tdo));
 BUF_X1 output75 (.A(net75),
    .Z(update_dr));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X2 FILLER_0_17 ();
 FILLCELL_X8 FILLER_0_42 ();
 FILLCELL_X1 FILLER_0_70 ();
 FILLCELL_X1 FILLER_0_74 ();
 FILLCELL_X1 FILLER_0_98 ();
 FILLCELL_X1 FILLER_0_102 ();
 FILLCELL_X2 FILLER_0_109 ();
 FILLCELL_X1 FILLER_0_111 ();
 FILLCELL_X2 FILLER_0_118 ();
 FILLCELL_X1 FILLER_0_120 ();
 FILLCELL_X8 FILLER_0_137 ();
 FILLCELL_X2 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_147 ();
 FILLCELL_X2 FILLER_0_158 ();
 FILLCELL_X32 FILLER_0_163 ();
 FILLCELL_X2 FILLER_0_195 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_19 ();
 FILLCELL_X8 FILLER_1_24 ();
 FILLCELL_X1 FILLER_1_32 ();
 FILLCELL_X8 FILLER_1_40 ();
 FILLCELL_X2 FILLER_1_55 ();
 FILLCELL_X8 FILLER_1_61 ();
 FILLCELL_X4 FILLER_1_69 ();
 FILLCELL_X2 FILLER_1_73 ();
 FILLCELL_X1 FILLER_1_85 ();
 FILLCELL_X4 FILLER_1_106 ();
 FILLCELL_X1 FILLER_1_110 ();
 FILLCELL_X4 FILLER_1_118 ();
 FILLCELL_X2 FILLER_1_122 ();
 FILLCELL_X4 FILLER_1_144 ();
 FILLCELL_X4 FILLER_1_168 ();
 FILLCELL_X4 FILLER_2_1 ();
 FILLCELL_X2 FILLER_2_5 ();
 FILLCELL_X1 FILLER_2_7 ();
 FILLCELL_X2 FILLER_2_35 ();
 FILLCELL_X16 FILLER_2_64 ();
 FILLCELL_X2 FILLER_2_80 ();
 FILLCELL_X1 FILLER_2_82 ();
 FILLCELL_X8 FILLER_2_93 ();
 FILLCELL_X1 FILLER_2_101 ();
 FILLCELL_X2 FILLER_2_122 ();
 FILLCELL_X1 FILLER_2_124 ();
 FILLCELL_X4 FILLER_2_132 ();
 FILLCELL_X2 FILLER_2_136 ();
 FILLCELL_X32 FILLER_2_158 ();
 FILLCELL_X4 FILLER_2_190 ();
 FILLCELL_X2 FILLER_2_194 ();
 FILLCELL_X1 FILLER_2_196 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X8 FILLER_3_17 ();
 FILLCELL_X4 FILLER_3_25 ();
 FILLCELL_X2 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_35 ();
 FILLCELL_X16 FILLER_3_43 ();
 FILLCELL_X1 FILLER_3_59 ();
 FILLCELL_X4 FILLER_3_80 ();
 FILLCELL_X2 FILLER_3_84 ();
 FILLCELL_X8 FILLER_3_113 ();
 FILLCELL_X8 FILLER_3_128 ();
 FILLCELL_X4 FILLER_3_136 ();
 FILLCELL_X2 FILLER_3_140 ();
 FILLCELL_X1 FILLER_3_156 ();
 FILLCELL_X8 FILLER_3_164 ();
 FILLCELL_X16 FILLER_3_179 ();
 FILLCELL_X2 FILLER_3_195 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X1 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_45 ();
 FILLCELL_X32 FILLER_4_89 ();
 FILLCELL_X2 FILLER_4_121 ();
 FILLCELL_X16 FILLER_4_137 ();
 FILLCELL_X2 FILLER_4_153 ();
 FILLCELL_X1 FILLER_4_155 ();
 FILLCELL_X1 FILLER_4_176 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_73 ();
 FILLCELL_X8 FILLER_5_94 ();
 FILLCELL_X16 FILLER_5_142 ();
 FILLCELL_X8 FILLER_5_165 ();
 FILLCELL_X4 FILLER_5_173 ();
 FILLCELL_X2 FILLER_5_177 ();
 FILLCELL_X8 FILLER_5_182 ();
 FILLCELL_X4 FILLER_5_190 ();
 FILLCELL_X4 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_5 ();
 FILLCELL_X8 FILLER_6_10 ();
 FILLCELL_X4 FILLER_6_25 ();
 FILLCELL_X1 FILLER_6_29 ();
 FILLCELL_X4 FILLER_6_34 ();
 FILLCELL_X4 FILLER_6_40 ();
 FILLCELL_X2 FILLER_6_44 ();
 FILLCELL_X1 FILLER_6_46 ();
 FILLCELL_X1 FILLER_6_67 ();
 FILLCELL_X4 FILLER_6_73 ();
 FILLCELL_X2 FILLER_6_77 ();
 FILLCELL_X1 FILLER_6_79 ();
 FILLCELL_X16 FILLER_6_83 ();
 FILLCELL_X2 FILLER_6_99 ();
 FILLCELL_X1 FILLER_6_101 ();
 FILLCELL_X16 FILLER_6_111 ();
 FILLCELL_X4 FILLER_6_127 ();
 FILLCELL_X8 FILLER_6_165 ();
 FILLCELL_X1 FILLER_6_173 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_17 ();
 FILLCELL_X1 FILLER_7_21 ();
 FILLCELL_X1 FILLER_7_60 ();
 FILLCELL_X2 FILLER_7_78 ();
 FILLCELL_X8 FILLER_7_85 ();
 FILLCELL_X4 FILLER_7_93 ();
 FILLCELL_X2 FILLER_7_97 ();
 FILLCELL_X16 FILLER_7_107 ();
 FILLCELL_X1 FILLER_7_123 ();
 FILLCELL_X16 FILLER_7_131 ();
 FILLCELL_X4 FILLER_7_147 ();
 FILLCELL_X2 FILLER_7_151 ();
 FILLCELL_X4 FILLER_7_187 ();
 FILLCELL_X2 FILLER_7_191 ();
 FILLCELL_X1 FILLER_7_193 ();
 FILLCELL_X2 FILLER_8_39 ();
 FILLCELL_X2 FILLER_8_43 ();
 FILLCELL_X1 FILLER_8_45 ();
 FILLCELL_X2 FILLER_8_65 ();
 FILLCELL_X1 FILLER_8_67 ();
 FILLCELL_X4 FILLER_8_73 ();
 FILLCELL_X2 FILLER_8_77 ();
 FILLCELL_X2 FILLER_8_88 ();
 FILLCELL_X8 FILLER_8_110 ();
 FILLCELL_X4 FILLER_8_118 ();
 FILLCELL_X16 FILLER_8_142 ();
 FILLCELL_X8 FILLER_8_165 ();
 FILLCELL_X1 FILLER_8_173 ();
 FILLCELL_X2 FILLER_9_21 ();
 FILLCELL_X1 FILLER_9_23 ();
 FILLCELL_X1 FILLER_9_45 ();
 FILLCELL_X1 FILLER_9_55 ();
 FILLCELL_X1 FILLER_9_69 ();
 FILLCELL_X1 FILLER_9_77 ();
 FILLCELL_X2 FILLER_9_85 ();
 FILLCELL_X8 FILLER_9_90 ();
 FILLCELL_X4 FILLER_9_98 ();
 FILLCELL_X8 FILLER_9_105 ();
 FILLCELL_X4 FILLER_9_113 ();
 FILLCELL_X4 FILLER_9_124 ();
 FILLCELL_X2 FILLER_9_128 ();
 FILLCELL_X1 FILLER_9_130 ();
 FILLCELL_X2 FILLER_9_158 ();
 FILLCELL_X1 FILLER_9_160 ();
 FILLCELL_X4 FILLER_9_188 ();
 FILLCELL_X2 FILLER_9_192 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_9 ();
 FILLCELL_X1 FILLER_10_11 ();
 FILLCELL_X2 FILLER_10_23 ();
 FILLCELL_X8 FILLER_10_29 ();
 FILLCELL_X4 FILLER_10_37 ();
 FILLCELL_X1 FILLER_10_41 ();
 FILLCELL_X4 FILLER_10_53 ();
 FILLCELL_X2 FILLER_10_57 ();
 FILLCELL_X1 FILLER_10_81 ();
 FILLCELL_X8 FILLER_10_91 ();
 FILLCELL_X4 FILLER_10_99 ();
 FILLCELL_X2 FILLER_10_103 ();
 FILLCELL_X8 FILLER_10_112 ();
 FILLCELL_X1 FILLER_10_120 ();
 FILLCELL_X16 FILLER_10_135 ();
 FILLCELL_X8 FILLER_10_151 ();
 FILLCELL_X2 FILLER_10_159 ();
 FILLCELL_X4 FILLER_10_168 ();
 FILLCELL_X2 FILLER_10_172 ();
 FILLCELL_X1 FILLER_10_174 ();
 FILLCELL_X8 FILLER_10_178 ();
 FILLCELL_X8 FILLER_10_189 ();
 FILLCELL_X2 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_3 ();
 FILLCELL_X8 FILLER_11_7 ();
 FILLCELL_X4 FILLER_11_15 ();
 FILLCELL_X2 FILLER_11_19 ();
 FILLCELL_X1 FILLER_11_21 ();
 FILLCELL_X1 FILLER_11_25 ();
 FILLCELL_X32 FILLER_11_53 ();
 FILLCELL_X1 FILLER_11_85 ();
 FILLCELL_X8 FILLER_11_106 ();
 FILLCELL_X2 FILLER_11_114 ();
 FILLCELL_X1 FILLER_11_116 ();
 FILLCELL_X16 FILLER_11_137 ();
 FILLCELL_X1 FILLER_11_153 ();
 FILLCELL_X8 FILLER_11_168 ();
 FILLCELL_X1 FILLER_11_176 ();
 FILLCELL_X1 FILLER_12_4 ();
 FILLCELL_X16 FILLER_12_12 ();
 FILLCELL_X4 FILLER_12_28 ();
 FILLCELL_X32 FILLER_12_35 ();
 FILLCELL_X8 FILLER_12_67 ();
 FILLCELL_X1 FILLER_12_75 ();
 FILLCELL_X4 FILLER_12_90 ();
 FILLCELL_X2 FILLER_12_94 ();
 FILLCELL_X4 FILLER_12_109 ();
 FILLCELL_X2 FILLER_12_113 ();
 FILLCELL_X4 FILLER_12_124 ();
 FILLCELL_X1 FILLER_12_137 ();
 FILLCELL_X1 FILLER_12_158 ();
 FILLCELL_X1 FILLER_12_189 ();
 FILLCELL_X1 FILLER_12_193 ();
 FILLCELL_X1 FILLER_13_28 ();
 FILLCELL_X2 FILLER_13_76 ();
 FILLCELL_X1 FILLER_13_78 ();
 FILLCELL_X8 FILLER_13_99 ();
 FILLCELL_X2 FILLER_13_107 ();
 FILLCELL_X1 FILLER_13_109 ();
 FILLCELL_X16 FILLER_13_130 ();
 FILLCELL_X8 FILLER_13_146 ();
 FILLCELL_X4 FILLER_13_154 ();
 FILLCELL_X2 FILLER_13_158 ();
 FILLCELL_X1 FILLER_13_160 ();
 FILLCELL_X16 FILLER_13_174 ();
 FILLCELL_X4 FILLER_13_190 ();
 FILLCELL_X2 FILLER_13_194 ();
 FILLCELL_X1 FILLER_13_196 ();
 FILLCELL_X2 FILLER_14_7 ();
 FILLCELL_X1 FILLER_14_9 ();
 FILLCELL_X2 FILLER_14_27 ();
 FILLCELL_X1 FILLER_14_29 ();
 FILLCELL_X32 FILLER_14_44 ();
 FILLCELL_X4 FILLER_14_76 ();
 FILLCELL_X2 FILLER_14_80 ();
 FILLCELL_X1 FILLER_14_82 ();
 FILLCELL_X16 FILLER_14_90 ();
 FILLCELL_X8 FILLER_14_106 ();
 FILLCELL_X4 FILLER_14_114 ();
 FILLCELL_X1 FILLER_14_118 ();
 FILLCELL_X2 FILLER_14_121 ();
 FILLCELL_X4 FILLER_14_177 ();
 FILLCELL_X8 FILLER_14_184 ();
 FILLCELL_X2 FILLER_14_192 ();
 FILLCELL_X1 FILLER_15_4 ();
 FILLCELL_X16 FILLER_15_12 ();
 FILLCELL_X2 FILLER_15_28 ();
 FILLCELL_X1 FILLER_15_30 ();
 FILLCELL_X16 FILLER_15_51 ();
 FILLCELL_X4 FILLER_15_67 ();
 FILLCELL_X2 FILLER_15_71 ();
 FILLCELL_X1 FILLER_15_73 ();
 FILLCELL_X32 FILLER_15_100 ();
 FILLCELL_X16 FILLER_15_132 ();
 FILLCELL_X8 FILLER_15_148 ();
 FILLCELL_X2 FILLER_15_156 ();
 FILLCELL_X8 FILLER_15_165 ();
 FILLCELL_X1 FILLER_15_173 ();
 FILLCELL_X2 FILLER_15_194 ();
 FILLCELL_X1 FILLER_15_196 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_25 ();
 FILLCELL_X2 FILLER_16_29 ();
 FILLCELL_X1 FILLER_16_31 ();
 FILLCELL_X2 FILLER_16_35 ();
 FILLCELL_X32 FILLER_16_64 ();
 FILLCELL_X8 FILLER_16_96 ();
 FILLCELL_X16 FILLER_16_131 ();
 FILLCELL_X4 FILLER_16_154 ();
 FILLCELL_X2 FILLER_16_158 ();
 FILLCELL_X1 FILLER_16_160 ();
 FILLCELL_X2 FILLER_16_168 ();
 FILLCELL_X1 FILLER_16_170 ();
 FILLCELL_X16 FILLER_17_45 ();
 FILLCELL_X8 FILLER_17_61 ();
 FILLCELL_X4 FILLER_17_69 ();
 FILLCELL_X1 FILLER_17_73 ();
 FILLCELL_X16 FILLER_17_81 ();
 FILLCELL_X4 FILLER_17_97 ();
 FILLCELL_X16 FILLER_17_108 ();
 FILLCELL_X8 FILLER_17_124 ();
 FILLCELL_X4 FILLER_17_132 ();
 FILLCELL_X8 FILLER_17_183 ();
 FILLCELL_X2 FILLER_17_191 ();
 FILLCELL_X1 FILLER_17_193 ();
 FILLCELL_X2 FILLER_18_4 ();
 FILLCELL_X1 FILLER_18_6 ();
 FILLCELL_X8 FILLER_18_14 ();
 FILLCELL_X4 FILLER_18_22 ();
 FILLCELL_X1 FILLER_18_26 ();
 FILLCELL_X16 FILLER_18_54 ();
 FILLCELL_X4 FILLER_18_70 ();
 FILLCELL_X16 FILLER_18_81 ();
 FILLCELL_X2 FILLER_18_97 ();
 FILLCELL_X1 FILLER_18_99 ();
 FILLCELL_X32 FILLER_18_120 ();
 FILLCELL_X4 FILLER_18_152 ();
 FILLCELL_X2 FILLER_18_156 ();
 FILLCELL_X8 FILLER_18_172 ();
 FILLCELL_X1 FILLER_18_180 ();
 FILLCELL_X8 FILLER_18_184 ();
 FILLCELL_X4 FILLER_18_192 ();
 FILLCELL_X1 FILLER_18_196 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_5 ();
 FILLCELL_X1 FILLER_19_7 ();
 FILLCELL_X2 FILLER_19_28 ();
 FILLCELL_X1 FILLER_19_30 ();
 FILLCELL_X32 FILLER_19_34 ();
 FILLCELL_X4 FILLER_19_66 ();
 FILLCELL_X2 FILLER_19_70 ();
 FILLCELL_X1 FILLER_19_72 ();
 FILLCELL_X8 FILLER_19_93 ();
 FILLCELL_X4 FILLER_19_101 ();
 FILLCELL_X32 FILLER_19_112 ();
 FILLCELL_X8 FILLER_19_144 ();
 FILLCELL_X1 FILLER_19_152 ();
 FILLCELL_X2 FILLER_19_167 ();
 FILLCELL_X1 FILLER_19_169 ();
 FILLCELL_X1 FILLER_20_4 ();
 FILLCELL_X2 FILLER_20_12 ();
 FILLCELL_X1 FILLER_20_14 ();
 FILLCELL_X2 FILLER_20_38 ();
 FILLCELL_X1 FILLER_20_67 ();
 FILLCELL_X1 FILLER_20_75 ();
 FILLCELL_X16 FILLER_20_110 ();
 FILLCELL_X2 FILLER_20_126 ();
 FILLCELL_X1 FILLER_20_135 ();
 FILLCELL_X1 FILLER_20_156 ();
 FILLCELL_X2 FILLER_20_177 ();
 FILLCELL_X4 FILLER_20_186 ();
 FILLCELL_X1 FILLER_20_190 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_5 ();
 FILLCELL_X1 FILLER_21_7 ();
 FILLCELL_X16 FILLER_21_22 ();
 FILLCELL_X8 FILLER_21_38 ();
 FILLCELL_X2 FILLER_21_46 ();
 FILLCELL_X1 FILLER_21_48 ();
 FILLCELL_X2 FILLER_21_56 ();
 FILLCELL_X16 FILLER_21_78 ();
 FILLCELL_X1 FILLER_21_94 ();
 FILLCELL_X4 FILLER_21_122 ();
 FILLCELL_X1 FILLER_21_126 ();
 FILLCELL_X32 FILLER_21_141 ();
 FILLCELL_X1 FILLER_21_173 ();
 FILLCELL_X1 FILLER_22_4 ();
 FILLCELL_X1 FILLER_22_12 ();
 FILLCELL_X2 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_42 ();
 FILLCELL_X1 FILLER_22_50 ();
 FILLCELL_X16 FILLER_22_58 ();
 FILLCELL_X1 FILLER_22_74 ();
 FILLCELL_X4 FILLER_22_89 ();
 FILLCELL_X2 FILLER_22_113 ();
 FILLCELL_X4 FILLER_22_155 ();
 FILLCELL_X1 FILLER_22_159 ();
 FILLCELL_X16 FILLER_22_180 ();
 FILLCELL_X1 FILLER_22_196 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_33 ();
 FILLCELL_X2 FILLER_23_37 ();
 FILLCELL_X4 FILLER_23_59 ();
 FILLCELL_X2 FILLER_23_63 ();
 FILLCELL_X1 FILLER_23_65 ();
 FILLCELL_X4 FILLER_23_93 ();
 FILLCELL_X2 FILLER_23_97 ();
 FILLCELL_X2 FILLER_23_106 ();
 FILLCELL_X1 FILLER_23_108 ();
 FILLCELL_X16 FILLER_23_116 ();
 FILLCELL_X2 FILLER_23_132 ();
 FILLCELL_X1 FILLER_23_134 ();
 FILLCELL_X16 FILLER_23_142 ();
 FILLCELL_X1 FILLER_23_158 ();
 FILLCELL_X8 FILLER_23_166 ();
 FILLCELL_X1 FILLER_23_174 ();
 FILLCELL_X16 FILLER_24_14 ();
 FILLCELL_X1 FILLER_24_30 ();
 FILLCELL_X1 FILLER_24_77 ();
 FILLCELL_X2 FILLER_24_105 ();
 FILLCELL_X2 FILLER_24_130 ();
 FILLCELL_X8 FILLER_24_166 ();
 FILLCELL_X4 FILLER_24_174 ();
 FILLCELL_X2 FILLER_24_178 ();
 FILLCELL_X4 FILLER_24_187 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_33 ();
 FILLCELL_X1 FILLER_25_41 ();
 FILLCELL_X2 FILLER_25_49 ();
 FILLCELL_X4 FILLER_25_57 ();
 FILLCELL_X1 FILLER_25_68 ();
 FILLCELL_X2 FILLER_25_72 ();
 FILLCELL_X1 FILLER_25_74 ();
 FILLCELL_X4 FILLER_25_81 ();
 FILLCELL_X1 FILLER_25_85 ();
 FILLCELL_X2 FILLER_25_89 ();
 FILLCELL_X1 FILLER_25_91 ();
 FILLCELL_X8 FILLER_25_95 ();
 FILLCELL_X1 FILLER_25_103 ();
 FILLCELL_X2 FILLER_25_120 ();
 FILLCELL_X1 FILLER_25_122 ();
 FILLCELL_X2 FILLER_25_126 ();
 FILLCELL_X8 FILLER_25_131 ();
 FILLCELL_X2 FILLER_25_139 ();
 FILLCELL_X1 FILLER_25_141 ();
 FILLCELL_X2 FILLER_25_148 ();
 FILLCELL_X1 FILLER_25_150 ();
 FILLCELL_X8 FILLER_25_184 ();
 FILLCELL_X4 FILLER_25_192 ();
 FILLCELL_X1 FILLER_25_196 ();
endmodule
