module parameterized_ring_counter (clk,
    enable,
    rst_n,
    count);
 input clk;
 input enable;
 input rst_n;
 output [3:0] count;

 wire _0_;
 wire _1_;
 wire _2_;
 wire _3_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4_ (.I0(net4),
    .I1(net7),
    .S(net2),
    .Z(_0_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5_ (.I0(net5),
    .I1(net4),
    .S(net2),
    .Z(_1_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6_ (.I0(net6),
    .I1(net5),
    .S(net2),
    .Z(_2_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7_ (.I0(net7),
    .I1(net6),
    .S(net2),
    .Z(_3_));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \counter_reg[0]$_DFFE_PN1P_  (.D(_0_),
    .SETN(net3),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[1]$_DFFE_PN0P_  (.D(_1_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[2]$_DFFE_PN0P_  (.D(_2_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[3]$_DFFE_PN0P_  (.D(_3_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 hold1 (.I(net3),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_65 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(rst_n),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net4),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net5),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net7),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_240 ();
endmodule
