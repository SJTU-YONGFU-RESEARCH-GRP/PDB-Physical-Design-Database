module sync_preset_register (clk,
    enable,
    rst_n,
    sync_preset,
    sync_rst,
    data_in,
    data_out);
 input clk;
 input enable;
 input rst_n;
 input sync_preset;
 input sync_rst;
 input [7:0] data_in;
 output [7:0] data_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _36_ (.A(net10),
    .ZN(_08_));
 NAND2_X4 _37_ (.A1(_08_),
    .A2(net9),
    .ZN(_09_));
 BUF_X4 _38_ (.A(sync_preset),
    .Z(_10_));
 BUF_X4 _39_ (.A(enable),
    .Z(_11_));
 MUX2_X1 _40_ (.A(net11),
    .B(net1),
    .S(_11_),
    .Z(_12_));
 NOR2_X1 _41_ (.A1(_10_),
    .A2(_12_),
    .ZN(_13_));
 NOR2_X1 _42_ (.A1(_09_),
    .A2(_13_),
    .ZN(_00_));
 MUX2_X1 _43_ (.A(net12),
    .B(net2),
    .S(_11_),
    .Z(_14_));
 NOR2_X1 _44_ (.A1(_10_),
    .A2(_14_),
    .ZN(_15_));
 NOR2_X1 _45_ (.A1(_09_),
    .A2(_15_),
    .ZN(_01_));
 MUX2_X1 _46_ (.A(net13),
    .B(net3),
    .S(_11_),
    .Z(_16_));
 NOR2_X1 _47_ (.A1(_10_),
    .A2(_16_),
    .ZN(_17_));
 NOR2_X1 _48_ (.A1(_09_),
    .A2(_17_),
    .ZN(_02_));
 MUX2_X1 _49_ (.A(net14),
    .B(net4),
    .S(_11_),
    .Z(_18_));
 NOR2_X1 _50_ (.A1(_10_),
    .A2(_18_),
    .ZN(_19_));
 NOR2_X1 _51_ (.A1(_09_),
    .A2(_19_),
    .ZN(_03_));
 MUX2_X1 _52_ (.A(net15),
    .B(net5),
    .S(_11_),
    .Z(_20_));
 NOR2_X1 _53_ (.A1(_10_),
    .A2(_20_),
    .ZN(_21_));
 NOR2_X1 _54_ (.A1(_09_),
    .A2(_21_),
    .ZN(_04_));
 MUX2_X1 _55_ (.A(net16),
    .B(net6),
    .S(_11_),
    .Z(_22_));
 NOR2_X1 _56_ (.A1(_10_),
    .A2(_22_),
    .ZN(_23_));
 NOR2_X1 _57_ (.A1(_09_),
    .A2(_23_),
    .ZN(_05_));
 MUX2_X1 _58_ (.A(net17),
    .B(net7),
    .S(_11_),
    .Z(_24_));
 NOR2_X1 _59_ (.A1(_10_),
    .A2(_24_),
    .ZN(_25_));
 NOR2_X1 _60_ (.A1(_09_),
    .A2(_25_),
    .ZN(_06_));
 MUX2_X1 _61_ (.A(net18),
    .B(net8),
    .S(_11_),
    .Z(_26_));
 NOR2_X1 _62_ (.A1(_10_),
    .A2(_26_),
    .ZN(_27_));
 NOR2_X1 _63_ (.A1(_09_),
    .A2(_27_),
    .ZN(_07_));
 DFF_X1 \data_out[0]$_SDFFE_PP0P_  (.D(_00_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net11),
    .QN(_35_));
 DFF_X1 \data_out[1]$_SDFFE_PP0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_34_));
 DFF_X1 \data_out[2]$_SDFFE_PP0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net13),
    .QN(_33_));
 DFF_X1 \data_out[3]$_SDFFE_PP0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net14),
    .QN(_32_));
 DFF_X1 \data_out[4]$_SDFFE_PP0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net15),
    .QN(_31_));
 DFF_X1 \data_out[5]$_SDFFE_PP0P_  (.D(_05_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_30_));
 DFF_X1 \data_out[6]$_SDFFE_PP0P_  (.D(_06_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_29_));
 DFF_X1 \data_out[7]$_SDFFE_PP0P_  (.D(_07_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_28_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_51 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X1 input9 (.A(rst_n),
    .Z(net9));
 BUF_X1 input10 (.A(sync_rst),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(data_out[0]));
 BUF_X1 output12 (.A(net12),
    .Z(data_out[1]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[2]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[3]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[4]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[5]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[6]));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X2 FILLER_0_65 ();
 FILLCELL_X1 FILLER_0_67 ();
 FILLCELL_X2 FILLER_0_74 ();
 FILLCELL_X1 FILLER_0_76 ();
 FILLCELL_X8 FILLER_0_89 ();
 FILLCELL_X4 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_103 ();
 FILLCELL_X32 FILLER_0_116 ();
 FILLCELL_X32 FILLER_0_148 ();
 FILLCELL_X8 FILLER_0_180 ();
 FILLCELL_X4 FILLER_0_188 ();
 FILLCELL_X1 FILLER_0_192 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X16 FILLER_1_33 ();
 FILLCELL_X8 FILLER_1_49 ();
 FILLCELL_X4 FILLER_1_57 ();
 FILLCELL_X2 FILLER_1_61 ();
 FILLCELL_X1 FILLER_1_90 ();
 FILLCELL_X32 FILLER_1_115 ();
 FILLCELL_X32 FILLER_1_147 ();
 FILLCELL_X8 FILLER_1_179 ();
 FILLCELL_X4 FILLER_1_187 ();
 FILLCELL_X2 FILLER_1_191 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_118 ();
 FILLCELL_X32 FILLER_2_150 ();
 FILLCELL_X8 FILLER_2_182 ();
 FILLCELL_X2 FILLER_2_190 ();
 FILLCELL_X1 FILLER_2_192 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X4 FILLER_3_65 ();
 FILLCELL_X1 FILLER_3_72 ();
 FILLCELL_X1 FILLER_3_82 ();
 FILLCELL_X2 FILLER_3_86 ();
 FILLCELL_X2 FILLER_3_91 ();
 FILLCELL_X1 FILLER_3_99 ();
 FILLCELL_X1 FILLER_3_103 ();
 FILLCELL_X32 FILLER_3_111 ();
 FILLCELL_X32 FILLER_3_143 ();
 FILLCELL_X16 FILLER_3_175 ();
 FILLCELL_X2 FILLER_3_191 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_81 ();
 FILLCELL_X32 FILLER_8_90 ();
 FILLCELL_X32 FILLER_8_122 ();
 FILLCELL_X32 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_186 ();
 FILLCELL_X2 FILLER_8_190 ();
 FILLCELL_X1 FILLER_8_192 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X16 FILLER_13_65 ();
 FILLCELL_X4 FILLER_13_81 ();
 FILLCELL_X32 FILLER_13_90 ();
 FILLCELL_X32 FILLER_13_122 ();
 FILLCELL_X32 FILLER_13_154 ();
 FILLCELL_X4 FILLER_13_186 ();
 FILLCELL_X2 FILLER_13_190 ();
 FILLCELL_X1 FILLER_13_192 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X8 FILLER_14_65 ();
 FILLCELL_X4 FILLER_14_76 ();
 FILLCELL_X2 FILLER_14_80 ();
 FILLCELL_X32 FILLER_14_85 ();
 FILLCELL_X32 FILLER_14_117 ();
 FILLCELL_X32 FILLER_14_149 ();
 FILLCELL_X8 FILLER_14_181 ();
 FILLCELL_X4 FILLER_14_189 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_36 ();
 FILLCELL_X1 FILLER_15_38 ();
 FILLCELL_X16 FILLER_15_42 ();
 FILLCELL_X2 FILLER_15_58 ();
 FILLCELL_X1 FILLER_15_60 ();
 FILLCELL_X32 FILLER_15_85 ();
 FILLCELL_X32 FILLER_15_117 ();
 FILLCELL_X32 FILLER_15_149 ();
 FILLCELL_X8 FILLER_15_181 ();
 FILLCELL_X4 FILLER_15_189 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X16 FILLER_18_65 ();
 FILLCELL_X2 FILLER_18_81 ();
 FILLCELL_X1 FILLER_18_83 ();
 FILLCELL_X32 FILLER_18_89 ();
 FILLCELL_X32 FILLER_18_121 ();
 FILLCELL_X32 FILLER_18_153 ();
 FILLCELL_X8 FILLER_18_185 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X16 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_81 ();
 FILLCELL_X2 FILLER_21_92 ();
 FILLCELL_X1 FILLER_21_94 ();
 FILLCELL_X32 FILLER_21_98 ();
 FILLCELL_X32 FILLER_21_130 ();
 FILLCELL_X16 FILLER_21_162 ();
 FILLCELL_X8 FILLER_21_178 ();
 FILLCELL_X4 FILLER_21_186 ();
 FILLCELL_X2 FILLER_21_190 ();
 FILLCELL_X1 FILLER_21_192 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_65 ();
 FILLCELL_X4 FILLER_22_73 ();
 FILLCELL_X2 FILLER_22_77 ();
 FILLCELL_X1 FILLER_22_82 ();
 FILLCELL_X32 FILLER_22_113 ();
 FILLCELL_X32 FILLER_22_145 ();
 FILLCELL_X16 FILLER_22_177 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X1 FILLER_23_65 ();
 FILLCELL_X4 FILLER_23_83 ();
 FILLCELL_X32 FILLER_23_114 ();
 FILLCELL_X32 FILLER_23_146 ();
 FILLCELL_X8 FILLER_23_178 ();
 FILLCELL_X4 FILLER_23_186 ();
 FILLCELL_X2 FILLER_23_190 ();
 FILLCELL_X1 FILLER_23_192 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X8 FILLER_24_65 ();
 FILLCELL_X4 FILLER_24_73 ();
 FILLCELL_X1 FILLER_24_77 ();
 FILLCELL_X8 FILLER_24_85 ();
 FILLCELL_X4 FILLER_24_93 ();
 FILLCELL_X2 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_99 ();
 FILLCELL_X2 FILLER_24_107 ();
 FILLCELL_X32 FILLER_24_112 ();
 FILLCELL_X32 FILLER_24_144 ();
 FILLCELL_X16 FILLER_24_176 ();
 FILLCELL_X1 FILLER_24_192 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_65 ();
 FILLCELL_X4 FILLER_25_73 ();
 FILLCELL_X16 FILLER_25_83 ();
 FILLCELL_X2 FILLER_25_99 ();
 FILLCELL_X2 FILLER_25_104 ();
 FILLCELL_X1 FILLER_25_106 ();
 FILLCELL_X32 FILLER_25_113 ();
 FILLCELL_X32 FILLER_25_145 ();
 FILLCELL_X16 FILLER_25_177 ();
endmodule
