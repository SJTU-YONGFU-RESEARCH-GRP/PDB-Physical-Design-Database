module parameterized_deserializer (clk,
    enable,
    load,
    rst_n,
    rx_busy,
    rx_done,
    serial_in,
    sync_detected,
    parallel_out);
 input clk;
 input enable;
 input load;
 input rst_n;
 output rx_busy;
 output rx_done;
 input serial_in;
 output sync_detected;
 output [7:0] parallel_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire clknet_0_clk;
 wire \bit_counter[0] ;
 wire \bit_counter[1] ;
 wire \bit_counter[2] ;
 wire \bit_counter[3] ;
 wire \clk_div_counter[0] ;
 wire \clk_div_counter[1] ;
 wire \clk_div_counter[2] ;
 wire \shift_reg[0] ;
 wire \shift_reg[1] ;
 wire \shift_reg[2] ;
 wire \shift_reg[3] ;
 wire \shift_reg[4] ;
 wire \shift_reg[5] ;
 wire \shift_reg[6] ;
 wire \shift_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net17;
 wire net18;

 gf180mcu_fd_sc_mcu9t5v0__buf_4 _082_ (.I(net2),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _083_ (.A1(net2),
    .A2(\state[1] ),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _084_ (.I(_047_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _085_ (.I(\state[0] ),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _086_ (.A1(_046_),
    .A2(net3),
    .B1(_048_),
    .B2(_049_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _087_ (.I(\bit_counter[3] ),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _088_ (.I(\clk_div_counter[2] ),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _089_ (.A1(\bit_counter[2] ),
    .A2(_071_),
    .A3(_051_),
    .A4(_075_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _090_ (.A1(_046_),
    .A2(_050_),
    .A3(\state[2] ),
    .A4(_052_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _091_ (.I(net3),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _092_ (.A1(_046_),
    .A2(_054_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _093_ (.A1(\state[1] ),
    .A2(_055_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _094_ (.A1(_053_),
    .A2(_056_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _095_ (.I(\state[2] ),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _096_ (.A1(_046_),
    .A2(_050_),
    .A3(_052_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _097_ (.A1(\state[0] ),
    .A2(net2),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _098_ (.A1(_057_),
    .A2(_058_),
    .B1(_059_),
    .B2(_054_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _099_ (.I(\clk_div_counter[0] ),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _100_ (.I(\clk_div_counter[1] ),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _101_ (.A1(net2),
    .A2(_051_),
    .A3(\state[2] ),
    .A4(_075_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _102_ (.I(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _103_ (.A1(\state[2] ),
    .A2(_059_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _104_ (.A1(\bit_counter[0] ),
    .A2(_060_),
    .A3(_062_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _105_ (.A1(\bit_counter[0] ),
    .A2(_061_),
    .B(_063_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _106_ (.I(_072_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _107_ (.A1(_060_),
    .A2(_062_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _108_ (.I(\bit_counter[1] ),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _109_ (.A1(_064_),
    .A2(_061_),
    .B1(_065_),
    .B2(_066_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _110_ (.A1(_071_),
    .A2(_051_),
    .A3(_075_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _111_ (.A1(_046_),
    .A2(_067_),
    .B(\bit_counter[2] ),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _112_ (.A1(\state[0] ),
    .A2(\state[2] ),
    .B(_046_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _113_ (.A1(\bit_counter[2] ),
    .A2(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _114_ (.A1(_057_),
    .A2(_052_),
    .A3(_068_),
    .B(_070_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _115_ (.A1(\bit_counter[2] ),
    .A2(\bit_counter[0] ),
    .A3(\bit_counter[1] ),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _116_ (.A1(_060_),
    .A2(_028_),
    .B(_062_),
    .C(\bit_counter[3] ),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _117_ (.A1(\bit_counter[3] ),
    .A2(_060_),
    .A3(_028_),
    .B(_029_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _118_ (.A1(\clk_div_counter[0] ),
    .A2(_079_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _119_ (.I0(\clk_div_counter[0] ),
    .I1(_030_),
    .S(_046_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _120_ (.A1(_046_),
    .A2(_076_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _121_ (.A1(_046_),
    .A2(_074_),
    .B1(_079_),
    .B2(_031_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _122_ (.I0(\clk_div_counter[2] ),
    .I1(_080_),
    .S(_046_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _123_ (.I0(\shift_reg[0] ),
    .I1(net6),
    .S(_048_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _124_ (.I0(\shift_reg[1] ),
    .I1(net7),
    .S(_048_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _125_ (.I0(\shift_reg[2] ),
    .I1(net8),
    .S(_048_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _126_ (.I0(\shift_reg[3] ),
    .I1(net9),
    .S(_048_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _127_ (.I0(\shift_reg[4] ),
    .I1(net10),
    .S(_048_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _128_ (.I0(\shift_reg[5] ),
    .I1(net11),
    .S(_048_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _129_ (.I0(\shift_reg[6] ),
    .I1(net12),
    .S(_048_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _130_ (.I0(\shift_reg[7] ),
    .I1(net13),
    .S(_047_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _131_ (.I(net14),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _132_ (.A1(net2),
    .A2(net3),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _133_ (.A1(net3),
    .A2(_032_),
    .B1(_033_),
    .B2(\state[1] ),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _134_ (.A1(net14),
    .A2(_048_),
    .B1(_034_),
    .B2(\state[0] ),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _135_ (.I(_035_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _136_ (.A1(net15),
    .A2(_059_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _137_ (.A1(_048_),
    .A2(_036_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _138_ (.I(net5),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _139_ (.I(\shift_reg[0] ),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _140_ (.A1(_037_),
    .A2(_061_),
    .B1(_065_),
    .B2(_038_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _141_ (.I(\shift_reg[1] ),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _142_ (.A1(_038_),
    .A2(_061_),
    .B1(_065_),
    .B2(_039_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _143_ (.I(\shift_reg[2] ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _144_ (.A1(_039_),
    .A2(_061_),
    .B1(_065_),
    .B2(_040_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _145_ (.I(\shift_reg[3] ),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _146_ (.A1(_040_),
    .A2(_061_),
    .B1(_065_),
    .B2(_041_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _147_ (.I(\shift_reg[4] ),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _148_ (.A1(_041_),
    .A2(_061_),
    .B1(_065_),
    .B2(_042_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _149_ (.I(\shift_reg[5] ),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _150_ (.A1(_042_),
    .A2(_061_),
    .B1(_065_),
    .B2(_043_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _151_ (.I(\shift_reg[6] ),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _152_ (.A1(_043_),
    .A2(_061_),
    .B1(_065_),
    .B2(_044_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _153_ (.I(\shift_reg[7] ),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _154_ (.A1(_044_),
    .A2(_061_),
    .B1(_065_),
    .B2(_045_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _155_ (.A(\bit_counter[0] ),
    .B(\bit_counter[1] ),
    .CO(_071_),
    .S(_072_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _156_ (.A(_073_),
    .B(_074_),
    .CO(_075_),
    .S(_076_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _157_ (.A(\clk_div_counter[0] ),
    .B(\clk_div_counter[1] ),
    .CO(_077_),
    .S(_078_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _158_ (.A(\clk_div_counter[2] ),
    .B(_077_),
    .CO(_079_),
    .S(_080_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _160_ (.I(net16),
    .Z(sync_detected));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[0]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\bit_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[1]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\bit_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[2]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\bit_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[3]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\bit_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_div_counter[0]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\clk_div_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_div_counter[1]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\clk_div_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_div_counter[2]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\clk_div_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[0]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[1]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[2]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[3]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[4]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[5]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[6]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parallel_out[7]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_busy$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_done$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[0]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[1]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[2]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[3]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[4]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[5]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[6]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[7]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \state[0]$_DFF_PN1_  (.D(_000_),
    .SETN(net4),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFF_PN0_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[2]$_DFF_PN0_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 hold1 (.I(net4),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(net18),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input3 (.I(net17),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(serial_in),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(parallel_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net7),
    .Z(parallel_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net8),
    .Z(parallel_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net9),
    .Z(parallel_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net10),
    .Z(parallel_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net11),
    .Z(parallel_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net12),
    .Z(parallel_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(parallel_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_busy));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_done));
 gf180mcu_fd_sc_mcu9t5v0__tiel _160__15 (.ZN(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(load),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_208 ();
endmodule
