module configurable_lfsr (clk,
    enable,
    load_seed,
    rst_n,
    serial_out,
    parallel_out,
    seed,
    tap_pattern);
 input clk;
 input enable;
 input load_seed;
 input rst_n;
 output serial_out;
 output [7:0] parallel_out;
 input [7:0] seed;
 input [7:0] tap_pattern;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net27;

 gf180mcu_fd_sc_mcu9t5v0__buf_4 _33_ (.I(enable),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _34_ (.I0(net26),
    .I1(net19),
    .S(_08_),
    .Z(_09_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _35_ (.I(load_seed),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _36_ (.I0(_09_),
    .I1(net2),
    .S(_10_),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _37_ (.I0(net19),
    .I1(net20),
    .S(_08_),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _38_ (.I0(_11_),
    .I1(net3),
    .S(_10_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _39_ (.I0(net20),
    .I1(net21),
    .S(_08_),
    .Z(_12_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _40_ (.I0(_12_),
    .I1(net4),
    .S(_10_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _41_ (.I0(net21),
    .I1(net22),
    .S(_08_),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _42_ (.I0(_13_),
    .I1(net5),
    .S(_10_),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _43_ (.I0(net22),
    .I1(net23),
    .S(_08_),
    .Z(_14_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _44_ (.I0(_14_),
    .I1(net6),
    .S(_10_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _45_ (.I0(net23),
    .I1(net24),
    .S(_08_),
    .Z(_15_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _46_ (.I0(_15_),
    .I1(net7),
    .S(_10_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _47_ (.I0(net24),
    .I1(net25),
    .S(_08_),
    .Z(_16_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _48_ (.I0(_16_),
    .I1(net8),
    .S(_10_),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _49_ (.I(_08_),
    .ZN(_17_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _50_ (.A1(net23),
    .A2(net15),
    .Z(_18_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _51_ (.A1(net21),
    .A2(net13),
    .Z(_19_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _52_ (.A1(_18_),
    .A2(_19_),
    .ZN(_20_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _53_ (.A1(net24),
    .A2(net16),
    .Z(_21_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _54_ (.A1(net22),
    .A2(net14),
    .Z(_22_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _55_ (.A1(_20_),
    .A2(_21_),
    .A3(_22_),
    .ZN(_23_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _56_ (.A1(net19),
    .A2(net11),
    .Z(_24_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _57_ (.A1(net10),
    .A2(net26),
    .Z(_25_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _58_ (.A1(_24_),
    .A2(_25_),
    .ZN(_26_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _59_ (.A1(net25),
    .A2(net17),
    .Z(_27_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _60_ (.A1(net20),
    .A2(net12),
    .Z(_28_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _61_ (.A1(_26_),
    .A2(_27_),
    .A3(_28_),
    .ZN(_29_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _62_ (.A1(_23_),
    .A2(_29_),
    .ZN(_30_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _63_ (.A1(_10_),
    .A2(_08_),
    .ZN(_31_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _64_ (.A1(_10_),
    .A2(net9),
    .B1(_31_),
    .B2(net25),
    .ZN(_32_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _65_ (.A1(_10_),
    .A2(_17_),
    .A3(_30_),
    .B(_32_),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _66_ (.I(net26),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[4]$_DFFE_PN0P_  (.D(_04_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[5]$_DFFE_PN0P_  (.D(_05_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[6]$_DFFE_PN0P_  (.D(_06_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg[7]$_DFFE_PN0P_  (.D(_07_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 hold1 (.I(net27),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(seed[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(seed[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(seed[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(seed[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(seed[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(seed[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(seed[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(seed[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tap_pattern[0]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tap_pattern[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(tap_pattern[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(tap_pattern[3]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(tap_pattern[4]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(tap_pattern[5]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(tap_pattern[6]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(tap_pattern[7]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(parallel_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(parallel_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(parallel_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(parallel_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(parallel_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(parallel_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(parallel_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(parallel_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net26),
    .Z(serial_out));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_208 ();
endmodule
