module floating_point_adder (clk,
    inexact,
    invalid_op,
    overflow,
    rst_n,
    underflow,
    valid_in,
    valid_out,
    a,
    b,
    result);
 input clk;
 output inexact;
 output invalid_op;
 output overflow;
 input rst_n;
 output underflow;
 input valid_in;
 output valid_out;
 input [31:0] a;
 input [31:0] b;
 output [31:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire a_exp_larger;
 wire a_sign_stage1;
 wire \add_result[10] ;
 wire \add_result[11] ;
 wire \add_result[12] ;
 wire \add_result[13] ;
 wire \add_result[14] ;
 wire \add_result[15] ;
 wire \add_result[16] ;
 wire \add_result[17] ;
 wire \add_result[18] ;
 wire \add_result[19] ;
 wire \add_result[20] ;
 wire \add_result[21] ;
 wire \add_result[22] ;
 wire \add_result[23] ;
 wire \add_result[24] ;
 wire \add_result[25] ;
 wire \add_result[26] ;
 wire \add_result[2] ;
 wire \add_result[3] ;
 wire \add_result[4] ;
 wire \add_result[5] ;
 wire \add_result[6] ;
 wire \add_result[7] ;
 wire \add_result[8] ;
 wire \add_result[9] ;
 wire \aligned_a_mant[0] ;
 wire \aligned_a_mant[10] ;
 wire \aligned_a_mant[11] ;
 wire \aligned_a_mant[12] ;
 wire \aligned_a_mant[13] ;
 wire \aligned_a_mant[14] ;
 wire \aligned_a_mant[15] ;
 wire \aligned_a_mant[16] ;
 wire \aligned_a_mant[17] ;
 wire \aligned_a_mant[18] ;
 wire \aligned_a_mant[19] ;
 wire \aligned_a_mant[1] ;
 wire \aligned_a_mant[20] ;
 wire \aligned_a_mant[21] ;
 wire \aligned_a_mant[22] ;
 wire \aligned_a_mant[23] ;
 wire \aligned_a_mant[24] ;
 wire \aligned_a_mant[25] ;
 wire \aligned_a_mant[2] ;
 wire \aligned_a_mant[3] ;
 wire \aligned_a_mant[4] ;
 wire \aligned_a_mant[5] ;
 wire \aligned_a_mant[6] ;
 wire \aligned_a_mant[7] ;
 wire \aligned_a_mant[8] ;
 wire \aligned_a_mant[9] ;
 wire \aligned_b_mant[0] ;
 wire \aligned_b_mant[10] ;
 wire \aligned_b_mant[11] ;
 wire \aligned_b_mant[12] ;
 wire \aligned_b_mant[13] ;
 wire \aligned_b_mant[14] ;
 wire \aligned_b_mant[15] ;
 wire \aligned_b_mant[16] ;
 wire \aligned_b_mant[17] ;
 wire \aligned_b_mant[18] ;
 wire \aligned_b_mant[19] ;
 wire \aligned_b_mant[1] ;
 wire \aligned_b_mant[20] ;
 wire \aligned_b_mant[21] ;
 wire \aligned_b_mant[22] ;
 wire \aligned_b_mant[23] ;
 wire \aligned_b_mant[24] ;
 wire \aligned_b_mant[25] ;
 wire \aligned_b_mant[2] ;
 wire \aligned_b_mant[3] ;
 wire \aligned_b_mant[4] ;
 wire \aligned_b_mant[5] ;
 wire \aligned_b_mant[6] ;
 wire \aligned_b_mant[7] ;
 wire \aligned_b_mant[8] ;
 wire \aligned_b_mant[9] ;
 wire b_sign_stage1;
 wire \final_exp[0] ;
 wire \final_exp[1] ;
 wire \final_exp[2] ;
 wire \final_exp[3] ;
 wire \final_exp[4] ;
 wire \final_exp[5] ;
 wire \final_exp[6] ;
 wire \final_exp[7] ;
 wire \final_mant[0] ;
 wire \final_mant[10] ;
 wire \final_mant[11] ;
 wire \final_mant[12] ;
 wire \final_mant[13] ;
 wire \final_mant[14] ;
 wire \final_mant[15] ;
 wire \final_mant[16] ;
 wire \final_mant[17] ;
 wire \final_mant[18] ;
 wire \final_mant[19] ;
 wire \final_mant[1] ;
 wire \final_mant[20] ;
 wire \final_mant[21] ;
 wire \final_mant[22] ;
 wire \final_mant[2] ;
 wire \final_mant[3] ;
 wire \final_mant[4] ;
 wire \final_mant[5] ;
 wire \final_mant[6] ;
 wire \final_mant[7] ;
 wire \final_mant[8] ;
 wire \final_mant[9] ;
 wire inexact_stage2;
 wire invalid_op_stage2;
 wire is_a_larger_stage1;
 wire \larger_exp_stage1[0] ;
 wire \larger_exp_stage1[1] ;
 wire \larger_exp_stage1[2] ;
 wire \larger_exp_stage1[3] ;
 wire \larger_exp_stage1[4] ;
 wire \larger_exp_stage1[5] ;
 wire \larger_exp_stage1[6] ;
 wire \larger_exp_stage1[7] ;
 wire \result_exp_stage2[0] ;
 wire \result_exp_stage2[1] ;
 wire \result_exp_stage2[2] ;
 wire \result_exp_stage2[3] ;
 wire \result_exp_stage2[4] ;
 wire \result_exp_stage2[5] ;
 wire \result_exp_stage2[6] ;
 wire \result_exp_stage2[7] ;
 wire result_sign_stage2;
 wire valid_stage1;
 wire valid_stage2;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;

 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1920_ (.A1(_1232_),
    .A2(_1322_),
    .A3(_1598_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1921_ (.A1(_1322_),
    .A2(_1598_),
    .B(_1325_),
    .C(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1922_ (.A1(_1321_),
    .A2(_1323_),
    .B(_1324_),
    .C(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1923_ (.A1(_1611_),
    .A2(_1567_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1924_ (.I(_1567_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1925_ (.A1(_1225_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1926_ (.A1(_1288_),
    .A2(_1315_),
    .B1(_1329_),
    .B2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1927_ (.A1(_1318_),
    .A2(_1319_),
    .B(_1605_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1928_ (.A1(_1232_),
    .A2(_1309_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _1929_ (.A1(_1321_),
    .A2(_1332_),
    .A3(_1333_),
    .A4(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1930_ (.A1(_1212_),
    .A2(_1223_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _1931_ (.A1(_1328_),
    .A2(_1335_),
    .A3(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1932_ (.I0(net3),
    .I1(net5),
    .I2(net35),
    .I3(net37),
    .S0(_1316_),
    .S1(_1337_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1933_ (.I(_1572_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1934_ (.I0(net35),
    .I1(net37),
    .S(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1935_ (.A1(_1229_),
    .A2(_1234_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1936_ (.A1(_1589_),
    .A2(_1341_),
    .B(_1581_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1937_ (.A1(_1611_),
    .A2(_1571_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1938_ (.A1(_1613_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1939_ (.I(_1607_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _1940_ (.A1(_1307_),
    .A2(_1344_),
    .B(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1941_ (.A1(_1237_),
    .A2(_1346_),
    .B(_1583_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1942_ (.A1(_1581_),
    .A2(_1236_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1943_ (.A1(_1230_),
    .A2(_1344_),
    .B(_1234_),
    .C(_1233_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1944_ (.A1(_1229_),
    .A2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1945_ (.A1(_1342_),
    .A2(_1347_),
    .B(_1348_),
    .C(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _1946_ (.A1(_1291_),
    .A2(_1292_),
    .A3(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1947_ (.A1(_1314_),
    .A2(_1338_),
    .B1(_1340_),
    .B2(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1948_ (.I0(net30),
    .I1(net32),
    .I2(net62),
    .I3(net64),
    .S0(_1316_),
    .S1(_1337_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1949_ (.I0(net62),
    .I1(net64),
    .S(_1339_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1950_ (.A1(_1314_),
    .A2(_1354_),
    .B1(_1355_),
    .B2(_1352_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1951_ (.A1(_1240_),
    .A2(_1246_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1952_ (.A1(_1263_),
    .A2(_1281_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1953_ (.A1(_1611_),
    .A2(_1330_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1954_ (.A1(_1225_),
    .A2(_1567_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _1955_ (.A1(_1357_),
    .A2(_1358_),
    .B1(_1359_),
    .B2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1956_ (.I(_1571_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1957_ (.A1(_1611_),
    .A2(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1958_ (.A1(_1225_),
    .A2(_1571_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1959_ (.A1(_1363_),
    .A2(_1364_),
    .B(_1291_),
    .C(_1292_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1960_ (.A1(_1361_),
    .A2(_1365_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1961_ (.I(_1366_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1962_ (.I0(_1353_),
    .I1(_1356_),
    .S(_1367_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1963_ (.A1(_1290_),
    .A2(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1964_ (.A1(_1318_),
    .A2(_1319_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1965_ (.I0(_1228_),
    .I1(_1370_),
    .S(_1283_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _1966_ (.A1(_1605_),
    .A2(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _1967_ (.I(_1283_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1968_ (.I0(_1309_),
    .I1(_1346_),
    .S(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _1969_ (.A1(_1232_),
    .A2(_1374_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _1970_ (.A1(_1372_),
    .A2(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1971_ (.A1(_1369_),
    .A2(_1376_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _1972_ (.I(_1572_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1973_ (.A1(_1225_),
    .A2(_1362_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1974_ (.A1(_1378_),
    .A2(_1291_),
    .A3(_1292_),
    .A4(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1975_ (.A1(_1378_),
    .A2(_1291_),
    .A3(_1292_),
    .A4(_1343_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _1976_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1329_),
    .B2(_1331_),
    .C(_1316_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _1977_ (.A1(_1380_),
    .A2(_1381_),
    .A3(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _1978_ (.A1(_1314_),
    .A2(_1352_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1979_ (.A1(_1298_),
    .A2(_1304_),
    .A3(_1312_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _1980_ (.A1(_1328_),
    .A2(_1335_),
    .A3(_1336_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1981_ (.A1(_1385_),
    .A2(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1982_ (.I(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1983_ (.I0(net16),
    .I1(_1204_),
    .S(_1288_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1984_ (.A1(_1284_),
    .A2(_1388_),
    .A3(_1389_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1985_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1986_ (.I0(_1679_),
    .I1(_1391_),
    .S(_1288_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1987_ (.A1(_1284_),
    .A2(_1388_),
    .B(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1988_ (.A1(_1390_),
    .A2(_1393_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1989_ (.A1(_1384_),
    .A2(_1394_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1990_ (.I(_1372_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _1991_ (.A1(_1232_),
    .A2(_1374_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1992_ (.A1(_1396_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1993_ (.A1(_1383_),
    .A2(_1395_),
    .A3(_1398_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1994_ (.I(_1690_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1995_ (.I(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1996_ (.I0(net43),
    .I1(net46),
    .S(_1315_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1997_ (.I0(net11),
    .I1(net14),
    .S(_1315_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1998_ (.A1(_1328_),
    .A2(_1335_),
    .A3(_1336_),
    .A4(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1999_ (.A1(_1386_),
    .A2(_1402_),
    .B(_1404_),
    .C(_1385_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2000_ (.I0(net43),
    .I1(net46),
    .S(_1339_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2001_ (.A1(_1351_),
    .A2(_1406_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2002_ (.I(_1373_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2003_ (.I0(_1405_),
    .I1(_1407_),
    .S(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2004_ (.I0(net7),
    .I1(net9),
    .S(_1315_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2005_ (.I0(net39),
    .I1(net41),
    .S(_1315_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2006_ (.I(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2007_ (.A1(_1328_),
    .A2(_1335_),
    .A3(_1336_),
    .B(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2008_ (.A1(_1337_),
    .A2(_1410_),
    .B(_1413_),
    .C(_1385_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2009_ (.I0(net39),
    .I1(net41),
    .S(_1339_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2010_ (.A1(_1351_),
    .A2(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2011_ (.I0(_1414_),
    .I1(_1416_),
    .S(_1408_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2012_ (.I0(_1409_),
    .I1(_1417_),
    .S(_1366_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2013_ (.A1(_1401_),
    .A2(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2014_ (.A1(_1378_),
    .A2(_1351_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2015_ (.I(_1315_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2016_ (.A1(_1421_),
    .A2(_1385_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2017_ (.I0(_1420_),
    .I1(_1422_),
    .S(_1283_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2018_ (.I(_1423_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2019_ (.A1(_1339_),
    .A2(_1351_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2020_ (.A1(_1315_),
    .A2(_1385_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2021_ (.I0(_1425_),
    .I1(_1426_),
    .S(_1283_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2022_ (.I(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2023_ (.A1(_1283_),
    .A2(_1388_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2024_ (.A1(net40),
    .A2(_1424_),
    .B1(_1428_),
    .B2(net42),
    .C(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2025_ (.I(_1373_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2026_ (.I(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2027_ (.A1(_1385_),
    .A2(_1386_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2028_ (.I(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2029_ (.I0(net8),
    .I1(net10),
    .S(_1316_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2030_ (.A1(_1432_),
    .A2(_1434_),
    .A3(_1435_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2031_ (.A1(_1366_),
    .A2(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2032_ (.A1(_1361_),
    .A2(_1365_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2033_ (.I(_1431_),
    .Z(a_exp_larger));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2034_ (.I(net12),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2035_ (.I(net15),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2036_ (.I0(_1439_),
    .I1(_1440_),
    .I2(_1667_),
    .I3(_1682_),
    .S0(_1315_),
    .S1(_1337_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2037_ (.I0(net44),
    .I1(net47),
    .S(_1339_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2038_ (.A1(_1291_),
    .A2(_1292_),
    .A3(_1351_),
    .A4(_1442_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2039_ (.A1(a_exp_larger),
    .A2(_1313_),
    .A3(_1441_),
    .B(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2040_ (.A1(_1438_),
    .A2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2041_ (.A1(_1430_),
    .A2(_1437_),
    .B(_1290_),
    .C(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2042_ (.A1(_1372_),
    .A2(_1375_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2043_ (.A1(_1419_),
    .A2(_1446_),
    .A3(_1447_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2044_ (.A1(_1377_),
    .A2(_1399_),
    .A3(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2045_ (.I(_1346_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2046_ (.A1(_1690_),
    .A2(_1378_),
    .B1(_1343_),
    .B2(_1379_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2047_ (.A1(_1307_),
    .A2(_1228_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2048_ (.A1(_1451_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2049_ (.A1(_1322_),
    .A2(_1601_),
    .B1(_1450_),
    .B2(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2050_ (.A1(_1605_),
    .A2(_1228_),
    .B(_1607_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2051_ (.A1(_1346_),
    .A2(_1453_),
    .B1(_1455_),
    .B2(_1593_),
    .C(_1232_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2052_ (.A1(_1232_),
    .A2(_1454_),
    .B(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2053_ (.I(_1601_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2054_ (.A1(_1458_),
    .A2(_1455_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2055_ (.I0(_1458_),
    .I1(_1459_),
    .S(_1593_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2056_ (.A1(_1352_),
    .A2(_1457_),
    .A3(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2057_ (.A1(_1408_),
    .A2(_1313_),
    .A3(_1328_),
    .A4(_1335_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2058_ (.A1(_1461_),
    .A2(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2059_ (.A1(_1212_),
    .A2(_1432_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2060_ (.A1(_1223_),
    .A2(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2061_ (.A1(_1463_),
    .A2(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2062_ (.I(_1438_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2063_ (.I(net4),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2064_ (.I(_1433_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2065_ (.A1(_1468_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2066_ (.I(_1433_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2067_ (.A1(_1408_),
    .A2(_1471_),
    .B(net36),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2068_ (.A1(_1378_),
    .A2(_1247_),
    .A3(_1282_),
    .A4(_1351_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2069_ (.A1(_1283_),
    .A2(_1422_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2070_ (.A1(_1470_),
    .A2(_1472_),
    .B(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2071_ (.I(net6),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2072_ (.A1(_1476_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2073_ (.A1(_1408_),
    .A2(_1471_),
    .B(net38),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2074_ (.A1(_1339_),
    .A2(_1247_),
    .A3(_1282_),
    .A4(_1351_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2075_ (.A1(_1283_),
    .A2(_1426_),
    .B(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2076_ (.A1(_1477_),
    .A2(_1478_),
    .B(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2077_ (.A1(_1475_),
    .A2(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2078_ (.I(net31),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2079_ (.A1(_1483_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2080_ (.A1(_1432_),
    .A2(_1471_),
    .B(net63),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2081_ (.A1(_1484_),
    .A2(_1485_),
    .B(_1474_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2082_ (.I(net33),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2083_ (.A1(_1487_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2084_ (.A1(_1432_),
    .A2(_1471_),
    .B(net65),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2085_ (.A1(_1488_),
    .A2(_1489_),
    .B(_1480_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2086_ (.A1(_1467_),
    .A2(_1486_),
    .A3(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2087_ (.A1(_1467_),
    .A2(_1482_),
    .B(_1491_),
    .C(_1401_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _2088_ (.I(_1372_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2089_ (.I(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2090_ (.A1(_1397_),
    .A2(_1463_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2091_ (.A1(_1494_),
    .A2(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2092_ (.A1(_1396_),
    .A2(_1495_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2093_ (.I(_1367_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2094_ (.A1(_1283_),
    .A2(_1387_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2095_ (.I0(net24),
    .I1(net56),
    .S(_1499_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2096_ (.I0(net28),
    .I1(net60),
    .S(_1499_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2097_ (.A1(_1424_),
    .A2(_1500_),
    .B1(_1501_),
    .B2(_1428_),
    .C(_1290_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2098_ (.I0(net27),
    .I1(net59),
    .S(_1499_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _2099_ (.I0(net29),
    .I1(net61),
    .S(_1499_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2100_ (.A1(_1424_),
    .A2(_1503_),
    .B1(_1504_),
    .B2(_1428_),
    .C(_1401_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2101_ (.I(_1288_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2102_ (.A1(net45),
    .A2(_1506_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2103_ (.A1(net34),
    .A2(_1400_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2104_ (.A1(a_exp_larger),
    .A2(_1434_),
    .B1(_1507_),
    .B2(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2105_ (.A1(net13),
    .A2(_1506_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2106_ (.A1(net2),
    .A2(_1400_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _2107_ (.A1(_1510_),
    .A2(_1511_),
    .B(_1284_),
    .C(_1388_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2108_ (.A1(_1509_),
    .A2(_1512_),
    .B(_1480_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2109_ (.A1(_1498_),
    .A2(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2110_ (.A1(_1498_),
    .A2(_1502_),
    .A3(_1505_),
    .B(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2111_ (.A1(_1492_),
    .A2(_1496_),
    .B1(_1497_),
    .B2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2112_ (.I(_1465_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2113_ (.A1(_1449_),
    .A2(_1466_),
    .B1(_1516_),
    .B2(_1517_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2114_ (.I0(net30),
    .I1(net62),
    .S(_1499_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _2115_ (.A1(_1424_),
    .A2(_1501_),
    .B1(_1518_),
    .B2(_1428_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2116_ (.A1(_1424_),
    .A2(_1503_),
    .B1(_1504_),
    .B2(_1428_),
    .C(_1290_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2117_ (.A1(_1290_),
    .A2(_1519_),
    .B(_1520_),
    .C(_1498_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _2118_ (.I0(_1316_),
    .I1(_1339_),
    .S(_1408_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2119_ (.I(_1499_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2120_ (.I0(net13),
    .I1(net24),
    .I2(net45),
    .I3(net56),
    .S0(_1506_),
    .S1(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2121_ (.A1(_1384_),
    .A2(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2122_ (.A1(_1522_),
    .A2(_1525_),
    .B(_1467_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2123_ (.I0(net2),
    .I1(net34),
    .S(_1523_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2124_ (.A1(_1506_),
    .A2(_1384_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2125_ (.A1(_1527_),
    .A2(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2126_ (.A1(_1383_),
    .A2(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2127_ (.A1(_1396_),
    .A2(_1397_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _2128_ (.A1(_1521_),
    .A2(_1526_),
    .B(_1530_),
    .C(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2129_ (.A1(net16),
    .A2(_1284_),
    .A3(_1388_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2130_ (.A1(_1284_),
    .A2(_1388_),
    .B(_1679_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2131_ (.A1(_1533_),
    .A2(_1534_),
    .B(_1522_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2132_ (.I(net14),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2133_ (.A1(_1536_),
    .A2(_1316_),
    .A3(_1408_),
    .A4(_1469_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2134_ (.A1(_1378_),
    .A2(_1291_),
    .A3(_1292_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2135_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1385_),
    .B2(_1386_),
    .C(_1316_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2136_ (.A1(_1538_),
    .A2(_1539_),
    .B(net46),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2137_ (.A1(_1537_),
    .A2(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2138_ (.A1(_1535_),
    .A2(_1541_),
    .B(_1498_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2139_ (.I(net9),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2140_ (.I(net11),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2141_ (.I0(_1543_),
    .I1(_1544_),
    .S(_1316_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2142_ (.A1(_1432_),
    .A2(_1471_),
    .A3(_1545_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2143_ (.A1(net41),
    .A2(_1421_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2144_ (.A1(net43),
    .A2(_1316_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2145_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1547_),
    .B2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2146_ (.A1(net41),
    .A2(_1378_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2147_ (.A1(net43),
    .A2(_1339_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2148_ (.A1(_1550_),
    .A2(_1551_),
    .B(_1357_),
    .C(_1358_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2149_ (.A1(a_exp_larger),
    .A2(_1434_),
    .B1(_1549_),
    .B2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2150_ (.A1(_1546_),
    .A2(_1553_),
    .B(_1467_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2151_ (.A1(_1542_),
    .A2(_1554_),
    .B(_1447_),
    .C(_1528_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2152_ (.A1(_1204_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2153_ (.A1(_1408_),
    .A2(_1471_),
    .B(_1391_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2154_ (.A1(_1400_),
    .A2(_1384_),
    .A3(_1556_),
    .A4(_1557_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2155_ (.A1(_1383_),
    .A2(_1558_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2156_ (.A1(_1401_),
    .A2(_1372_),
    .A3(_1375_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2157_ (.A1(_1430_),
    .A2(_1437_),
    .B(_1445_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2158_ (.A1(_1398_),
    .A2(_1559_),
    .B1(_1560_),
    .B2(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2159_ (.A1(_1372_),
    .A2(_1375_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2160_ (.I(net3),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2161_ (.A1(_1564_),
    .A2(_1408_),
    .A3(_1469_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2162_ (.A1(_1432_),
    .A2(_1434_),
    .B(net35),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2163_ (.A1(_0122_),
    .A2(_0123_),
    .B(_1480_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2164_ (.I(net32),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2165_ (.A1(_0125_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2166_ (.A1(_1432_),
    .A2(_1434_),
    .B(net64),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2167_ (.A1(_0126_),
    .A2(_0127_),
    .B(_1474_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2168_ (.A1(_1289_),
    .A2(_1366_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2169_ (.A1(_1506_),
    .A2(_1438_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2170_ (.I(net7),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2171_ (.A1(_0131_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2172_ (.A1(_1432_),
    .A2(_1471_),
    .B(net39),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2173_ (.A1(_0132_),
    .A2(_0133_),
    .B(_1480_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2174_ (.I(net5),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2175_ (.A1(_0135_),
    .A2(_1431_),
    .A3(_1469_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2176_ (.A1(_1432_),
    .A2(_1471_),
    .B(net37),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2177_ (.A1(_0136_),
    .A2(_0137_),
    .B(_1474_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _2178_ (.A1(_0124_),
    .A2(_0128_),
    .A3(_0129_),
    .B1(_0130_),
    .B2(_0134_),
    .B3(_0138_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2179_ (.A1(_1400_),
    .A2(_1366_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2180_ (.A1(_1400_),
    .A2(_1438_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _2181_ (.A1(_0140_),
    .A2(_1486_),
    .A3(_1490_),
    .B1(_0141_),
    .B2(_1481_),
    .B3(_1475_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2182_ (.A1(_1563_),
    .A2(_0139_),
    .A3(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2183_ (.A1(_1555_),
    .A2(_1562_),
    .A3(_0143_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2184_ (.A1(_1532_),
    .A2(_0144_),
    .B(_1466_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2185_ (.A1(_1484_),
    .A2(_1485_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _2186_ (.A1(_1424_),
    .A2(_1504_),
    .B1(_0145_),
    .B2(_1428_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2187_ (.A1(_1509_),
    .A2(_1512_),
    .B(_1522_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2188_ (.A1(net59),
    .A2(_1506_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2189_ (.A1(net56),
    .A2(_1400_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2190_ (.A1(a_exp_larger),
    .A2(_1434_),
    .B1(_0148_),
    .B2(_0149_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2191_ (.A1(net27),
    .A2(_1506_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2192_ (.A1(net24),
    .A2(_1400_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2193_ (.A1(_0151_),
    .A2(_0152_),
    .B(_1284_),
    .C(_1388_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _2194_ (.I0(_1421_),
    .I1(_1378_),
    .S(a_exp_larger),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2195_ (.A1(_0150_),
    .A2(_0153_),
    .B(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2196_ (.A1(_0147_),
    .A2(_0155_),
    .B(_1498_),
    .C(_1384_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2197_ (.A1(_1519_),
    .A2(_0141_),
    .B1(_0146_),
    .B2(_0130_),
    .C(_0156_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2198_ (.A1(_0124_),
    .A2(_0128_),
    .B(_1401_),
    .C(_1367_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2199_ (.A1(_1400_),
    .A2(_1438_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2200_ (.A1(_0134_),
    .A2(_0138_),
    .B(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2201_ (.I(_1438_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2202_ (.A1(_1488_),
    .A2(_1489_),
    .B(_1474_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2203_ (.A1(_1470_),
    .A2(_1472_),
    .B(_1480_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2204_ (.I0(net6),
    .I1(net8),
    .I2(net38),
    .I3(net40),
    .S0(_1315_),
    .S1(_1337_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2205_ (.I0(net38),
    .I1(net40),
    .S(_1339_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _2206_ (.A1(_1314_),
    .A2(_0164_),
    .B1(_0165_),
    .B2(_1352_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2207_ (.A1(_1438_),
    .A2(_0166_),
    .B(_1400_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2208_ (.A1(_0161_),
    .A2(_0162_),
    .A3(_0163_),
    .B(_0167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2209_ (.A1(_0158_),
    .A2(_0160_),
    .A3(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2210_ (.A1(_1531_),
    .A2(_0157_),
    .B1(_0169_),
    .B2(_1376_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2211_ (.I0(_1440_),
    .I1(_1536_),
    .I2(_1682_),
    .I3(_1685_),
    .S0(_1690_),
    .S1(_1523_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2212_ (.A1(_1390_),
    .A2(_1393_),
    .B(_1522_),
    .C(_1384_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2213_ (.A1(_1474_),
    .A2(_0171_),
    .B(_0172_),
    .C(_0161_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2214_ (.A1(net44),
    .A2(_1506_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2215_ (.A1(net43),
    .A2(_1690_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2216_ (.A1(_1284_),
    .A2(_1388_),
    .B1(_0174_),
    .B2(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2217_ (.A1(net12),
    .A2(_1506_),
    .A3(_1284_),
    .A4(_1388_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2218_ (.A1(net11),
    .A2(_1690_),
    .A3(_1284_),
    .A4(_1388_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2219_ (.A1(_0176_),
    .A2(_0177_),
    .A3(_0178_),
    .B(_1428_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2220_ (.A1(_1367_),
    .A2(_0179_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2221_ (.I(net10),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2222_ (.I0(_0181_),
    .I1(_1543_),
    .I2(_1673_),
    .I3(_1676_),
    .S0(_1690_),
    .S1(_1523_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2223_ (.A1(_1383_),
    .A2(_1384_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2224_ (.A1(_0182_),
    .A2(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2225_ (.A1(_0173_),
    .A2(_0180_),
    .B(_0184_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _2226_ (.A1(_1494_),
    .A2(_1397_),
    .A3(_1466_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2227_ (.A1(net34),
    .A2(_1287_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2228_ (.A1(_1466_),
    .A2(_0170_),
    .B1(_0185_),
    .B2(_0186_),
    .C(_0187_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2229_ (.I0(net27),
    .I1(net28),
    .I2(net59),
    .I3(net60),
    .S0(_1506_),
    .S1(_1523_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2230_ (.A1(_1424_),
    .A2(_1524_),
    .B1(_0188_),
    .B2(_1428_),
    .C(_1467_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2231_ (.A1(_1290_),
    .A2(_1467_),
    .A3(_1356_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2232_ (.A1(_0159_),
    .A2(_0146_),
    .B(_0189_),
    .C(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2233_ (.I0(_1353_),
    .I1(_1417_),
    .S(_0161_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2234_ (.A1(_0161_),
    .A2(_0166_),
    .B(_1289_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2235_ (.A1(_1467_),
    .A2(_0162_),
    .A3(_0163_),
    .B(_0193_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2236_ (.A1(_1401_),
    .A2(_0192_),
    .B(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2237_ (.A1(_1531_),
    .A2(_0191_),
    .B1(_0195_),
    .B2(_1376_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2238_ (.I0(net15),
    .I1(net16),
    .I2(net47),
    .I3(net48),
    .S0(_1288_),
    .S1(_1523_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2239_ (.A1(_1522_),
    .A2(_1558_),
    .B1(_0197_),
    .B2(_1424_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2240_ (.A1(_1439_),
    .A2(_1432_),
    .A3(_1471_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2241_ (.A1(a_exp_larger),
    .A2(_1434_),
    .B(net44),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2242_ (.A1(_0199_),
    .A2(_0200_),
    .B(_1480_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2243_ (.A1(_0181_),
    .A2(_1408_),
    .A3(_1471_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2244_ (.A1(a_exp_larger),
    .A2(_1434_),
    .B(net42),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2245_ (.A1(_0202_),
    .A2(_0203_),
    .B(_1474_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2246_ (.A1(_1289_),
    .A2(_1409_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2247_ (.A1(_1289_),
    .A2(_0201_),
    .A3(_0204_),
    .B(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _2248_ (.I0(_0198_),
    .I1(_0206_),
    .S(_1367_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2249_ (.A1(net45),
    .A2(_1287_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2250_ (.A1(_1466_),
    .A2(_0196_),
    .B1(_0207_),
    .B2(_0186_),
    .C(_0208_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2251_ (.A1(_1212_),
    .A2(_1285_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2252_ (.I(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2253_ (.A1(_1465_),
    .A2(_1495_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2254_ (.I(_0211_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2255_ (.A1(_1424_),
    .A2(_1500_),
    .B1(_1501_),
    .B2(_1428_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2256_ (.A1(_1486_),
    .A2(_1490_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2257_ (.A1(_1424_),
    .A2(_1503_),
    .B1(_1504_),
    .B2(_1428_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2258_ (.I0(_1356_),
    .I1(_0213_),
    .I2(_0214_),
    .I3(_0215_),
    .S0(_1367_),
    .S1(_1290_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _2259_ (.A1(_1643_),
    .A2(_1474_),
    .B1(_1480_),
    .B2(_1673_),
    .C(_1523_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2260_ (.A1(_0217_),
    .A2(_1436_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2261_ (.I0(_1353_),
    .I1(_1417_),
    .I2(_1482_),
    .I3(_0218_),
    .S0(_0161_),
    .S1(_1289_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2262_ (.I0(_0216_),
    .I1(_0219_),
    .S(_1493_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2263_ (.A1(_1438_),
    .A2(_0154_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2264_ (.A1(_1289_),
    .A2(_1444_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2265_ (.A1(_1289_),
    .A2(_1409_),
    .B(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _2266_ (.A1(_1395_),
    .A2(_0221_),
    .B1(_0223_),
    .B2(_1498_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _2267_ (.A1(_1628_),
    .A2(_0210_),
    .B1(_0212_),
    .B2(_0220_),
    .C1(_0224_),
    .C2(_0186_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2268_ (.I(net16),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2269_ (.A1(_0225_),
    .A2(a_exp_larger),
    .A3(_1434_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2270_ (.A1(a_exp_larger),
    .A2(_1434_),
    .B(net48),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2271_ (.A1(_0226_),
    .A2(_0227_),
    .B(_0154_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2272_ (.A1(_1537_),
    .A2(_1540_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2273_ (.A1(_0228_),
    .A2(_0229_),
    .B(_1528_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2274_ (.A1(_1401_),
    .A2(_1444_),
    .B(_1467_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2275_ (.A1(_0230_),
    .A2(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2276_ (.A1(_0154_),
    .A2(_1558_),
    .B(_1498_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2277_ (.A1(_0232_),
    .A2(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2278_ (.I0(_0215_),
    .I1(_0214_),
    .S(_0161_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2279_ (.I0(_0218_),
    .I1(_1482_),
    .S(_1367_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2280_ (.A1(_0124_),
    .A2(_0128_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2281_ (.I0(_1519_),
    .I1(_0237_),
    .S(_1438_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2282_ (.A1(_0134_),
    .A2(_0138_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2283_ (.A1(_1314_),
    .A2(_1352_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2284_ (.A1(_1546_),
    .A2(_1553_),
    .B(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2285_ (.A1(_0161_),
    .A2(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2286_ (.A1(_1498_),
    .A2(_0239_),
    .B(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _2287_ (.I0(_0235_),
    .I1(_0236_),
    .I2(_0238_),
    .I3(_0243_),
    .S0(_1493_),
    .S1(_1290_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2288_ (.A1(net59),
    .A2(_1287_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2289_ (.A1(_0186_),
    .A2(_0234_),
    .B1(_0244_),
    .B2(_0212_),
    .C(_0245_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2290_ (.A1(_1474_),
    .A2(_0182_),
    .B(_0179_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2291_ (.A1(_1289_),
    .A2(_0134_),
    .A3(_0138_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2292_ (.A1(_1289_),
    .A2(_0166_),
    .B(_0161_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2293_ (.A1(_1467_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2294_ (.A1(_0162_),
    .A2(_0163_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2295_ (.I0(_1519_),
    .I1(_0237_),
    .I2(_0146_),
    .I3(_0250_),
    .S0(_0161_),
    .S1(_1290_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2296_ (.I0(_0249_),
    .I1(_0251_),
    .S(_1396_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2297_ (.A1(_1474_),
    .A2(_0171_),
    .B(_0172_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2298_ (.A1(_1498_),
    .A2(_0253_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _2299_ (.A1(_1640_),
    .A2(_0210_),
    .B1(_0211_),
    .B2(_0252_),
    .C1(_0254_),
    .C2(_0186_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2300_ (.A1(_1366_),
    .A2(_0166_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2301_ (.A1(_1367_),
    .A2(_0201_),
    .A3(_0204_),
    .B(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2302_ (.I0(_1418_),
    .I1(_0256_),
    .S(_1401_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2303_ (.I0(_1353_),
    .I1(_1356_),
    .I2(_0250_),
    .I3(_0146_),
    .S0(_1367_),
    .S1(_1401_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2304_ (.I0(_0257_),
    .I1(_0258_),
    .S(_1396_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _2305_ (.A1(_1467_),
    .A2(_0198_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _2306_ (.A1(_1637_),
    .A2(_0210_),
    .B1(_0211_),
    .B2(_0259_),
    .C1(_0260_),
    .C2(_0186_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _2307_ (.A1(_1390_),
    .A2(_1393_),
    .B(_1383_),
    .C(_1384_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2308_ (.A1(_1375_),
    .A2(_0261_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2309_ (.A1(_1369_),
    .A2(_1375_),
    .A3(_1492_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2310_ (.A1(_1419_),
    .A2(_1446_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2311_ (.A1(_1563_),
    .A2(_1466_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2312_ (.A1(net62),
    .A2(_1287_),
    .B1(_0264_),
    .B2(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2313_ (.A1(_1494_),
    .A2(_1466_),
    .A3(_0263_),
    .B(_0266_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2314_ (.A1(_1383_),
    .A2(_1558_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2315_ (.A1(_0139_),
    .A2(_0142_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2316_ (.A1(_1535_),
    .A2(_1541_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2317_ (.A1(_1438_),
    .A2(_1528_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2318_ (.A1(_1429_),
    .A2(_1549_),
    .A3(_1552_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2319_ (.A1(_1543_),
    .A2(_1421_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2320_ (.A1(_1544_),
    .A2(_1316_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2321_ (.A1(_0272_),
    .A2(_0273_),
    .B(_1429_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2322_ (.A1(_1367_),
    .A2(_1528_),
    .A3(_0271_),
    .A4(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2323_ (.A1(_1401_),
    .A2(_1561_),
    .B1(_0269_),
    .B2(_0270_),
    .C(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2324_ (.I0(_0268_),
    .I1(_0276_),
    .S(_1493_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _2325_ (.A1(_1631_),
    .A2(_0210_),
    .B1(_0267_),
    .B2(_0186_),
    .C1(_0211_),
    .C2(_0277_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2326_ (.I(_0209_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2327_ (.A1(_0158_),
    .A2(_0160_),
    .A3(_0168_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2328_ (.I0(_0279_),
    .I1(_0185_),
    .S(_1494_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2329_ (.A1(_1664_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0280_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2330_ (.A1(_1494_),
    .A2(_0207_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2331_ (.A1(_1494_),
    .A2(_0195_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2332_ (.A1(_0212_),
    .A2(_0281_),
    .A3(_0282_),
    .B1(_0210_),
    .B2(_1661_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2333_ (.I0(_0219_),
    .I1(_0224_),
    .S(_1494_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2334_ (.A1(_1658_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0283_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2335_ (.A1(_0230_),
    .A2(_0231_),
    .B(_0233_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2336_ (.A1(_1475_),
    .A2(_1481_),
    .B(_1498_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2337_ (.A1(_0161_),
    .A2(_1436_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2338_ (.A1(_0217_),
    .A2(_0286_),
    .B(_1290_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2339_ (.A1(_0134_),
    .A2(_0138_),
    .A3(_0129_),
    .B1(_0130_),
    .B2(_0241_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2340_ (.A1(_0285_),
    .A2(_0287_),
    .B(_0288_),
    .C(_1493_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2341_ (.A1(_1494_),
    .A2(_0284_),
    .B(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2342_ (.A1(_1655_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0290_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2343_ (.I0(_0249_),
    .I1(_0254_),
    .S(_1494_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2344_ (.A1(_1652_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0291_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2345_ (.I0(_0257_),
    .I1(_0260_),
    .S(_1494_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2346_ (.A1(_1649_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0292_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2347_ (.A1(_1396_),
    .A2(_0261_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2348_ (.A1(_1396_),
    .A2(_0264_),
    .B(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2349_ (.A1(_1646_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0294_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2350_ (.I0(_0267_),
    .I1(_0276_),
    .S(_1396_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2351_ (.A1(_1643_),
    .A2(_0278_),
    .B1(_0212_),
    .B2(_0295_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2352_ (.A1(_1465_),
    .A2(_1497_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2353_ (.A1(_1676_),
    .A2(_0278_),
    .B1(_0296_),
    .B2(_0185_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2354_ (.A1(_1673_),
    .A2(_0278_),
    .B1(_0296_),
    .B2(_0207_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2355_ (.A1(_1670_),
    .A2(_0278_),
    .B1(_0296_),
    .B2(_0224_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2356_ (.A1(_1667_),
    .A2(_0210_),
    .B1(_0296_),
    .B2(_0234_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2357_ (.A1(_1685_),
    .A2(_0210_),
    .B1(_0296_),
    .B2(_0254_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2358_ (.A1(_1682_),
    .A2(_0210_),
    .B1(_0296_),
    .B2(_0260_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2359_ (.A1(_1679_),
    .A2(_0210_),
    .B1(_0261_),
    .B2(_0296_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2360_ (.A1(_1497_),
    .A2(_1559_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2361_ (.A1(_1220_),
    .A2(_1221_),
    .A3(_1222_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2362_ (.A1(_0298_),
    .A2(_1464_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2363_ (.A1(_1464_),
    .A2(_0297_),
    .B1(_0299_),
    .B2(_1391_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2364_ (.A1(_1377_),
    .A2(_1399_),
    .A3(_1448_),
    .B(_1463_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2365_ (.I(_1212_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2366_ (.A1(_0301_),
    .A2(_1285_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2367_ (.A1(_1516_),
    .A2(_0300_),
    .B(_0302_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2368_ (.A1(_1532_),
    .A2(_0144_),
    .B(_1523_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2369_ (.A1(net2),
    .A2(_0209_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2370_ (.A1(_1429_),
    .A2(_1447_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2371_ (.A1(_0185_),
    .A2(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2372_ (.A1(_1523_),
    .A2(_0170_),
    .B(_0303_),
    .C(_0305_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2373_ (.A1(net13),
    .A2(_0209_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2374_ (.A1(_0207_),
    .A2(_0304_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2375_ (.A1(_1523_),
    .A2(_0196_),
    .B(_0306_),
    .C(_0307_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2376_ (.A1(_1397_),
    .A2(_1429_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2377_ (.I(_0308_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2378_ (.A1(net24),
    .A2(_1285_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2379_ (.A1(_0224_),
    .A2(_0304_),
    .B1(_0309_),
    .B2(_0220_),
    .C(_0310_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2380_ (.I(_1495_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2381_ (.A1(_1429_),
    .A2(_1447_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2382_ (.A1(net27),
    .A2(_1285_),
    .B1(_0284_),
    .B2(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2383_ (.A1(_0302_),
    .A2(_0311_),
    .A3(_0244_),
    .B(_0313_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2384_ (.A1(net28),
    .A2(_1285_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2385_ (.A1(_0254_),
    .A2(_0304_),
    .B1(_0309_),
    .B2(_0252_),
    .C(_0314_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2386_ (.A1(net29),
    .A2(_1285_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2387_ (.A1(_0260_),
    .A2(_0304_),
    .B1(_0309_),
    .B2(_0259_),
    .C(_0315_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2388_ (.A1(net30),
    .A2(_0210_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2389_ (.A1(_1396_),
    .A2(_1429_),
    .A3(_0262_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2390_ (.A1(_1369_),
    .A2(_1375_),
    .A3(_1492_),
    .B(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2391_ (.A1(_1429_),
    .A2(_0264_),
    .A3(_1376_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2392_ (.A1(_0316_),
    .A2(_0318_),
    .A3(_0319_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _2393_ (.A1(_1483_),
    .A2(_1287_),
    .B1(_0267_),
    .B2(_0304_),
    .C1(_0308_),
    .C2(_0277_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2394_ (.I(_1286_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2395_ (.A1(_0125_),
    .A2(_0320_),
    .B1(_0280_),
    .B2(_0309_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2396_ (.A1(_0281_),
    .A2(_0282_),
    .A3(_0308_),
    .B1(_1287_),
    .B2(_1487_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2397_ (.A1(_1564_),
    .A2(_0320_),
    .B1(_0283_),
    .B2(_0309_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2398_ (.A1(_1468_),
    .A2(_0320_),
    .B1(_0290_),
    .B2(_0309_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2399_ (.A1(_0135_),
    .A2(_0320_),
    .B1(_0291_),
    .B2(_0309_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2400_ (.A1(_1476_),
    .A2(_0320_),
    .B1(_0292_),
    .B2(_0309_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2401_ (.A1(_0131_),
    .A2(_0320_),
    .B1(_0294_),
    .B2(_0309_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2402_ (.A1(net8),
    .A2(_0209_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2403_ (.A1(_0295_),
    .A2(_0309_),
    .B(_0321_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2404_ (.A1(net9),
    .A2(_1285_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2405_ (.A1(_1396_),
    .A2(_1495_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2406_ (.A1(_1285_),
    .A2(_0323_),
    .A3(_0185_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2407_ (.A1(_0322_),
    .A2(_0324_),
    .B(_0301_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _2408_ (.A1(_0302_),
    .A2(_0323_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2409_ (.A1(_0181_),
    .A2(_0320_),
    .B1(_0207_),
    .B2(_0325_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2410_ (.A1(_1544_),
    .A2(_0320_),
    .B1(_0224_),
    .B2(_0325_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2411_ (.A1(_1439_),
    .A2(_0320_),
    .B1(_0234_),
    .B2(_0325_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2412_ (.A1(_1536_),
    .A2(_0320_),
    .B1(_0254_),
    .B2(_0325_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2413_ (.A1(_1440_),
    .A2(_1287_),
    .B1(_0260_),
    .B2(_0325_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2414_ (.A1(_0225_),
    .A2(_1287_),
    .B1(_0261_),
    .B2(_0325_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2415_ (.A1(_1204_),
    .A2(_1285_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2416_ (.A1(_0267_),
    .A2(_0325_),
    .B(_0326_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2417_ (.I(\add_result[26] ),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2418_ (.I(\add_result[25] ),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2419_ (.A1(\add_result[15] ),
    .A2(\add_result[18] ),
    .A3(\add_result[17] ),
    .A4(\add_result[19] ),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2420_ (.A1(\add_result[4] ),
    .A2(\add_result[24] ),
    .A3(_0328_),
    .A4(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2421_ (.I(\add_result[20] ),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2422_ (.I(\add_result[21] ),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2423_ (.I(\add_result[22] ),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _2424_ (.I(\add_result[23] ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2425_ (.A1(_0333_),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2426_ (.A1(\add_result[6] ),
    .A2(\add_result[5] ),
    .A3(\add_result[8] ),
    .A4(\add_result[14] ),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2427_ (.A1(_0331_),
    .A2(_0332_),
    .A3(_0335_),
    .A4(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2428_ (.A1(\add_result[7] ),
    .A2(\add_result[10] ),
    .A3(\add_result[9] ),
    .A4(\add_result[12] ),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2429_ (.A1(\add_result[3] ),
    .A2(\add_result[11] ),
    .A3(\add_result[13] ),
    .A4(\add_result[16] ),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2430_ (.A1(_0338_),
    .A2(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2431_ (.A1(_0327_),
    .A2(_0330_),
    .A3(_0337_),
    .A4(_0340_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2432_ (.A1(inexact_stage2),
    .A2(_0341_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _2433_ (.I(\add_result[25] ),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _2434_ (.I(\add_result[26] ),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2435_ (.A1(_0342_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _2436_ (.A1(\add_result[24] ),
    .A2(_0335_),
    .A3(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _2437_ (.I(_0345_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2438_ (.I(\add_result[24] ),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2439_ (.A1(_0342_),
    .A2(_0343_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2440_ (.A1(_0331_),
    .A2(_0332_),
    .B(_0334_),
    .C(_0333_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2441_ (.A1(_0346_),
    .A2(_0347_),
    .A3(_0348_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2442_ (.I(\add_result[21] ),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2443_ (.A1(\add_result[20] ),
    .A2(_0349_),
    .B(\add_result[22] ),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2444_ (.A1(\add_result[23] ),
    .A2(_0350_),
    .B(_0346_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2445_ (.A1(_0347_),
    .A2(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2446_ (.I(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2447_ (.I(_0353_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2448_ (.A1(_0330_),
    .A2(_0337_),
    .A3(_0340_),
    .B(_0343_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2449_ (.I(_1710_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2450_ (.A1(_0355_),
    .A2(_1712_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2451_ (.A1(_1704_),
    .A2(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2452_ (.A1(_1703_),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2453_ (.A1(_1697_),
    .A2(_0358_),
    .B(_1696_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2454_ (.A1(\result_exp_stage2[5] ),
    .A2(\result_exp_stage2[4] ),
    .A3(\result_exp_stage2[3] ),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2455_ (.A1(\result_exp_stage2[6] ),
    .A2(_0360_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2456_ (.A1(\result_exp_stage2[7] ),
    .A2(_0359_),
    .A3(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2457_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2458_ (.A1(_0328_),
    .A2(_0354_),
    .A3(_0363_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2459_ (.I(\result_exp_stage2[0] ),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2460_ (.I(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2461_ (.I(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2462_ (.I(_0366_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2463_ (.I(\result_exp_stage2[1] ),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2464_ (.I(\result_exp_stage2[2] ),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2465_ (.I(_1709_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2466_ (.A1(net22),
    .A2(net21),
    .A3(net25),
    .A4(net23),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2467_ (.A1(net18),
    .A2(net17),
    .A3(net20),
    .A4(net19),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2468_ (.A1(_0367_),
    .A2(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2469_ (.A1(net54),
    .A2(net53),
    .A3(net57),
    .A4(net55),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2470_ (.A1(net50),
    .A2(net49),
    .A3(net52),
    .A4(net51),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2471_ (.A1(_0370_),
    .A2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2472_ (.A1(_0369_),
    .A2(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2473_ (.I(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2474_ (.I(\aligned_a_mant[0] ),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2475_ (.I(\aligned_b_mant[0] ),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2476_ (.I(_1734_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2477_ (.A1(_0375_),
    .A2(_0376_),
    .A3(_1730_),
    .B(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2478_ (.I(is_a_larger_stage1),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2479_ (.I0(_1729_),
    .I1(_1732_),
    .S(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2480_ (.A1(_0375_),
    .A2(\aligned_b_mant[0] ),
    .A3(_1729_),
    .A4(is_a_larger_stage1),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2481_ (.I(is_a_larger_stage1),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2482_ (.I(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2483_ (.I(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2484_ (.A1(\aligned_a_mant[0] ),
    .A2(_0376_),
    .A3(_1732_),
    .A4(_0384_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2485_ (.A1(_1730_),
    .A2(_0380_),
    .B(_0381_),
    .C(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _2486_ (.A1(a_sign_stage1),
    .A2(b_sign_stage1),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2487_ (.I(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2488_ (.I0(_0378_),
    .I1(_0386_),
    .S(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2489_ (.A1(_1722_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2490_ (.A1(_0374_),
    .A2(_0390_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2491_ (.A1(a_sign_stage1),
    .A2(b_sign_stage1),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2492_ (.I(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2493_ (.I(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2494_ (.I(_1722_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2495_ (.A1(_0394_),
    .A2(_0378_),
    .B(_1726_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2496_ (.I(_0387_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2497_ (.I(_1732_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2498_ (.A1(\aligned_a_mant[0] ),
    .A2(_0376_),
    .B(_1730_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2499_ (.A1(_0397_),
    .A2(_0398_),
    .B(_0394_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2500_ (.A1(_0384_),
    .A2(_1724_),
    .A3(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2501_ (.I(_1729_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2502_ (.A1(_0375_),
    .A2(\aligned_b_mant[0] ),
    .B(_1730_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2503_ (.A1(_0401_),
    .A2(_0402_),
    .B(_0394_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2504_ (.A1(_0379_),
    .A2(_1721_),
    .A3(_0403_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2505_ (.A1(_0396_),
    .A2(_0400_),
    .A3(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2506_ (.A1(_0393_),
    .A2(_0395_),
    .B(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2507_ (.A1(_1738_),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2508_ (.A1(_0374_),
    .A2(_0407_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2509_ (.I(_1742_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2510_ (.A1(_1738_),
    .A2(_0395_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2511_ (.I(_1740_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2512_ (.A1(_1724_),
    .A2(_0399_),
    .B(_1738_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2513_ (.A1(_0410_),
    .A2(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2514_ (.I(_1737_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2515_ (.A1(_1721_),
    .A2(_0403_),
    .B(_1738_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2516_ (.A1(_0413_),
    .A2(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2517_ (.I(_0384_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2518_ (.I0(_0412_),
    .I1(_0415_),
    .S(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2519_ (.I0(_0409_),
    .I1(_0417_),
    .S(_0388_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2520_ (.A1(_1746_),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2521_ (.A1(_0374_),
    .A2(_0419_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2522_ (.I(_1746_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2523_ (.A1(_0420_),
    .A2(_0409_),
    .B(_1750_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2524_ (.I(_1748_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2525_ (.A1(_0420_),
    .A2(_0412_),
    .B(_0422_),
    .C(_0379_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2526_ (.I(_1745_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2527_ (.A1(_0420_),
    .A2(_0415_),
    .B(_0424_),
    .C(_0416_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2528_ (.A1(_0396_),
    .A2(_0423_),
    .A3(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2529_ (.A1(_0393_),
    .A2(_0421_),
    .B(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2530_ (.A1(_1754_),
    .A2(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2531_ (.A1(_0374_),
    .A2(_0428_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2532_ (.I(_1762_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2533_ (.I(_1730_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2534_ (.A1(\aligned_a_mant[0] ),
    .A2(\aligned_b_mant[0] ),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2535_ (.A1(_0430_),
    .A2(_0431_),
    .B(_1734_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2536_ (.I(_1726_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2537_ (.A1(_1722_),
    .A2(_0432_),
    .B(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _2538_ (.A1(_1738_),
    .A2(_1746_),
    .A3(_1754_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2539_ (.A1(_1742_),
    .A2(_0420_),
    .B(_1750_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2540_ (.I(_1758_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2541_ (.A1(_1754_),
    .A2(_0436_),
    .B(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2542_ (.A1(_0434_),
    .A2(_0435_),
    .B(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2543_ (.A1(_1746_),
    .A2(_1754_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2544_ (.A1(_1754_),
    .A2(_1748_),
    .B(_1756_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2545_ (.A1(_0412_),
    .A2(_0440_),
    .B(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2546_ (.A1(_1754_),
    .A2(_1745_),
    .B(_1753_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2547_ (.A1(_0415_),
    .A2(_0440_),
    .B(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2548_ (.I0(_0442_),
    .I1(_0444_),
    .S(_0416_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2549_ (.I0(_0439_),
    .I1(_0445_),
    .S(_0388_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2550_ (.A1(_0429_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2551_ (.A1(_0374_),
    .A2(_0447_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2552_ (.A1(_0429_),
    .A2(_0440_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2553_ (.A1(_0410_),
    .A2(_0411_),
    .B(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _2554_ (.A1(_0429_),
    .A2(_0441_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _2555_ (.A1(_0383_),
    .A2(_1764_),
    .A3(_0449_),
    .A4(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2556_ (.A1(_0413_),
    .A2(_0414_),
    .B(_0448_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _2557_ (.A1(_0429_),
    .A2(_0443_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _2558_ (.A1(is_a_larger_stage1),
    .A2(_1761_),
    .A3(_0452_),
    .A4(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2559_ (.I(_1766_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2560_ (.A1(_1762_),
    .A2(_0439_),
    .B(_0392_),
    .C(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2561_ (.A1(_0393_),
    .A2(_0451_),
    .A3(_0454_),
    .B(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2562_ (.A1(_1770_),
    .A2(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2563_ (.A1(_0374_),
    .A2(_0458_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2564_ (.A1(_1762_),
    .A2(_0455_),
    .B(_1770_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _2565_ (.A1(_1774_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2566_ (.A1(_1766_),
    .A2(_1774_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2567_ (.A1(_0434_),
    .A2(_0435_),
    .B(_0461_),
    .C(_0438_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2568_ (.A1(_0460_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2569_ (.A1(_1764_),
    .A2(_0449_),
    .A3(_0450_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2570_ (.A1(_1770_),
    .A2(_0464_),
    .B(_1772_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2571_ (.A1(_1761_),
    .A2(_0452_),
    .A3(_0453_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2572_ (.A1(_1770_),
    .A2(_0466_),
    .B(_1769_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2573_ (.I0(_0465_),
    .I1(_0467_),
    .S(_0384_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2574_ (.I0(_0463_),
    .I1(_0468_),
    .S(_0396_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2575_ (.A1(_1778_),
    .A2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2576_ (.A1(_0374_),
    .A2(_0470_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2577_ (.A1(_1778_),
    .A2(_0460_),
    .A3(_0462_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2578_ (.A1(_1782_),
    .A2(_0471_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2579_ (.A1(_1764_),
    .A2(_1772_),
    .A3(_1780_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2580_ (.A1(_1770_),
    .A2(_1772_),
    .A3(_1780_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2581_ (.A1(_1778_),
    .A2(_1780_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2582_ (.A1(_0474_),
    .A2(_0475_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2583_ (.A1(_0449_),
    .A2(_0450_),
    .A3(_0473_),
    .B(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2584_ (.A1(_1761_),
    .A2(_1769_),
    .A3(_1777_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2585_ (.A1(_1770_),
    .A2(_1769_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2586_ (.A1(_1778_),
    .A2(_0479_),
    .B(_1777_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2587_ (.I(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2588_ (.A1(_0452_),
    .A2(_0453_),
    .A3(_0478_),
    .B(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2589_ (.I0(_0477_),
    .I1(_0482_),
    .S(_0384_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2590_ (.I0(_0472_),
    .I1(_0483_),
    .S(_0396_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2591_ (.A1(_1786_),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2592_ (.A1(_0374_),
    .A2(_0485_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _2593_ (.I(_1786_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2594_ (.A1(_0486_),
    .A2(_0472_),
    .B(_1790_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2595_ (.I(_1785_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2596_ (.A1(_0486_),
    .A2(_0482_),
    .B(_0488_),
    .C(_0416_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2597_ (.I(_1788_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2598_ (.A1(is_a_larger_stage1),
    .A2(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2599_ (.A1(_0486_),
    .A2(_0477_),
    .B(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2600_ (.A1(_0387_),
    .A2(_0489_),
    .A3(_0492_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2601_ (.A1(_0393_),
    .A2(_0487_),
    .B(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2602_ (.A1(_1794_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2603_ (.A1(_0374_),
    .A2(_0495_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _2604_ (.I(_0373_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2605_ (.I(_1802_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2606_ (.A1(_1770_),
    .A2(_1778_),
    .A3(_1786_),
    .A4(_1794_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2607_ (.A1(_1794_),
    .A2(_1785_),
    .B(_1793_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2608_ (.I(_1794_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2609_ (.A1(_1778_),
    .A2(_1769_),
    .B(_1777_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2610_ (.A1(_0486_),
    .A2(_0500_),
    .A3(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2611_ (.A1(_0383_),
    .A2(_0499_),
    .A3(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2612_ (.A1(_1778_),
    .A2(_1772_),
    .B(_1780_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2613_ (.A1(_0486_),
    .A2(_0504_),
    .B(_0490_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2614_ (.A1(_1794_),
    .A2(_0505_),
    .B(_1796_),
    .C(_0383_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2615_ (.A1(_0451_),
    .A2(_0454_),
    .A3(_0498_),
    .B1(_0503_),
    .B2(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2616_ (.A1(_1794_),
    .A2(_0487_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2617_ (.A1(_1798_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2618_ (.I0(_0507_),
    .I1(_0509_),
    .S(_0392_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2619_ (.A1(_0497_),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2620_ (.A1(_0496_),
    .A2(_0511_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2621_ (.I(_1810_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2622_ (.A1(_1786_),
    .A2(_1794_),
    .A3(_1802_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2623_ (.I(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2624_ (.I(_1782_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2625_ (.I(_1790_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2626_ (.A1(_0515_),
    .A2(_1786_),
    .B(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2627_ (.A1(_0500_),
    .A2(_0517_),
    .B(_1798_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2628_ (.I(_1806_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2629_ (.A1(_1802_),
    .A2(_0518_),
    .B(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2630_ (.A1(_0471_),
    .A2(_0514_),
    .B(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2631_ (.A1(_1802_),
    .A2(_1796_),
    .B(_1804_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2632_ (.A1(_0491_),
    .A2(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2633_ (.A1(_0477_),
    .A2(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2634_ (.A1(_1794_),
    .A2(_1802_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2635_ (.A1(_1802_),
    .A2(_1793_),
    .B(_1801_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2636_ (.I0(_0522_),
    .I1(_0526_),
    .S(_0383_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2637_ (.A1(_0383_),
    .A2(_0488_),
    .A3(_0526_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2638_ (.A1(_0523_),
    .A2(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _2639_ (.A1(_0525_),
    .A2(_0527_),
    .B1(_0528_),
    .B2(_0482_),
    .C1(_0486_),
    .C2(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2640_ (.A1(_0524_),
    .A2(_0530_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2641_ (.I0(_0521_),
    .I1(_0531_),
    .S(_0396_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2642_ (.A1(_0512_),
    .A2(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2643_ (.A1(_0496_),
    .A2(_0533_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2644_ (.I(_1814_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2645_ (.A1(_1810_),
    .A2(_0521_),
    .B(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2646_ (.A1(_0486_),
    .A2(_0500_),
    .A3(_0497_),
    .A4(_0512_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2647_ (.A1(_1794_),
    .A2(_1788_),
    .B(_1796_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2648_ (.I(_1804_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2649_ (.A1(_0497_),
    .A2(_0537_),
    .B(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2650_ (.A1(_1810_),
    .A2(_0539_),
    .B(_1812_),
    .C(_0383_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2651_ (.A1(_0477_),
    .A2(_0536_),
    .B(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2652_ (.A1(is_a_larger_stage1),
    .A2(_1809_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2653_ (.A1(_0497_),
    .A2(_0499_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2654_ (.A1(_1801_),
    .A2(_0543_),
    .B(_1810_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2655_ (.A1(_0482_),
    .A2(_0536_),
    .B(_0542_),
    .C(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2656_ (.A1(_0541_),
    .A2(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2657_ (.I0(_0535_),
    .I1(_0546_),
    .S(_0396_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2658_ (.A1(_1818_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2659_ (.A1(_0496_),
    .A2(_0548_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2660_ (.I(_1826_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2661_ (.I(_1818_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2662_ (.A1(_0550_),
    .A2(_0535_),
    .B(_1822_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2663_ (.I(_1820_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2664_ (.A1(_0512_),
    .A2(_0550_),
    .A3(_0525_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2665_ (.A1(_0512_),
    .A2(_0522_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2666_ (.A1(_1812_),
    .A2(_0554_),
    .B(_1818_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2667_ (.A1(is_a_larger_stage1),
    .A2(_0552_),
    .A3(_0553_),
    .A4(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2668_ (.A1(_0512_),
    .A2(_0526_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2669_ (.A1(_1809_),
    .A2(_0557_),
    .B(_1818_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2670_ (.I(_1817_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2671_ (.A1(_0382_),
    .A2(_0559_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2672_ (.A1(_0488_),
    .A2(_0553_),
    .B(_0558_),
    .C(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2673_ (.A1(_0556_),
    .A2(_0561_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2674_ (.A1(_0482_),
    .A2(_0553_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2675_ (.A1(is_a_larger_stage1),
    .A2(_0490_),
    .A3(_0552_),
    .A4(_0555_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2676_ (.I(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2677_ (.A1(_0562_),
    .A2(_0564_),
    .B(_1786_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2678_ (.A1(_0477_),
    .A2(_0565_),
    .B(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2679_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2680_ (.A1(_0392_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2681_ (.A1(_0392_),
    .A2(_0551_),
    .B(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2682_ (.A1(_0549_),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2683_ (.A1(_0496_),
    .A2(_0571_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2684_ (.I(_1830_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2685_ (.A1(_0549_),
    .A2(_0551_),
    .B(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2686_ (.A1(_1802_),
    .A2(_1810_),
    .A3(_1818_),
    .A4(_0549_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2687_ (.A1(_1810_),
    .A2(_1801_),
    .B(_1809_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2688_ (.A1(_0550_),
    .A2(_0575_),
    .B(_0559_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2689_ (.A1(_0549_),
    .A2(_0576_),
    .B(_1825_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2690_ (.A1(_1810_),
    .A2(_1804_),
    .B(_1812_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2691_ (.A1(_0550_),
    .A2(_0578_),
    .B(_0552_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2692_ (.A1(_0549_),
    .A2(_0579_),
    .B(_1828_),
    .C(_0383_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2693_ (.A1(_0384_),
    .A2(_0577_),
    .B(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2694_ (.A1(_0507_),
    .A2(_0574_),
    .B(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2695_ (.I0(_0573_),
    .I1(_0582_),
    .S(_0396_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2696_ (.A1(_1834_),
    .A2(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2697_ (.A1(_0496_),
    .A2(_0584_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2698_ (.I(_1842_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _2699_ (.I(_1834_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2700_ (.A1(_0586_),
    .A2(_0573_),
    .B(_0388_),
    .C(_1838_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2701_ (.A1(_1810_),
    .A2(_1818_),
    .A3(_0549_),
    .A4(_1834_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2702_ (.I(_1826_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2703_ (.A1(_1818_),
    .A2(_1812_),
    .B(_1820_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2704_ (.I(_1828_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2705_ (.A1(_0589_),
    .A2(_0590_),
    .B(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2706_ (.A1(_1834_),
    .A2(_0592_),
    .B(_1836_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2707_ (.A1(_1818_),
    .A2(_1809_),
    .B(_1817_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2708_ (.I(_1825_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2709_ (.A1(_0589_),
    .A2(_0594_),
    .B(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2710_ (.A1(_1834_),
    .A2(_0596_),
    .B(_1833_),
    .C(is_a_larger_stage1),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _2711_ (.A1(_0379_),
    .A2(_0593_),
    .B(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2712_ (.A1(_0531_),
    .A2(_0588_),
    .B(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2713_ (.A1(_0393_),
    .A2(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2714_ (.A1(_0585_),
    .A2(_0587_),
    .A3(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2715_ (.A1(_0587_),
    .A2(_0600_),
    .B(_0585_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2716_ (.A1(_0373_),
    .A2(_0601_),
    .A3(_0602_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2717_ (.I(_1850_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2718_ (.A1(_1818_),
    .A2(_1826_),
    .A3(_1834_),
    .A4(_1842_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2719_ (.A1(_0512_),
    .A2(_0520_),
    .B(_1814_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2720_ (.A1(_0604_),
    .A2(_0605_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2721_ (.A1(_1738_),
    .A2(_1746_),
    .A3(_1754_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2722_ (.I(_1754_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2723_ (.I(_1750_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2724_ (.A1(_0408_),
    .A2(_1746_),
    .B(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2725_ (.A1(_0608_),
    .A2(_0610_),
    .B(_0461_),
    .C(_1758_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2726_ (.A1(_0395_),
    .A2(_0607_),
    .B(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2727_ (.A1(_1778_),
    .A2(_1810_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _2728_ (.A1(_0460_),
    .A2(_0513_),
    .A3(_0604_),
    .A4(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2729_ (.I(_1838_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2730_ (.I(_1822_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2731_ (.A1(_0616_),
    .A2(_1826_),
    .B(_0572_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2732_ (.A1(_0586_),
    .A2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2733_ (.A1(_0615_),
    .A2(_0618_),
    .B(_1842_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2734_ (.A1(_0612_),
    .A2(_0614_),
    .B(_0619_),
    .C(_1846_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2735_ (.A1(_0606_),
    .A2(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2736_ (.A1(_0549_),
    .A2(_1820_),
    .B(_1828_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2737_ (.I(_1836_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2738_ (.A1(_0586_),
    .A2(_0622_),
    .B(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2739_ (.A1(_0585_),
    .A2(_0624_),
    .B(_1844_),
    .C(_0384_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2740_ (.A1(_0549_),
    .A2(_1817_),
    .B(_1825_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2741_ (.I(_1833_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2742_ (.A1(_0586_),
    .A2(_0626_),
    .B(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2743_ (.A1(_0585_),
    .A2(_0628_),
    .B(_1841_),
    .C(_0379_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2744_ (.A1(_1818_),
    .A2(_0549_),
    .A3(_1834_),
    .A4(_0585_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _2745_ (.A1(_0625_),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0546_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2746_ (.I0(_0621_),
    .I1(_0631_),
    .S(_0396_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2747_ (.A1(_0603_),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2748_ (.A1(_0496_),
    .A2(_0633_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _2749_ (.I(_1858_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _2750_ (.A1(_0604_),
    .A2(_0605_),
    .B(_0620_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2751_ (.A1(_0603_),
    .A2(_0635_),
    .B(_1854_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2752_ (.I(_1852_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2753_ (.A1(_0586_),
    .A2(_0591_),
    .B(_0623_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2754_ (.A1(_0585_),
    .A2(_0638_),
    .B(_1844_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2755_ (.A1(_0603_),
    .A2(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2756_ (.A1(_0379_),
    .A2(_0637_),
    .A3(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2757_ (.I(_1849_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2758_ (.A1(_0586_),
    .A2(_0595_),
    .B(_0627_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2759_ (.A1(_0585_),
    .A2(_0643_),
    .B(_1841_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2760_ (.A1(_0603_),
    .A2(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2761_ (.A1(_0384_),
    .A2(_0642_),
    .A3(_0645_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2762_ (.A1(_1834_),
    .A2(_0585_),
    .A3(_1850_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2763_ (.A1(_0549_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2764_ (.A1(_0641_),
    .A2(_0646_),
    .B1(_0648_),
    .B2(_0568_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2765_ (.I0(_0636_),
    .I1(_0649_),
    .S(_0396_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2766_ (.A1(_0634_),
    .A2(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2767_ (.A1(_0496_),
    .A2(_0651_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2768_ (.I(_1866_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2769_ (.I(_1862_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2770_ (.I(_1858_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2771_ (.A1(_0654_),
    .A2(_0636_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2772_ (.A1(_0653_),
    .A2(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2773_ (.A1(_0585_),
    .A2(_1836_),
    .B(_1844_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2774_ (.A1(_0603_),
    .A2(_0657_),
    .B(_0637_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2775_ (.A1(_0654_),
    .A2(_0658_),
    .B(_1860_),
    .C(_0416_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2776_ (.A1(_0585_),
    .A2(_1833_),
    .B(_1841_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2777_ (.A1(_0603_),
    .A2(_0660_),
    .B(_0642_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2778_ (.A1(_0654_),
    .A2(_0661_),
    .B(_1857_),
    .C(_0379_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2779_ (.A1(_0654_),
    .A2(_0647_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2780_ (.A1(_0659_),
    .A2(_0662_),
    .B1(_0663_),
    .B2(_0582_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2781_ (.I0(_0656_),
    .I1(_0664_),
    .S(_0388_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2782_ (.A1(_0652_),
    .A2(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2783_ (.A1(_0496_),
    .A2(_0666_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2784_ (.I(_1870_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _2785_ (.A1(_1850_),
    .A2(_0654_),
    .A3(_1866_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2786_ (.A1(_1854_),
    .A2(_0634_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2787_ (.A1(_0653_),
    .A2(_0669_),
    .B(_1866_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2788_ (.A1(_0635_),
    .A2(_0668_),
    .B(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2789_ (.A1(_0667_),
    .A2(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2790_ (.A1(_1842_),
    .A2(_1850_),
    .A3(_0654_),
    .A4(_1866_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2791_ (.A1(_0588_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2792_ (.A1(_0477_),
    .A2(_0523_),
    .B(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2793_ (.A1(_1850_),
    .A2(_1841_),
    .B(_1849_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2794_ (.I(_1857_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2795_ (.A1(_0634_),
    .A2(_0676_),
    .B(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2796_ (.A1(_0652_),
    .A2(_0678_),
    .B(_1865_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2797_ (.A1(_1850_),
    .A2(_1844_),
    .B(_1852_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2798_ (.I(_1860_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2799_ (.A1(_0634_),
    .A2(_0680_),
    .B(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2800_ (.A1(_0652_),
    .A2(_0682_),
    .B(_1868_),
    .C(_0383_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2801_ (.A1(_0384_),
    .A2(_0679_),
    .B(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2802_ (.A1(_0598_),
    .A2(_0673_),
    .B1(_0675_),
    .B2(_0530_),
    .C(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2803_ (.I0(_0672_),
    .I1(_0685_),
    .S(_0396_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2804_ (.A1(_1874_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2805_ (.A1(_0496_),
    .A2(_0687_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _2806_ (.I(_1882_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2807_ (.A1(_0688_),
    .A2(_0373_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2808_ (.A1(_1882_),
    .A2(_0373_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2809_ (.A1(_1850_),
    .A2(_0654_),
    .A3(_0652_),
    .A4(_1874_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2810_ (.A1(_0631_),
    .A2(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2811_ (.I(_1868_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2812_ (.A1(_0654_),
    .A2(_1852_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2813_ (.A1(_1860_),
    .A2(_0694_),
    .B(_0652_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2814_ (.A1(_0693_),
    .A2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2815_ (.A1(_1874_),
    .A2(_0696_),
    .B(_1876_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2816_ (.I(_1865_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2817_ (.A1(_0654_),
    .A2(_1849_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2818_ (.A1(_1857_),
    .A2(_0699_),
    .B(_0652_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2819_ (.A1(_0698_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2820_ (.A1(_1874_),
    .A2(_0701_),
    .B(_1873_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2821_ (.I0(_0697_),
    .I1(_0702_),
    .S(_0384_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2822_ (.A1(_0388_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2823_ (.I(_1874_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2824_ (.A1(_0705_),
    .A2(_0672_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2825_ (.A1(_1878_),
    .A2(_0706_),
    .B(_0393_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2826_ (.A1(_0692_),
    .A2(_0704_),
    .B(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2827_ (.I0(_0689_),
    .I1(_0690_),
    .S(_0708_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2828_ (.I(_1890_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2829_ (.A1(_0709_),
    .A2(_0373_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2830_ (.A1(_0369_),
    .A2(_0372_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2831_ (.A1(_0709_),
    .A2(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2832_ (.A1(_1870_),
    .A2(_1878_),
    .A3(_1886_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2833_ (.A1(_0635_),
    .A2(_0668_),
    .B(_0670_),
    .C(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2834_ (.A1(_0705_),
    .A2(_1878_),
    .A3(_1886_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2835_ (.A1(_0688_),
    .A2(_1886_),
    .B(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2836_ (.A1(_0714_),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2837_ (.A1(_1874_),
    .A2(_1882_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _2838_ (.A1(_0654_),
    .A2(_0652_),
    .A3(_0649_),
    .A4(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2839_ (.A1(_0652_),
    .A2(_1860_),
    .B(_1868_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2840_ (.I(_1876_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2841_ (.A1(_0705_),
    .A2(_0720_),
    .B(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2842_ (.A1(_1882_),
    .A2(_0722_),
    .B(_1884_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2843_ (.A1(_0652_),
    .A2(_1857_),
    .B(_1865_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2844_ (.I(_1873_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2845_ (.A1(_0705_),
    .A2(_0724_),
    .B(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2846_ (.A1(_1882_),
    .A2(_0726_),
    .B(_1881_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2847_ (.I0(_0723_),
    .I1(_0727_),
    .S(_0416_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2848_ (.A1(_0388_),
    .A2(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2849_ (.A1(_0393_),
    .A2(_0717_),
    .B1(_0719_),
    .B2(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2850_ (.I0(_0710_),
    .I1(_0712_),
    .S(_0730_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _2851_ (.I(_1898_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2852_ (.A1(_0731_),
    .A2(_0373_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2853_ (.A1(_1898_),
    .A2(_0373_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2854_ (.A1(_0652_),
    .A2(_0709_),
    .A3(_0664_),
    .A4(_0718_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2855_ (.A1(_1874_),
    .A2(_1865_),
    .B(_1873_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2856_ (.I(_1881_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2857_ (.A1(_0688_),
    .A2(_0735_),
    .B(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2858_ (.A1(_0709_),
    .A2(_0737_),
    .B(_1889_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2859_ (.A1(_1874_),
    .A2(_1868_),
    .B(_1876_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2860_ (.I(_1884_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2861_ (.A1(_0688_),
    .A2(_0739_),
    .B(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2862_ (.A1(_0709_),
    .A2(_0741_),
    .B(_1892_),
    .C(_0416_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2863_ (.A1(_0416_),
    .A2(_0738_),
    .B(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2864_ (.I(_1894_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2865_ (.A1(_0709_),
    .A2(_0714_),
    .A3(_0716_),
    .B(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2866_ (.A1(_0393_),
    .A2(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2867_ (.A1(_0393_),
    .A2(_0734_),
    .A3(_0743_),
    .B(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2868_ (.I0(_0732_),
    .I1(_0733_),
    .S(_0747_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2869_ (.A1(_0731_),
    .A2(_0745_),
    .B(_1902_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2870_ (.I(_1900_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2871_ (.A1(_0688_),
    .A2(_0721_),
    .B(_0740_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2872_ (.A1(_0709_),
    .A2(_0750_),
    .B(_1892_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2873_ (.A1(_0731_),
    .A2(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2874_ (.A1(_0379_),
    .A2(_0749_),
    .A3(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2875_ (.I(_1897_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2876_ (.A1(_0688_),
    .A2(_0725_),
    .B(_0736_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2877_ (.A1(_0709_),
    .A2(_0755_),
    .B(_1889_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2878_ (.A1(_0731_),
    .A2(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2879_ (.A1(_0416_),
    .A2(_0754_),
    .A3(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2880_ (.A1(_0709_),
    .A2(_1898_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2881_ (.A1(_0718_),
    .A2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2882_ (.A1(_0753_),
    .A2(_0758_),
    .B1(_0760_),
    .B2(_0685_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2883_ (.I0(_0748_),
    .I1(_0761_),
    .S(_0388_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2884_ (.A1(_1906_),
    .A2(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2885_ (.A1(_0496_),
    .A2(_0763_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2886_ (.I(_1914_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2887_ (.A1(_1906_),
    .A2(_0387_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2888_ (.A1(_1882_),
    .A2(_0691_),
    .A3(_0759_),
    .A4(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2889_ (.I(_1910_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2890_ (.A1(_0767_),
    .A2(_0392_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2891_ (.A1(_1882_),
    .A2(_0759_),
    .A3(_0765_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2892_ (.A1(_0709_),
    .A2(_1884_),
    .B(_1892_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2893_ (.A1(_0731_),
    .A2(_0770_),
    .B(_0749_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2894_ (.A1(_1906_),
    .A2(_0771_),
    .B(_1908_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2895_ (.A1(_1890_),
    .A2(_1881_),
    .B(_1889_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2896_ (.A1(_0731_),
    .A2(_0773_),
    .B(_0754_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2897_ (.A1(_1906_),
    .A2(_0774_),
    .B(_1905_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2898_ (.I0(_0772_),
    .I1(_0775_),
    .S(_0383_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2899_ (.A1(_1906_),
    .A2(_0767_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2900_ (.I0(_0776_),
    .I1(_0777_),
    .S(_0392_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2901_ (.A1(_0703_),
    .A2(_0769_),
    .B(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2902_ (.A1(_0631_),
    .A2(_0766_),
    .B1(_0768_),
    .B2(_0748_),
    .C(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2903_ (.A1(_0764_),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2904_ (.A1(_0374_),
    .A2(_0781_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2905_ (.A1(_0719_),
    .A2(_0728_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2906_ (.A1(_1906_),
    .A2(_1914_),
    .A3(_0388_),
    .A4(_0759_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2907_ (.I(_1908_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2908_ (.A1(_1898_),
    .A2(_1892_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2909_ (.A1(_1900_),
    .A2(_0785_),
    .B(_1906_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2910_ (.A1(_0784_),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2911_ (.A1(_1914_),
    .A2(_0787_),
    .B(_1916_),
    .C(_0416_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2912_ (.I(_1905_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2913_ (.A1(_1898_),
    .A2(_1889_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2914_ (.A1(_1897_),
    .A2(_0790_),
    .B(_1906_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2915_ (.A1(_0789_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2916_ (.A1(_1914_),
    .A2(_0792_),
    .B(_1913_),
    .C(_0379_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2917_ (.A1(_0393_),
    .A2(_0788_),
    .A3(_0793_),
    .B(_0373_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2918_ (.A1(_1906_),
    .A2(_0748_),
    .B(_0767_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2919_ (.A1(_0764_),
    .A2(_0795_),
    .B(_0388_),
    .C(_1918_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2920_ (.A1(_0782_),
    .A2(_0783_),
    .B(_0794_),
    .C(_0796_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2921_ (.A1(_1220_),
    .A2(_1221_),
    .A3(_1222_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2922_ (.A1(net58),
    .A2(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2923_ (.I0(b_sign_stage1),
    .I1(a_sign_stage1),
    .S(_0379_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2924_ (.I0(_0798_),
    .I1(_0799_),
    .S(_0372_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2925_ (.A1(_1209_),
    .A2(_1210_),
    .A3(_1211_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2926_ (.I(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2927_ (.A1(_1577_),
    .A2(_0797_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2928_ (.I0(_0803_),
    .I1(net26),
    .S(_0372_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2929_ (.A1(_0802_),
    .A2(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2930_ (.A1(_0367_),
    .A2(_0368_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2931_ (.I0(_0800_),
    .I1(_0805_),
    .S(_0806_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2932_ (.I(\result_exp_stage2[4] ),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2933_ (.I(\result_exp_stage2[3] ),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2934_ (.I(\result_exp_stage2[2] ),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2935_ (.A1(\result_exp_stage2[5] ),
    .A2(_0807_),
    .A3(_0808_),
    .A4(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2936_ (.A1(\result_exp_stage2[6] ),
    .A2(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _2937_ (.A1(\result_exp_stage2[7] ),
    .A2(_1716_),
    .A3(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2938_ (.A1(_0327_),
    .A2(_0812_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2939_ (.I(net25),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2940_ (.I(net23),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2941_ (.I(net22),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2942_ (.I(net21),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2943_ (.I(net20),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2944_ (.I(net19),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2945_ (.I(net18),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2946_ (.I(_1689_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2947_ (.I(net17),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2948_ (.I(\aligned_a_mant[2] ),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2949_ (.I(\aligned_a_mant[1] ),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2950_ (.I(\aligned_a_mant[3] ),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2951_ (.I(\aligned_a_mant[4] ),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2952_ (.I(\aligned_a_mant[5] ),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2953_ (.I(\aligned_a_mant[6] ),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2954_ (.I(\aligned_a_mant[7] ),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2955_ (.I(\aligned_a_mant[8] ),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2956_ (.I(\aligned_a_mant[9] ),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2957_ (.I(\aligned_a_mant[10] ),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2958_ (.I(\aligned_a_mant[11] ),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2959_ (.I(\aligned_a_mant[12] ),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2960_ (.I(\aligned_a_mant[13] ),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2961_ (.I(\aligned_a_mant[14] ),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2962_ (.I(\aligned_a_mant[15] ),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2963_ (.I(\aligned_a_mant[16] ),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2964_ (.I(\aligned_a_mant[17] ),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2965_ (.I(\aligned_a_mant[18] ),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2966_ (.I(\aligned_a_mant[19] ),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2967_ (.I(\aligned_a_mant[20] ),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2968_ (.I(\aligned_a_mant[21] ),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2969_ (.I(\aligned_a_mant[22] ),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2970_ (.I(\aligned_a_mant[23] ),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2971_ (.I(\aligned_a_mant[24] ),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2972_ (.I(\aligned_a_mant[25] ),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2973_ (.I(net57),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2974_ (.I(net55),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2975_ (.I(net54),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2976_ (.I(net53),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2977_ (.I(net52),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2978_ (.I(net51),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2979_ (.I(net50),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2980_ (.I(net49),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2981_ (.I(_0345_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2982_ (.I(_1702_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2983_ (.I(_0813_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2984_ (.I(_0352_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2985_ (.I(\aligned_b_mant[2] ),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2986_ (.I(\aligned_b_mant[1] ),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2987_ (.I(\aligned_b_mant[3] ),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2988_ (.I(\aligned_b_mant[4] ),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2989_ (.I(\aligned_b_mant[5] ),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2990_ (.I(\aligned_b_mant[6] ),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2991_ (.I(\aligned_b_mant[7] ),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2992_ (.I(\aligned_b_mant[8] ),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2993_ (.I(\aligned_b_mant[9] ),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2994_ (.I(\aligned_b_mant[10] ),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2995_ (.I(\aligned_b_mant[11] ),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2996_ (.I(\aligned_b_mant[12] ),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2997_ (.I(\aligned_b_mant[13] ),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2998_ (.I(\aligned_b_mant[14] ),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2999_ (.I(\aligned_b_mant[15] ),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3000_ (.I(\aligned_b_mant[16] ),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3001_ (.I(\aligned_b_mant[17] ),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3002_ (.I(\aligned_b_mant[18] ),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3003_ (.I(\aligned_b_mant[19] ),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3004_ (.I(\aligned_b_mant[20] ),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3005_ (.I(\aligned_b_mant[21] ),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3006_ (.I(\aligned_b_mant[22] ),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3007_ (.I(\aligned_b_mant[23] ),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3008_ (.I(\aligned_b_mant[24] ),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3009_ (.I(\aligned_b_mant[25] ),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _3010_ (.A1(\result_exp_stage2[7] ),
    .A2(_0359_),
    .A3(_0361_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3011_ (.A1(_0342_),
    .A2(_0814_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _3012_ (.A1(_0354_),
    .A2(_0815_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3013_ (.I0(_1707_),
    .I1(_1710_),
    .S(_0342_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3014_ (.A1(_0343_),
    .A2(_0366_),
    .A3(_0812_),
    .B1(_0816_),
    .B2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3015_ (.I(net66),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3016_ (.I0(\final_exp[0] ),
    .I1(_0818_),
    .S(_0819_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3017_ (.I(_1715_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3018_ (.I(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3019_ (.I(_0816_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3020_ (.I0(_1576_),
    .I1(\result_exp_stage2[1] ),
    .S(_0328_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3021_ (.A1(_0327_),
    .A2(_0821_),
    .B1(_0822_),
    .B2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3022_ (.I(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3023_ (.I0(\final_exp[1] ),
    .I1(_0825_),
    .S(_0819_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3024_ (.A1(_1697_),
    .A2(_1575_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3025_ (.I0(_1694_),
    .I1(_0826_),
    .S(_0342_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3026_ (.A1(_0809_),
    .A2(_1718_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3027_ (.I(\add_result[26] ),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3028_ (.A1(_0812_),
    .A2(_0828_),
    .B(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3029_ (.A1(_0816_),
    .A2(_0827_),
    .B(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3030_ (.I0(\final_exp[2] ),
    .I1(_0831_),
    .S(_0819_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3031_ (.A1(_1573_),
    .A2(_1704_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3032_ (.A1(_1705_),
    .A2(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3033_ (.A1(_1697_),
    .A2(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3034_ (.A1(_0328_),
    .A2(_1699_),
    .A3(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3035_ (.A1(_0808_),
    .A2(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3036_ (.A1(\result_exp_stage2[1] ),
    .A2(_0366_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3037_ (.A1(_0809_),
    .A2(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3038_ (.A1(_0808_),
    .A2(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3039_ (.A1(_0812_),
    .A2(_0839_),
    .B(_0829_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3040_ (.A1(_0816_),
    .A2(_0836_),
    .B(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3041_ (.I0(\final_exp[3] ),
    .I1(_0841_),
    .S(_0819_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3042_ (.A1(_0328_),
    .A2(_0808_),
    .A3(_1699_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3043_ (.A1(_1697_),
    .A2(_1575_),
    .B(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3044_ (.A1(_0807_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3045_ (.A1(_0808_),
    .A2(_0809_),
    .A3(_1718_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3046_ (.A1(_0807_),
    .A2(_0845_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3047_ (.A1(_0812_),
    .A2(_0846_),
    .B(_0829_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3048_ (.A1(_0816_),
    .A2(_0844_),
    .B(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3049_ (.I0(\final_exp[4] ),
    .I1(_0848_),
    .S(_0819_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3050_ (.A1(_0807_),
    .A2(_0808_),
    .A3(_0835_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3051_ (.A1(\result_exp_stage2[5] ),
    .A2(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3052_ (.A1(_0807_),
    .A2(_0808_),
    .A3(_0809_),
    .A4(_0837_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3053_ (.A1(\result_exp_stage2[5] ),
    .A2(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3054_ (.A1(_0812_),
    .A2(_0852_),
    .B(\add_result[26] ),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3055_ (.A1(_0816_),
    .A2(_0850_),
    .B(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3056_ (.I0(\final_exp[5] ),
    .I1(_0854_),
    .S(_0819_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3057_ (.A1(\result_exp_stage2[5] ),
    .A2(_0807_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3058_ (.A1(_0855_),
    .A2(_0843_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3059_ (.A1(\result_exp_stage2[6] ),
    .A2(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3060_ (.A1(_1718_),
    .A2(_0810_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3061_ (.A1(\result_exp_stage2[6] ),
    .A2(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3062_ (.A1(_0812_),
    .A2(_0859_),
    .B(\add_result[26] ),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3063_ (.A1(_0816_),
    .A2(_0857_),
    .B(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3064_ (.I0(\final_exp[6] ),
    .I1(_0861_),
    .S(_0819_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3065_ (.I(_0343_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3066_ (.I(\result_exp_stage2[7] ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3067_ (.A1(_0863_),
    .A2(_1716_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3068_ (.A1(_0811_),
    .A2(_0837_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3069_ (.I0(_0863_),
    .I1(_0864_),
    .S(_0865_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3070_ (.A1(_0361_),
    .A2(_0835_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3071_ (.A1(\result_exp_stage2[7] ),
    .A2(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _3072_ (.A1(_0862_),
    .A2(_0866_),
    .B1(_0868_),
    .B2(_0816_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3073_ (.I0(\final_exp[7] ),
    .I1(_0869_),
    .S(_0819_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3074_ (.A1(_0863_),
    .A2(_1714_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _3075_ (.A1(_0809_),
    .A2(_0361_),
    .A3(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3076_ (.A1(_0814_),
    .A2(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3077_ (.A1(_0328_),
    .A2(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3078_ (.I(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3079_ (.I(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3080_ (.A1(\result_exp_stage2[2] ),
    .A2(_1714_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3081_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3082_ (.A1(_0807_),
    .A2(_1714_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3083_ (.A1(\result_exp_stage2[1] ),
    .A2(_0364_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3084_ (.A1(\result_exp_stage2[4] ),
    .A2(_1714_),
    .A3(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3085_ (.I0(_0878_),
    .I1(_0880_),
    .S(\result_exp_stage2[5] ),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3086_ (.A1(_0808_),
    .A2(_0809_),
    .A3(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3087_ (.A1(\result_exp_stage2[1] ),
    .A2(_0364_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3088_ (.A1(_1714_),
    .A2(_0883_),
    .B(_1694_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3089_ (.A1(_0808_),
    .A2(_0884_),
    .B(_0855_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _3090_ (.A1(_0882_),
    .A2(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3091_ (.A1(\result_exp_stage2[3] ),
    .A2(\result_exp_stage2[2] ),
    .A3(_0879_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3092_ (.A1(_0809_),
    .A2(_0879_),
    .B(\result_exp_stage2[3] ),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3093_ (.A1(_0887_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3094_ (.A1(_0886_),
    .A2(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3095_ (.A1(_0877_),
    .A2(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3096_ (.A1(_0365_),
    .A2(\add_result[2] ),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3097_ (.A1(_0360_),
    .A2(_0884_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3098_ (.A1(_0863_),
    .A2(_1714_),
    .A3(_0879_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3099_ (.I0(_0894_),
    .I1(_0870_),
    .S(\result_exp_stage2[6] ),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _3100_ (.A1(\result_exp_stage2[7] ),
    .A2(\result_exp_stage2[6] ),
    .A3(_0893_),
    .B1(_0895_),
    .B2(_0809_),
    .B3(_0360_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3101_ (.A1(_0820_),
    .A2(_0892_),
    .A3(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3102_ (.A1(_0815_),
    .A2(_0891_),
    .A3(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3103_ (.A1(\add_result[2] ),
    .A2(_0875_),
    .B(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3104_ (.A1(\add_result[3] ),
    .A2(_0327_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3105_ (.A1(_0354_),
    .A2(_0899_),
    .B(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3106_ (.I0(\final_mant[0] ),
    .I1(_0901_),
    .S(_0819_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3107_ (.I(_0896_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3108_ (.I(_0902_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3109_ (.I0(\add_result[5] ),
    .I1(\add_result[6] ),
    .S(_0364_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3110_ (.I0(\add_result[7] ),
    .I1(\add_result[8] ),
    .S(_0364_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3111_ (.I0(_0904_),
    .I1(_0905_),
    .S(_1715_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3112_ (.I0(\add_result[9] ),
    .I1(\add_result[10] ),
    .S(_0364_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3113_ (.I0(\add_result[11] ),
    .I1(\add_result[12] ),
    .S(_0364_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3114_ (.I0(_0907_),
    .I1(_0908_),
    .S(_1715_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3115_ (.I0(_0906_),
    .I1(_0909_),
    .S(_0877_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3116_ (.A1(_0890_),
    .A2(_0903_),
    .A3(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3117_ (.I0(\add_result[6] ),
    .I1(\add_result[5] ),
    .S(_1708_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3118_ (.I0(\add_result[8] ),
    .I1(\add_result[7] ),
    .S(_1708_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3119_ (.I(_0813_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3120_ (.I0(_0912_),
    .I1(_0913_),
    .S(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3121_ (.I0(\add_result[10] ),
    .I1(\add_result[9] ),
    .S(_1708_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3122_ (.I0(\add_result[12] ),
    .I1(\add_result[11] ),
    .S(_1708_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3123_ (.I0(_0916_),
    .I1(_0917_),
    .S(_0914_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3124_ (.I0(_0915_),
    .I1(_0918_),
    .S(_0345_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3125_ (.I(_0362_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3126_ (.I0(_0911_),
    .I1(_0919_),
    .S(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3127_ (.I(_0342_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3128_ (.A1(\add_result[12] ),
    .A2(_0874_),
    .B1(_0921_),
    .B2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3129_ (.A1(\add_result[13] ),
    .A2(_0327_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3130_ (.A1(_0327_),
    .A2(_0923_),
    .B(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3131_ (.I0(\final_mant[10] ),
    .I1(_0925_),
    .S(_0819_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _3132_ (.I(net66),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3133_ (.I(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3134_ (.I(\add_result[14] ),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _3135_ (.I(_0890_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3136_ (.I0(\add_result[6] ),
    .I1(\add_result[7] ),
    .S(_0365_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3137_ (.I0(\add_result[8] ),
    .I1(\add_result[9] ),
    .S(_0365_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3138_ (.I0(_0930_),
    .I1(_0931_),
    .S(_0820_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3139_ (.I0(\add_result[10] ),
    .I1(\add_result[11] ),
    .S(_0366_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3140_ (.I0(\add_result[12] ),
    .I1(\add_result[13] ),
    .S(_0366_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3141_ (.I0(_0933_),
    .I1(_0934_),
    .S(_0821_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3142_ (.I0(_0932_),
    .I1(_0935_),
    .S(_0877_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3143_ (.A1(_0929_),
    .A2(_0903_),
    .A3(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3144_ (.I0(\add_result[6] ),
    .I1(\add_result[7] ),
    .S(_1711_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3145_ (.I0(\add_result[8] ),
    .I1(\add_result[9] ),
    .S(_1711_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3146_ (.I0(_0938_),
    .I1(_0939_),
    .S(_0914_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3147_ (.I0(\add_result[10] ),
    .I1(\add_result[11] ),
    .S(_1711_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3148_ (.I0(\add_result[12] ),
    .I1(\add_result[13] ),
    .S(_1711_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3149_ (.I0(_0941_),
    .I1(_0942_),
    .S(_1574_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3150_ (.I0(_0940_),
    .I1(_0943_),
    .S(_1698_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3151_ (.I0(_0937_),
    .I1(_0944_),
    .S(_0363_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3152_ (.I(_0342_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3153_ (.A1(\add_result[13] ),
    .A2(_0875_),
    .B1(_0945_),
    .B2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3154_ (.I0(_0928_),
    .I1(_0947_),
    .S(_0862_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3155_ (.A1(_0927_),
    .A2(\final_mant[11] ),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3156_ (.A1(_0927_),
    .A2(_0948_),
    .B(_0949_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3157_ (.I0(_0905_),
    .I1(_0907_),
    .S(_1715_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3158_ (.I0(\add_result[13] ),
    .I1(\add_result[14] ),
    .S(_0364_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3159_ (.I0(_0908_),
    .I1(_0951_),
    .S(_1715_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3160_ (.I0(_0950_),
    .I1(_0952_),
    .S(_0876_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3161_ (.A1(_0890_),
    .A2(_0903_),
    .A3(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3162_ (.I0(_0913_),
    .I1(_0916_),
    .S(_0914_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3163_ (.I0(\add_result[14] ),
    .I1(\add_result[13] ),
    .S(_0353_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3164_ (.I0(_0917_),
    .I1(_0956_),
    .S(_0914_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3165_ (.I0(_0955_),
    .I1(_0957_),
    .S(_0345_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3166_ (.I0(_0954_),
    .I1(_0958_),
    .S(_0920_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3167_ (.A1(\add_result[14] ),
    .A2(_0874_),
    .B1(_0959_),
    .B2(_0922_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3168_ (.A1(\add_result[15] ),
    .A2(_0327_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3169_ (.A1(_0327_),
    .A2(_0960_),
    .B(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3170_ (.I(net66),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3171_ (.I0(\final_mant[12] ),
    .I1(_0962_),
    .S(_0963_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3172_ (.I(\add_result[16] ),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3173_ (.I0(_0931_),
    .I1(_0933_),
    .S(_0820_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3174_ (.I0(\add_result[14] ),
    .I1(\add_result[15] ),
    .S(_0365_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3175_ (.I0(_0934_),
    .I1(_0966_),
    .S(_0820_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3176_ (.I(_0876_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3177_ (.I0(_0965_),
    .I1(_0967_),
    .S(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3178_ (.A1(_0929_),
    .A2(_0903_),
    .A3(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3179_ (.I0(_0939_),
    .I1(_0941_),
    .S(_1574_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3180_ (.I0(\add_result[14] ),
    .I1(\add_result[15] ),
    .S(_1711_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3181_ (.I0(_0942_),
    .I1(_0972_),
    .S(_1574_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3182_ (.I0(_0971_),
    .I1(_0973_),
    .S(_1698_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3183_ (.I0(_0970_),
    .I1(_0974_),
    .S(_0363_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3184_ (.A1(\add_result[15] ),
    .A2(_0875_),
    .B1(_0975_),
    .B2(_0946_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3185_ (.I0(_0964_),
    .I1(_0976_),
    .S(_0862_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3186_ (.A1(_0926_),
    .A2(\final_mant[13] ),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3187_ (.A1(_0927_),
    .A2(_0977_),
    .B(_0978_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3188_ (.I(\add_result[17] ),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3189_ (.I0(\add_result[15] ),
    .I1(\add_result[16] ),
    .S(_0364_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3190_ (.I0(_0951_),
    .I1(_0980_),
    .S(_1715_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3191_ (.I0(_0909_),
    .I1(_0981_),
    .S(_0876_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3192_ (.A1(_0929_),
    .A2(_0903_),
    .A3(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3193_ (.I0(\add_result[16] ),
    .I1(\add_result[15] ),
    .S(_1708_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3194_ (.I0(_0956_),
    .I1(_0984_),
    .S(_1574_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3195_ (.I0(_0918_),
    .I1(_0985_),
    .S(_1698_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3196_ (.I0(_0983_),
    .I1(_0986_),
    .S(_0363_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3197_ (.A1(\add_result[16] ),
    .A2(_0875_),
    .B1(_0987_),
    .B2(_0946_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3198_ (.I0(_0979_),
    .I1(_0988_),
    .S(_0862_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3199_ (.A1(_0926_),
    .A2(\final_mant[14] ),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3200_ (.A1(_0927_),
    .A2(_0989_),
    .B(_0990_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3201_ (.I0(\add_result[16] ),
    .I1(\add_result[17] ),
    .S(_0366_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3202_ (.I0(_0966_),
    .I1(_0991_),
    .S(_0821_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3203_ (.I0(_0935_),
    .I1(_0992_),
    .S(_0877_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3204_ (.A1(_0929_),
    .A2(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3205_ (.I0(\add_result[16] ),
    .I1(\add_result[17] ),
    .S(_1711_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3206_ (.I0(_0972_),
    .I1(_0995_),
    .S(_0914_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3207_ (.I0(_0943_),
    .I1(_0996_),
    .S(_0345_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3208_ (.I0(_0994_),
    .I1(_0997_),
    .S(_0920_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3209_ (.A1(\add_result[17] ),
    .A2(_0874_),
    .B1(_0998_),
    .B2(_0922_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3210_ (.A1(\add_result[18] ),
    .A2(_0829_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3211_ (.A1(_0327_),
    .A2(_0999_),
    .B(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3212_ (.I0(\final_mant[15] ),
    .I1(_1001_),
    .S(_0963_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3213_ (.I(\add_result[19] ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3214_ (.A1(_0878_),
    .A2(_0883_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3215_ (.A1(_0807_),
    .A2(_0879_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3216_ (.I0(_1003_),
    .I1(_1004_),
    .S(\result_exp_stage2[3] ),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3217_ (.A1(_0807_),
    .A2(_0808_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3218_ (.A1(_1006_),
    .A2(_0884_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _3219_ (.A1(_0809_),
    .A2(_1005_),
    .B(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3220_ (.I(_0902_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3221_ (.I0(\add_result[17] ),
    .I1(\add_result[18] ),
    .S(_0365_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3222_ (.I0(_0980_),
    .I1(_1010_),
    .S(_0821_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3223_ (.I0(_0952_),
    .I1(_1011_),
    .S(_0877_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3224_ (.A1(_1009_),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3225_ (.A1(_1714_),
    .A2(_0887_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3226_ (.A1(_0888_),
    .A2(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _3227_ (.A1(_0878_),
    .A2(_0887_),
    .B1(_1015_),
    .B2(_0807_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3228_ (.I0(\add_result[3] ),
    .I1(\add_result[4] ),
    .S(_0364_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3229_ (.I0(_1017_),
    .I1(_0904_),
    .S(_1715_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3230_ (.I0(_1018_),
    .I1(_0950_),
    .S(_0968_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3231_ (.A1(_1009_),
    .A2(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3232_ (.A1(\result_exp_stage2[5] ),
    .A2(_0889_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3233_ (.A1(_0968_),
    .A2(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3234_ (.A1(_0897_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _3235_ (.A1(_1008_),
    .A2(_1013_),
    .B1(_1016_),
    .B2(_1020_),
    .C1(_1023_),
    .C2(_0886_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3236_ (.I0(\add_result[18] ),
    .I1(\add_result[17] ),
    .S(_1708_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3237_ (.I0(_0984_),
    .I1(_1025_),
    .S(_0914_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3238_ (.I0(_0957_),
    .I1(_1026_),
    .S(_1698_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3239_ (.I0(_1024_),
    .I1(_1027_),
    .S(_0363_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3240_ (.A1(\add_result[18] ),
    .A2(_0875_),
    .B1(_1028_),
    .B2(_0946_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3241_ (.I0(_1002_),
    .I1(_1029_),
    .S(_0862_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3242_ (.A1(_0926_),
    .A2(\final_mant[16] ),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3243_ (.A1(_0927_),
    .A2(_1030_),
    .B(_1031_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3244_ (.I(_0331_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3245_ (.I0(\add_result[18] ),
    .I1(\add_result[19] ),
    .S(_0366_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3246_ (.I0(_0991_),
    .I1(_1033_),
    .S(_0821_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3247_ (.I0(_0967_),
    .I1(_1034_),
    .S(_0877_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3248_ (.A1(_1009_),
    .A2(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3249_ (.I0(\add_result[4] ),
    .I1(\add_result[5] ),
    .S(_0365_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3250_ (.I0(_1037_),
    .I1(_0930_),
    .S(_0820_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3251_ (.I0(_1038_),
    .I1(_0965_),
    .S(_0968_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3252_ (.A1(_1009_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3253_ (.I0(\add_result[2] ),
    .I1(\add_result[3] ),
    .S(_0365_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3254_ (.A1(_0821_),
    .A2(_1009_),
    .A3(_1022_),
    .A4(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _3255_ (.A1(_1008_),
    .A2(_1036_),
    .B1(_1040_),
    .B2(_1016_),
    .C1(_1042_),
    .C2(_0886_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3256_ (.I0(\add_result[18] ),
    .I1(\add_result[19] ),
    .S(_1711_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3257_ (.I0(_0995_),
    .I1(_1044_),
    .S(_1574_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3258_ (.I0(_0973_),
    .I1(_1045_),
    .S(_1698_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3259_ (.I0(_1043_),
    .I1(_1046_),
    .S(_0363_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3260_ (.A1(\add_result[19] ),
    .A2(_0875_),
    .B1(_1047_),
    .B2(_0946_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3261_ (.I0(_1032_),
    .I1(_1048_),
    .S(_0862_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3262_ (.A1(_0926_),
    .A2(\final_mant[17] ),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3263_ (.A1(_0927_),
    .A2(_1049_),
    .B(_1050_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3264_ (.A1(_0903_),
    .A2(_0910_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3265_ (.I0(\add_result[19] ),
    .I1(_0331_),
    .S(_0365_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3266_ (.I0(_1010_),
    .I1(_1052_),
    .S(_0820_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3267_ (.I0(_0981_),
    .I1(_1053_),
    .S(_0968_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3268_ (.A1(_1009_),
    .A2(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3269_ (.I0(_0892_),
    .I1(_1017_),
    .S(_1715_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3270_ (.A1(_0902_),
    .A2(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3271_ (.A1(_1022_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _3272_ (.A1(_1051_),
    .A2(_1016_),
    .B1(_1055_),
    .B2(_1008_),
    .C1(_1058_),
    .C2(_0886_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3273_ (.I0(\add_result[18] ),
    .I1(\add_result[17] ),
    .I2(_0331_),
    .I3(\add_result[19] ),
    .S0(_1708_),
    .S1(_0914_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3274_ (.I0(_0985_),
    .I1(_1060_),
    .S(_1698_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3275_ (.I0(_1059_),
    .I1(_1061_),
    .S(_0363_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3276_ (.A1(_0331_),
    .A2(_0875_),
    .B1(_1062_),
    .B2(_0946_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3277_ (.I0(_0349_),
    .I1(_1063_),
    .S(_0862_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3278_ (.A1(_0926_),
    .A2(\final_mant[18] ),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3279_ (.A1(_0927_),
    .A2(_1064_),
    .B(_1065_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3280_ (.A1(_0903_),
    .A2(_0936_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3281_ (.I0(_0331_),
    .I1(_0332_),
    .S(_0366_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3282_ (.I0(_0966_),
    .I1(_0991_),
    .I2(_1033_),
    .I3(_1067_),
    .S0(_0821_),
    .S1(_0877_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3283_ (.A1(_1009_),
    .A2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3284_ (.I0(_1041_),
    .I1(_1037_),
    .S(_0820_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3285_ (.A1(_0902_),
    .A2(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3286_ (.A1(_1022_),
    .A2(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _3287_ (.A1(_1066_),
    .A2(_1016_),
    .B1(_1069_),
    .B2(_1008_),
    .C1(_1072_),
    .C2(_0886_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3288_ (.I0(_0331_),
    .I1(_0332_),
    .S(_1711_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3289_ (.I0(_1044_),
    .I1(_1074_),
    .S(_1574_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3290_ (.I0(_0996_),
    .I1(_1075_),
    .S(_0345_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3291_ (.I0(_1073_),
    .I1(_1076_),
    .S(_0363_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3292_ (.A1(_0332_),
    .A2(_0875_),
    .B1(_1077_),
    .B2(_0946_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3293_ (.I0(_0333_),
    .I1(_1078_),
    .S(_0862_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3294_ (.A1(_0926_),
    .A2(\final_mant[19] ),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3295_ (.A1(_0927_),
    .A2(_1079_),
    .B(_1080_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3296_ (.A1(\add_result[24] ),
    .A2(\add_result[2] ),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3297_ (.I0(\add_result[3] ),
    .I1(_1081_),
    .S(_0347_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3298_ (.A1(_0821_),
    .A2(_0891_),
    .A3(_0903_),
    .A4(_1041_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3299_ (.I0(_1082_),
    .I1(_1083_),
    .S(_0814_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3300_ (.A1(\add_result[3] ),
    .A2(_0874_),
    .B1(_1084_),
    .B2(_0922_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3301_ (.A1(\add_result[4] ),
    .A2(_0829_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3302_ (.A1(_0354_),
    .A2(_1085_),
    .B(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3303_ (.I0(\final_mant[1] ),
    .I1(_1087_),
    .S(_0963_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3304_ (.A1(_0328_),
    .A2(_0872_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3305_ (.I(_0886_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3306_ (.A1(_0902_),
    .A2(_1018_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3307_ (.I0(_0897_),
    .I1(_1090_),
    .S(_0968_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3308_ (.A1(_1021_),
    .A2(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3309_ (.A1(_0902_),
    .A2(_0953_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3310_ (.I0(_0332_),
    .I1(\add_result[22] ),
    .S(_0365_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3311_ (.I0(_0980_),
    .I1(_1010_),
    .I2(_1052_),
    .I3(_1094_),
    .S0(_0820_),
    .S1(_0968_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3312_ (.A1(_0902_),
    .A2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3313_ (.A1(_1093_),
    .A2(_1016_),
    .B1(_1096_),
    .B2(_1008_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3314_ (.I(_0871_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _3315_ (.A1(_1089_),
    .A2(_1092_),
    .B(_1097_),
    .C(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3316_ (.I0(_0331_),
    .I1(\add_result[19] ),
    .I2(\add_result[22] ),
    .I3(_0332_),
    .S0(_1708_),
    .S1(_1574_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3317_ (.A1(_1695_),
    .A2(_1026_),
    .B(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3318_ (.I0(_1099_),
    .I1(_1101_),
    .S(_0920_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _3319_ (.A1(_0333_),
    .A2(_1088_),
    .B1(_1102_),
    .B2(_0328_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3320_ (.I0(\add_result[23] ),
    .I1(_1103_),
    .S(_0343_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3321_ (.I0(\final_mant[20] ),
    .I1(_1104_),
    .S(_0963_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3322_ (.A1(_1009_),
    .A2(_0969_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3323_ (.I0(\add_result[22] ),
    .I1(\add_result[23] ),
    .S(_0366_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3324_ (.I0(_0991_),
    .I1(_1033_),
    .I2(_1067_),
    .I3(_1106_),
    .S0(_0821_),
    .S1(_0877_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3325_ (.A1(_1009_),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3326_ (.A1(_1105_),
    .A2(_1016_),
    .B1(_1108_),
    .B2(_1008_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3327_ (.A1(_1098_),
    .A2(_1109_),
    .B(_0920_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3328_ (.A1(_0331_),
    .A2(_0334_),
    .B(\add_result[24] ),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3329_ (.A1(_0332_),
    .A2(_0346_),
    .B(_0344_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3330_ (.A1(_0333_),
    .A2(_0344_),
    .A3(_1111_),
    .B1(_1112_),
    .B2(_0334_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3331_ (.A1(_1695_),
    .A2(_1045_),
    .B(_1113_),
    .C(_0814_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3332_ (.A1(_0328_),
    .A2(_1110_),
    .A3(_1114_),
    .B1(_1088_),
    .B2(_0334_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3333_ (.I0(\add_result[24] ),
    .I1(_1115_),
    .S(_0343_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3334_ (.I0(\final_mant[21] ),
    .I1(_1116_),
    .S(_0963_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3335_ (.I0(_0332_),
    .I1(\add_result[23] ),
    .I2(\add_result[22] ),
    .I3(\add_result[24] ),
    .S0(_0820_),
    .S1(_0366_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3336_ (.I0(_1053_),
    .I1(_1117_),
    .S(_0968_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3337_ (.A1(_1009_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3338_ (.A1(_0902_),
    .A2(_0906_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3339_ (.I0(_1057_),
    .I1(_1120_),
    .S(_0968_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3340_ (.A1(_1021_),
    .A2(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3341_ (.A1(_0902_),
    .A2(_0982_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3342_ (.A1(_1123_),
    .A2(_1016_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3343_ (.A1(_1098_),
    .A2(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _3344_ (.A1(_1008_),
    .A2(_1119_),
    .B1(_1122_),
    .B2(_0886_),
    .C(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3345_ (.A1(_0334_),
    .A2(_1060_),
    .B(\add_result[22] ),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _3346_ (.A1(_0333_),
    .A2(_0332_),
    .A3(\add_result[23] ),
    .B(_0347_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3347_ (.A1(\add_result[23] ),
    .A2(_0344_),
    .B(\add_result[24] ),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _3348_ (.A1(\add_result[24] ),
    .A2(_1127_),
    .A3(_1128_),
    .B(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3349_ (.I0(_1126_),
    .I1(_1130_),
    .S(_0920_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _3350_ (.A1(\add_result[24] ),
    .A2(_0874_),
    .B1(_1131_),
    .B2(_0922_),
    .C(\add_result[26] ),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3351_ (.A1(_0946_),
    .A2(_0327_),
    .B(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3352_ (.I0(\final_mant[22] ),
    .I1(_1133_),
    .S(_0963_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3353_ (.I(\add_result[5] ),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3354_ (.A1(\add_result[2] ),
    .A2(_1711_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3355_ (.I0(\add_result[4] ),
    .I1(\add_result[3] ),
    .S(_1708_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3356_ (.I0(_1135_),
    .I1(_1136_),
    .S(_0914_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3357_ (.A1(_1698_),
    .A2(_0920_),
    .A3(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3358_ (.A1(_0814_),
    .A2(_0891_),
    .A3(_1057_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3359_ (.A1(_1138_),
    .A2(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3360_ (.A1(\add_result[4] ),
    .A2(_0874_),
    .B1(_1140_),
    .B2(_0922_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _3361_ (.A1(_1134_),
    .A2(_0862_),
    .B1(_0354_),
    .B2(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3362_ (.I0(\final_mant[2] ),
    .I1(_1142_),
    .S(_0963_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3363_ (.A1(\add_result[5] ),
    .A2(_0871_),
    .B1(_0891_),
    .B2(_1071_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3364_ (.I0(\add_result[3] ),
    .I1(\add_result[2] ),
    .S(_0353_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3365_ (.I0(\add_result[4] ),
    .I1(\add_result[5] ),
    .S(_0352_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3366_ (.I0(_1144_),
    .I1(_1145_),
    .S(_0914_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3367_ (.A1(_1698_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3368_ (.I0(_1143_),
    .I1(_1147_),
    .S(_0920_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3369_ (.I0(_1134_),
    .I1(_1148_),
    .S(_0342_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3370_ (.A1(\add_result[6] ),
    .A2(_0829_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3371_ (.A1(_0354_),
    .A2(_1149_),
    .B(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3372_ (.I0(\final_mant[3] ),
    .I1(_1151_),
    .S(_0963_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3373_ (.I0(_0912_),
    .I1(_1136_),
    .S(_1702_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3374_ (.A1(_1695_),
    .A2(_1574_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _3375_ (.A1(_1698_),
    .A2(_1152_),
    .B1(_1153_),
    .B2(_1135_),
    .C(_0814_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3376_ (.A1(_1098_),
    .A2(_1154_),
    .B(_0922_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3377_ (.A1(_0929_),
    .A2(_1091_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3378_ (.A1(_0814_),
    .A2(_1156_),
    .B(_1154_),
    .C(_0328_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3379_ (.A1(\add_result[6] ),
    .A2(_1155_),
    .B(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3380_ (.A1(\add_result[7] ),
    .A2(_0829_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3381_ (.A1(_0354_),
    .A2(_1158_),
    .B(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3382_ (.I0(\final_mant[4] ),
    .I1(_1160_),
    .S(_0963_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3383_ (.I0(_0938_),
    .I1(_1145_),
    .S(_1702_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3384_ (.A1(_1574_),
    .A2(_1144_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3385_ (.I0(_1161_),
    .I1(_1162_),
    .S(_1695_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3386_ (.A1(_0877_),
    .A2(_1037_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3387_ (.I0(\add_result[3] ),
    .I1(\add_result[7] ),
    .I2(\add_result[2] ),
    .I3(\add_result[6] ),
    .S0(_0968_),
    .S1(_1707_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3388_ (.I0(_1164_),
    .I1(_1165_),
    .S(_0821_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3389_ (.A1(_0929_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3390_ (.I0(_1163_),
    .I1(_1167_),
    .S(_0814_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3391_ (.A1(\add_result[7] ),
    .A2(_0874_),
    .B1(_1168_),
    .B2(_0922_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3392_ (.A1(\add_result[8] ),
    .A2(_0829_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3393_ (.A1(_0354_),
    .A2(_1169_),
    .B(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3394_ (.I0(\final_mant[5] ),
    .I1(_1171_),
    .S(_0963_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3395_ (.A1(_0929_),
    .A2(_1121_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3396_ (.I0(_0915_),
    .I1(_1137_),
    .S(_1695_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3397_ (.I0(_1172_),
    .I1(_1173_),
    .S(_0920_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3398_ (.A1(\add_result[8] ),
    .A2(_0874_),
    .B1(_1174_),
    .B2(_0922_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3399_ (.A1(\add_result[9] ),
    .A2(_0829_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3400_ (.A1(_0354_),
    .A2(_1175_),
    .B(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3401_ (.I0(\final_mant[6] ),
    .I1(_1177_),
    .S(net66),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3402_ (.A1(_0902_),
    .A2(_0932_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3403_ (.I0(_1071_),
    .I1(_1178_),
    .S(_0877_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3404_ (.A1(_0929_),
    .A2(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3405_ (.I0(_0940_),
    .I1(_1146_),
    .S(_1695_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3406_ (.I0(_1180_),
    .I1(_1181_),
    .S(_0920_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3407_ (.A1(\add_result[9] ),
    .A2(_0874_),
    .B1(_1182_),
    .B2(_0922_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3408_ (.A1(\add_result[10] ),
    .A2(_0829_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3409_ (.A1(_0354_),
    .A2(_1183_),
    .B(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3410_ (.I0(\final_mant[7] ),
    .I1(_1185_),
    .S(net66),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3411_ (.I(\add_result[11] ),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3412_ (.A1(_0929_),
    .A2(_0903_),
    .A3(_1019_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3413_ (.I0(_0955_),
    .I1(_1152_),
    .S(_1695_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3414_ (.I0(_1187_),
    .I1(_1188_),
    .S(_0363_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3415_ (.A1(\add_result[10] ),
    .A2(_0875_),
    .B1(_1189_),
    .B2(_0946_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3416_ (.I0(_1186_),
    .I1(_1190_),
    .S(_0862_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3417_ (.A1(_0926_),
    .A2(\final_mant[8] ),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3418_ (.A1(_0927_),
    .A2(_1191_),
    .B(_1192_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3419_ (.I(\add_result[12] ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3420_ (.A1(_0929_),
    .A2(_0903_),
    .A3(_1039_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3421_ (.I0(_0971_),
    .I1(_1161_),
    .S(_1695_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3422_ (.I0(_1194_),
    .I1(_1195_),
    .S(_0363_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3423_ (.A1(\add_result[11] ),
    .A2(_0875_),
    .B1(_1196_),
    .B2(_0946_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3424_ (.I0(_1193_),
    .I1(_1197_),
    .S(_0343_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3425_ (.A1(_0926_),
    .A2(\final_mant[9] ),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3426_ (.A1(_0927_),
    .A2(_1198_),
    .B(_1199_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3427_ (.A1(_1578_),
    .A2(_0806_),
    .B(_0298_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3428_ (.A1(_0801_),
    .A2(_0806_),
    .B(invalid_op_stage2),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3429_ (.A1(_0372_),
    .A2(_1200_),
    .B(_1201_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3430_ (.A1(\aligned_a_mant[1] ),
    .A2(\aligned_a_mant[0] ),
    .A3(\aligned_b_mant[1] ),
    .A4(\aligned_b_mant[0] ),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3431_ (.A1(net22),
    .A2(net21),
    .A3(net25),
    .A4(net23),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3432_ (.A1(net18),
    .A2(net17),
    .A3(net20),
    .A4(net19),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3433_ (.A1(_1202_),
    .A2(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3434_ (.A1(net13),
    .A2(net2),
    .A3(net27),
    .A4(net16),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3435_ (.A1(net9),
    .A2(net11),
    .A3(net15),
    .A4(net14),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3436_ (.A1(net3),
    .A2(net7),
    .A3(net10),
    .A4(net12),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3437_ (.A1(net6),
    .A2(net5),
    .A3(net8),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3438_ (.A1(_1205_),
    .A2(_1206_),
    .A3(_1207_),
    .A4(_1208_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3439_ (.A1(net28),
    .A2(net30),
    .A3(net33),
    .A4(net32),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3440_ (.A1(net24),
    .A2(net29),
    .A3(net31),
    .A4(net4),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _3441_ (.A1(_1204_),
    .A2(_1209_),
    .A3(_1210_),
    .A4(_1211_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3442_ (.A1(net54),
    .A2(net53),
    .A3(net57),
    .A4(net55),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3443_ (.A1(net50),
    .A2(net49),
    .A3(net52),
    .A4(net51),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3444_ (.A1(_1213_),
    .A2(_1214_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3445_ (.A1(net45),
    .A2(net34),
    .A3(net59),
    .A4(net48),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3446_ (.A1(net41),
    .A2(net43),
    .A3(net47),
    .A4(net46),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3447_ (.A1(net35),
    .A2(net39),
    .A3(net42),
    .A4(net44),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3448_ (.A1(net38),
    .A2(net37),
    .A3(net40),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3449_ (.A1(_1216_),
    .A2(_1217_),
    .A3(_1218_),
    .A4(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3450_ (.A1(net60),
    .A2(net62),
    .A3(net65),
    .A4(net64),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3451_ (.A1(net56),
    .A2(net61),
    .A3(net63),
    .A4(net36),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3452_ (.A1(_1215_),
    .A2(_1220_),
    .A3(_1221_),
    .A4(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3453_ (.I(_1581_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3454_ (.I(_1611_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3455_ (.I(_1616_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3456_ (.A1(_1611_),
    .A2(_1617_),
    .B(_1613_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _3457_ (.A1(_1225_),
    .A2(_1689_),
    .A3(_1226_),
    .B(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3458_ (.I(_1587_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3459_ (.A1(_1599_),
    .A2(_1605_),
    .A3(_1593_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3460_ (.A1(_1229_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3461_ (.I(_1599_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3462_ (.A1(_1232_),
    .A2(_1593_),
    .A3(_1607_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3463_ (.A1(_1593_),
    .A2(_1601_),
    .B(_1595_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3464_ (.A1(_1233_),
    .A2(_1234_),
    .B(_1229_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _3465_ (.A1(_1228_),
    .A2(_1231_),
    .B(_1235_),
    .C(_1589_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3466_ (.A1(_1587_),
    .A2(_1599_),
    .A3(_1581_),
    .A4(_1593_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3467_ (.A1(_1611_),
    .A2(_1605_),
    .A3(_1690_),
    .A4(_1616_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3468_ (.A1(_1237_),
    .A2(_1238_),
    .B(_1583_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3469_ (.A1(_1224_),
    .A2(_1236_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3470_ (.A1(_1669_),
    .A2(_1668_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3471_ (.A1(_1687_),
    .A2(_1681_),
    .A3(_1684_),
    .A4(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3472_ (.I(_1681_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3473_ (.A1(_1684_),
    .A2(_1686_),
    .B(_1683_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _3474_ (.A1(_1243_),
    .A2(_1244_),
    .B(_1238_),
    .C(_1237_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3475_ (.A1(_1680_),
    .A2(_1242_),
    .A3(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3476_ (.A1(_1240_),
    .A2(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3477_ (.A1(_1635_),
    .A2(_1638_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3478_ (.I(_1623_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _3479_ (.A1(_1249_),
    .A2(_1624_),
    .B(_1630_),
    .C(_1621_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3480_ (.A1(_1620_),
    .A2(_1630_),
    .B(_1629_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3481_ (.A1(_1627_),
    .A2(_1639_),
    .A3(_1642_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3482_ (.A1(_1250_),
    .A2(_1251_),
    .B(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3483_ (.A1(_1626_),
    .A2(_1642_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3484_ (.A1(_1641_),
    .A2(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3485_ (.A1(_1639_),
    .A2(_1255_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3486_ (.A1(_1645_),
    .A2(_1672_),
    .A3(_1675_),
    .A4(_1678_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3487_ (.A1(_1648_),
    .A2(_1651_),
    .A3(_1654_),
    .A4(_1657_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3488_ (.A1(_1257_),
    .A2(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3489_ (.A1(_1633_),
    .A2(_1660_),
    .A3(_1663_),
    .A4(_1666_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3490_ (.A1(_1636_),
    .A2(_1635_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3491_ (.A1(_1259_),
    .A2(_1260_),
    .A3(_1261_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _3492_ (.A1(_1248_),
    .A2(_1253_),
    .A3(_1256_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3493_ (.A1(_1648_),
    .A2(_1651_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3494_ (.A1(_1656_),
    .A2(_1654_),
    .B(_1653_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3495_ (.A1(_1648_),
    .A2(_1650_),
    .B(_1647_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3496_ (.A1(_1264_),
    .A2(_1265_),
    .B(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3497_ (.A1(_1257_),
    .A2(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3498_ (.A1(_1660_),
    .A2(_1663_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3499_ (.A1(_1632_),
    .A2(_1666_),
    .B(_1665_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3500_ (.A1(_1662_),
    .A2(_1660_),
    .B(_1659_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3501_ (.A1(_1269_),
    .A2(_1270_),
    .B(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3502_ (.A1(_1259_),
    .A2(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3503_ (.A1(_1687_),
    .A2(_1681_),
    .A3(_1684_),
    .A4(_1668_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3504_ (.A1(_1671_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3505_ (.I(_1675_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3506_ (.A1(_1644_),
    .A2(_1678_),
    .B(_1677_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3507_ (.I(_1674_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3508_ (.A1(_1276_),
    .A2(_1277_),
    .B(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3509_ (.A1(_1672_),
    .A2(_1279_),
    .B(_1245_),
    .C(_1680_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3510_ (.A1(_1268_),
    .A2(_1273_),
    .A3(_1275_),
    .A4(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3511_ (.A1(_1263_),
    .A2(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _3512_ (.A1(_1247_),
    .A2(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3513_ (.I(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _3514_ (.A1(_1223_),
    .A2(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _3515_ (.A1(_1212_),
    .A2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3516_ (.I(_1286_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3517_ (.I0(net17),
    .I1(net49),
    .S(_1287_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3518_ (.I0(net18),
    .I1(net50),
    .S(_1287_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3519_ (.I0(net19),
    .I1(net51),
    .S(_1286_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3520_ (.I0(net20),
    .I1(net52),
    .S(_1286_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3521_ (.I0(net21),
    .I1(net53),
    .S(_1286_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3522_ (.I0(net22),
    .I1(net54),
    .S(_1286_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3523_ (.I0(net23),
    .I1(net55),
    .S(_1286_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3524_ (.I0(net25),
    .I1(net57),
    .S(_1286_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3525_ (.I(net2),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3526_ (.I(net45),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3527_ (.I(net56),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3528_ (.I(net59),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3529_ (.I(net60),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3530_ (.I(net61),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3531_ (.I(net62),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3532_ (.I(net63),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3533_ (.I(net64),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3534_ (.I(net65),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3535_ (.I(net35),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3536_ (.I(net36),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3537_ (.I(net37),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3538_ (.I(net38),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3539_ (.I(net39),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3540_ (.I(net40),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3541_ (.I(net41),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3542_ (.I(net42),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3543_ (.I(net43),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3544_ (.I(net44),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3545_ (.I(net46),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3546_ (.I(net47),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3547_ (.I(net48),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _3548_ (.I(_1690_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3549_ (.I(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3550_ (.I(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3551_ (.I(_1247_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3552_ (.I(_1282_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3553_ (.A1(_1593_),
    .A2(_1598_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3554_ (.A1(_1232_),
    .A2(_1593_),
    .A3(_1604_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3555_ (.A1(_1611_),
    .A2(_1567_),
    .B(_1610_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3556_ (.A1(_1230_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3557_ (.A1(_1592_),
    .A2(_1293_),
    .A3(_1294_),
    .A4(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3558_ (.A1(_1587_),
    .A2(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3559_ (.A1(_1229_),
    .A2(_1230_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3560_ (.I(_1692_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3561_ (.A1(_1566_),
    .A2(_1616_),
    .B(_1610_),
    .C(_1615_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3562_ (.A1(_1611_),
    .A2(_1610_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _3563_ (.A1(_1592_),
    .A2(_1293_),
    .A3(_1294_),
    .B(_1587_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _3564_ (.A1(_1299_),
    .A2(_1300_),
    .A3(_1301_),
    .B(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3565_ (.A1(_1224_),
    .A2(_1586_),
    .A3(_1303_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3566_ (.A1(_1586_),
    .A2(_1592_),
    .A3(_1293_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _3567_ (.A1(_1587_),
    .A2(_1586_),
    .B(_1305_),
    .C(_1581_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3568_ (.I(_1605_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3569_ (.I(_1604_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3570_ (.A1(_1307_),
    .A2(_1295_),
    .B(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3571_ (.A1(_1237_),
    .A2(_1309_),
    .B(_1580_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3572_ (.A1(_1224_),
    .A2(_1586_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _3573_ (.A1(_1224_),
    .A2(_1303_),
    .B1(_1306_),
    .B2(_1310_),
    .C(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3574_ (.A1(_1298_),
    .A2(_1304_),
    .A3(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _3575_ (.A1(_1291_),
    .A2(_1292_),
    .B(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3576_ (.I(_1568_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _3577_ (.I(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3578_ (.A1(_1610_),
    .A2(_1615_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3579_ (.A1(_1692_),
    .A2(_1226_),
    .B(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3580_ (.A1(_1611_),
    .A2(_1610_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3581_ (.A1(_1605_),
    .A2(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3582_ (.A1(_1318_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3583_ (.I(_1593_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3584_ (.A1(_1322_),
    .A2(_1598_),
    .A3(_1604_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3585_ (.A1(_1232_),
    .A2(_1322_),
    .A3(_1318_),
    .A4(_1320_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3586_ (.A1(_1232_),
    .A2(_1322_),
    .A3(_1604_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _3587_ (.A(_1565_),
    .B(net50),
    .CI(_1566_),
    .CO(_1567_),
    .S(_1568_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _3588_ (.A(net18),
    .B(_1569_),
    .CI(_1570_),
    .CO(_1571_),
    .S(_1572_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _3589_ (.A(\result_exp_stage2[1] ),
    .B(_1573_),
    .CI(_1574_),
    .CO(_1575_),
    .S(_1576_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3590_ (.A(net26),
    .B(net58),
    .CO(_1577_),
    .S(_1578_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3591_ (.A(_1579_),
    .B(net57),
    .CO(_1580_),
    .S(_1581_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3592_ (.A(net25),
    .B(_1582_),
    .CO(_1583_),
    .S(_1584_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3593_ (.A(_1585_),
    .B(net55),
    .CO(_1586_),
    .S(_1587_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3594_ (.A(net23),
    .B(_1588_),
    .CO(_1589_),
    .S(_1590_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3595_ (.A(_1591_),
    .B(net54),
    .CO(_1592_),
    .S(_1593_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3596_ (.A(net22),
    .B(_1594_),
    .CO(_1595_),
    .S(_1596_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3597_ (.A(_1597_),
    .B(net53),
    .CO(_1598_),
    .S(_1599_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3598_ (.A(net21),
    .B(_1600_),
    .CO(_1601_),
    .S(_1602_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3599_ (.A(_1603_),
    .B(net52),
    .CO(_1604_),
    .S(_1605_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3600_ (.A(net20),
    .B(_1606_),
    .CO(_1607_),
    .S(_1608_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3601_ (.A(_1609_),
    .B(net51),
    .CO(_1610_),
    .S(_1611_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3602_ (.A(net19),
    .B(_1612_),
    .CO(_1613_),
    .S(_1614_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3603_ (.A(_1565_),
    .B(net50),
    .CO(_1615_),
    .S(_1616_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3604_ (.A(net18),
    .B(_1569_),
    .CO(_1617_),
    .S(_1618_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3605_ (.A(net13),
    .B(_1619_),
    .CO(_1620_),
    .S(_1621_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3606_ (.A(_1622_),
    .B(net34),
    .CO(_1623_),
    .S(_1624_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3607_ (.A(net27),
    .B(_1625_),
    .CO(_1626_),
    .S(_1627_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3608_ (.A(net24),
    .B(_1628_),
    .CO(_1629_),
    .S(_1630_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3609_ (.A(net31),
    .B(_1631_),
    .CO(_1632_),
    .S(_1633_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3610_ (.A(net30),
    .B(_1634_),
    .CO(_1635_),
    .S(_1636_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3611_ (.A(net29),
    .B(_1637_),
    .CO(_1638_),
    .S(_1639_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3612_ (.A(net28),
    .B(_1640_),
    .CO(_1641_),
    .S(_1642_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3613_ (.A(net8),
    .B(_1643_),
    .CO(_1644_),
    .S(_1645_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3614_ (.A(net7),
    .B(_1646_),
    .CO(_1647_),
    .S(_1648_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3615_ (.A(net6),
    .B(_1649_),
    .CO(_1650_),
    .S(_1651_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3616_ (.A(net5),
    .B(_1652_),
    .CO(_1653_),
    .S(_1654_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3617_ (.A(net4),
    .B(_1655_),
    .CO(_1656_),
    .S(_1657_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3618_ (.A(net3),
    .B(_1658_),
    .CO(_1659_),
    .S(_1660_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3619_ (.A(net33),
    .B(_1661_),
    .CO(_1662_),
    .S(_1663_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3620_ (.A(net32),
    .B(_1664_),
    .CO(_1665_),
    .S(_1666_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3621_ (.A(net12),
    .B(_1667_),
    .CO(_1668_),
    .S(_1669_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3622_ (.A(net11),
    .B(_1670_),
    .CO(_1671_),
    .S(_1672_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3623_ (.A(net10),
    .B(_1673_),
    .CO(_1674_),
    .S(_1675_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3624_ (.A(net9),
    .B(_1676_),
    .CO(_1677_),
    .S(_1678_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3625_ (.A(net16),
    .B(_1679_),
    .CO(_1680_),
    .S(_1681_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3626_ (.A(net15),
    .B(_1682_),
    .CO(_1683_),
    .S(_1684_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3627_ (.A(net14),
    .B(_1685_),
    .CO(_1686_),
    .S(_1687_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3628_ (.A(_1688_),
    .B(net49),
    .CO(_1689_),
    .S(_1690_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3629_ (.A(net17),
    .B(_1691_),
    .CO(_1692_),
    .S(_1693_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3630_ (.A(_1694_),
    .B(_1695_),
    .CO(_1696_),
    .S(_1697_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3631_ (.A(\result_exp_stage2[2] ),
    .B(_1698_),
    .CO(_1699_),
    .S(_1700_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3632_ (.A(_1701_),
    .B(_1702_),
    .CO(_1703_),
    .S(_1704_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3633_ (.A(\result_exp_stage2[1] ),
    .B(_1574_),
    .CO(_1705_),
    .S(_1706_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3634_ (.A(_1707_),
    .B(_1708_),
    .CO(_1709_),
    .S(_1710_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3635_ (.A(\result_exp_stage2[0] ),
    .B(_1711_),
    .CO(_1712_),
    .S(_1713_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3636_ (.A(_1707_),
    .B(_1701_),
    .CO(_1714_),
    .S(_1715_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3637_ (.A(_1707_),
    .B(\result_exp_stage2[1] ),
    .CO(_1716_),
    .S(_1717_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3638_ (.A(\result_exp_stage2[0] ),
    .B(\result_exp_stage2[1] ),
    .CO(_1718_),
    .S(_1719_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3639_ (.A(_1720_),
    .B(\aligned_b_mant[2] ),
    .CO(_1721_),
    .S(_1722_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3640_ (.A(\aligned_a_mant[2] ),
    .B(_1723_),
    .CO(_1724_),
    .S(_1725_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3641_ (.A(\aligned_a_mant[2] ),
    .B(\aligned_b_mant[2] ),
    .CO(_1726_),
    .S(_1727_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3642_ (.A(_1728_),
    .B(\aligned_b_mant[1] ),
    .CO(_1729_),
    .S(_1730_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3643_ (.A(\aligned_a_mant[1] ),
    .B(_1731_),
    .CO(_1732_),
    .S(_1733_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3644_ (.A(\aligned_a_mant[1] ),
    .B(\aligned_b_mant[1] ),
    .CO(_1734_),
    .S(_1735_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3645_ (.A(_1736_),
    .B(\aligned_b_mant[3] ),
    .CO(_1737_),
    .S(_1738_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3646_ (.A(\aligned_a_mant[3] ),
    .B(_1739_),
    .CO(_1740_),
    .S(_1741_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3647_ (.A(\aligned_a_mant[3] ),
    .B(\aligned_b_mant[3] ),
    .CO(_1742_),
    .S(_1743_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3648_ (.A(_1744_),
    .B(\aligned_b_mant[4] ),
    .CO(_1745_),
    .S(_1746_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3649_ (.A(\aligned_a_mant[4] ),
    .B(_1747_),
    .CO(_1748_),
    .S(_1749_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3650_ (.A(\aligned_a_mant[4] ),
    .B(\aligned_b_mant[4] ),
    .CO(_1750_),
    .S(_1751_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3651_ (.A(_1752_),
    .B(\aligned_b_mant[5] ),
    .CO(_1753_),
    .S(_1754_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3652_ (.A(\aligned_a_mant[5] ),
    .B(_1755_),
    .CO(_1756_),
    .S(_1757_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3653_ (.A(\aligned_a_mant[5] ),
    .B(\aligned_b_mant[5] ),
    .CO(_1758_),
    .S(_1759_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3654_ (.A(_1760_),
    .B(\aligned_b_mant[6] ),
    .CO(_1761_),
    .S(_1762_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3655_ (.A(\aligned_a_mant[6] ),
    .B(_1763_),
    .CO(_1764_),
    .S(_1765_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3656_ (.A(\aligned_a_mant[6] ),
    .B(\aligned_b_mant[6] ),
    .CO(_1766_),
    .S(_1767_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3657_ (.A(_1768_),
    .B(\aligned_b_mant[7] ),
    .CO(_1769_),
    .S(_1770_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3658_ (.A(\aligned_a_mant[7] ),
    .B(_1771_),
    .CO(_1772_),
    .S(_1773_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3659_ (.A(\aligned_a_mant[7] ),
    .B(\aligned_b_mant[7] ),
    .CO(_1774_),
    .S(_1775_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3660_ (.A(_1776_),
    .B(\aligned_b_mant[8] ),
    .CO(_1777_),
    .S(_1778_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3661_ (.A(\aligned_a_mant[8] ),
    .B(_1779_),
    .CO(_1780_),
    .S(_1781_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3662_ (.A(\aligned_a_mant[8] ),
    .B(\aligned_b_mant[8] ),
    .CO(_1782_),
    .S(_1783_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3663_ (.A(_1784_),
    .B(\aligned_b_mant[9] ),
    .CO(_1785_),
    .S(_1786_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3664_ (.A(\aligned_a_mant[9] ),
    .B(_1787_),
    .CO(_1788_),
    .S(_1789_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3665_ (.A(\aligned_a_mant[9] ),
    .B(\aligned_b_mant[9] ),
    .CO(_1790_),
    .S(_1791_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3666_ (.A(_1792_),
    .B(\aligned_b_mant[10] ),
    .CO(_1793_),
    .S(_1794_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3667_ (.A(\aligned_a_mant[10] ),
    .B(_1795_),
    .CO(_1796_),
    .S(_1797_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3668_ (.A(\aligned_a_mant[10] ),
    .B(\aligned_b_mant[10] ),
    .CO(_1798_),
    .S(_1799_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3669_ (.A(_1800_),
    .B(\aligned_b_mant[11] ),
    .CO(_1801_),
    .S(_1802_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3670_ (.A(\aligned_a_mant[11] ),
    .B(_1803_),
    .CO(_1804_),
    .S(_1805_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3671_ (.A(\aligned_a_mant[11] ),
    .B(\aligned_b_mant[11] ),
    .CO(_1806_),
    .S(_1807_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3672_ (.A(_1808_),
    .B(\aligned_b_mant[12] ),
    .CO(_1809_),
    .S(_1810_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3673_ (.A(\aligned_a_mant[12] ),
    .B(_1811_),
    .CO(_1812_),
    .S(_1813_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3674_ (.A(\aligned_a_mant[12] ),
    .B(\aligned_b_mant[12] ),
    .CO(_1814_),
    .S(_1815_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3675_ (.A(_1816_),
    .B(\aligned_b_mant[13] ),
    .CO(_1817_),
    .S(_1818_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3676_ (.A(\aligned_a_mant[13] ),
    .B(_1819_),
    .CO(_1820_),
    .S(_1821_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3677_ (.A(\aligned_a_mant[13] ),
    .B(\aligned_b_mant[13] ),
    .CO(_1822_),
    .S(_1823_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3678_ (.A(_1824_),
    .B(\aligned_b_mant[14] ),
    .CO(_1825_),
    .S(_1826_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3679_ (.A(\aligned_a_mant[14] ),
    .B(_1827_),
    .CO(_1828_),
    .S(_1829_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3680_ (.A(\aligned_a_mant[14] ),
    .B(\aligned_b_mant[14] ),
    .CO(_1830_),
    .S(_1831_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3681_ (.A(_1832_),
    .B(\aligned_b_mant[15] ),
    .CO(_1833_),
    .S(_1834_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3682_ (.A(\aligned_a_mant[15] ),
    .B(_1835_),
    .CO(_1836_),
    .S(_1837_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3683_ (.A(\aligned_a_mant[15] ),
    .B(\aligned_b_mant[15] ),
    .CO(_1838_),
    .S(_1839_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3684_ (.A(_1840_),
    .B(\aligned_b_mant[16] ),
    .CO(_1841_),
    .S(_1842_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3685_ (.A(\aligned_a_mant[16] ),
    .B(_1843_),
    .CO(_1844_),
    .S(_1845_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3686_ (.A(\aligned_a_mant[16] ),
    .B(\aligned_b_mant[16] ),
    .CO(_1846_),
    .S(_1847_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3687_ (.A(_1848_),
    .B(\aligned_b_mant[17] ),
    .CO(_1849_),
    .S(_1850_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3688_ (.A(\aligned_a_mant[17] ),
    .B(_1851_),
    .CO(_1852_),
    .S(_1853_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3689_ (.A(\aligned_a_mant[17] ),
    .B(\aligned_b_mant[17] ),
    .CO(_1854_),
    .S(_1855_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3690_ (.A(_1856_),
    .B(\aligned_b_mant[18] ),
    .CO(_1857_),
    .S(_1858_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3691_ (.A(\aligned_a_mant[18] ),
    .B(_1859_),
    .CO(_1860_),
    .S(_1861_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3692_ (.A(\aligned_a_mant[18] ),
    .B(\aligned_b_mant[18] ),
    .CO(_1862_),
    .S(_1863_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3693_ (.A(_1864_),
    .B(\aligned_b_mant[19] ),
    .CO(_1865_),
    .S(_1866_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3694_ (.A(\aligned_a_mant[19] ),
    .B(_1867_),
    .CO(_1868_),
    .S(_1869_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3695_ (.A(\aligned_a_mant[19] ),
    .B(\aligned_b_mant[19] ),
    .CO(_1870_),
    .S(_1871_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3696_ (.A(_1872_),
    .B(\aligned_b_mant[20] ),
    .CO(_1873_),
    .S(_1874_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3697_ (.A(\aligned_a_mant[20] ),
    .B(_1875_),
    .CO(_1876_),
    .S(_1877_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3698_ (.A(\aligned_a_mant[20] ),
    .B(\aligned_b_mant[20] ),
    .CO(_1878_),
    .S(_1879_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3699_ (.A(_1880_),
    .B(\aligned_b_mant[21] ),
    .CO(_1881_),
    .S(_1882_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3700_ (.A(\aligned_a_mant[21] ),
    .B(_1883_),
    .CO(_1884_),
    .S(_1885_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3701_ (.A(\aligned_a_mant[21] ),
    .B(\aligned_b_mant[21] ),
    .CO(_1886_),
    .S(_1887_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3702_ (.A(_1888_),
    .B(\aligned_b_mant[22] ),
    .CO(_1889_),
    .S(_1890_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3703_ (.A(\aligned_a_mant[22] ),
    .B(_1891_),
    .CO(_1892_),
    .S(_1893_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3704_ (.A(\aligned_a_mant[22] ),
    .B(\aligned_b_mant[22] ),
    .CO(_1894_),
    .S(_1895_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3705_ (.A(_1896_),
    .B(\aligned_b_mant[23] ),
    .CO(_1897_),
    .S(_1898_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3706_ (.A(\aligned_a_mant[23] ),
    .B(_1899_),
    .CO(_1900_),
    .S(_1901_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3707_ (.A(\aligned_a_mant[23] ),
    .B(\aligned_b_mant[23] ),
    .CO(_1902_),
    .S(_1903_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3708_ (.A(_1904_),
    .B(\aligned_b_mant[24] ),
    .CO(_1905_),
    .S(_1906_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3709_ (.A(\aligned_a_mant[24] ),
    .B(_1907_),
    .CO(_1908_),
    .S(_1909_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3710_ (.A(\aligned_a_mant[24] ),
    .B(\aligned_b_mant[24] ),
    .CO(_1910_),
    .S(_1911_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3711_ (.A(_1912_),
    .B(\aligned_b_mant[25] ),
    .CO(_1913_),
    .S(_1914_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3712_ (.A(\aligned_a_mant[25] ),
    .B(_1915_),
    .CO(_1916_),
    .S(_1917_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3713_ (.A(\aligned_a_mant[25] ),
    .B(\aligned_b_mant[25] ),
    .CO(_1918_),
    .S(_1919_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \a_sign_stage1$_DFF_PN0_  (.D(net26),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(a_sign_stage1));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[10]$_DFF_PN0_  (.D(_0000_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\add_result[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[11]$_DFF_PN0_  (.D(_0001_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\add_result[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[12]$_DFF_PN0_  (.D(_0002_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\add_result[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[13]$_DFF_PN0_  (.D(_0003_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\add_result[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[14]$_DFF_PN0_  (.D(_0004_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\add_result[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[15]$_DFF_PN0_  (.D(_0005_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\add_result[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[16]$_DFF_PN0_  (.D(_0006_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\add_result[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[17]$_DFF_PN0_  (.D(_0007_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[18]$_DFF_PN0_  (.D(_0008_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[19]$_DFF_PN0_  (.D(_0009_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[20]$_DFF_PN0_  (.D(_0010_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\add_result[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[21]$_DFF_PN0_  (.D(_0011_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[22]$_DFF_PN0_  (.D(_0012_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[23]$_DFF_PN0_  (.D(_0013_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[24]$_DFF_PN0_  (.D(_0014_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[25]$_DFF_PN0_  (.D(_0015_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[26]$_DFF_PN0_  (.D(_0016_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\add_result[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[2]$_DFF_PN0_  (.D(_0017_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\add_result[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[3]$_DFF_PN0_  (.D(_0018_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\add_result[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[4]$_DFF_PN0_  (.D(_0019_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\add_result[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[5]$_DFF_PN0_  (.D(_0020_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\add_result[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[6]$_DFF_PN0_  (.D(_0021_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\add_result[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[7]$_DFF_PN0_  (.D(_0022_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\add_result[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \add_result[8]$_DFF_PN0_  (.D(_0023_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\add_result[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \add_result[9]$_DFF_PN0_  (.D(_0024_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\add_result[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[0]$_DFF_PN0_  (.D(_0025_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[10]$_DFF_PN0_  (.D(_0026_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[11]$_DFF_PN0_  (.D(_0027_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[12]$_DFF_PN0_  (.D(_0028_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_a_mant[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[13]$_DFF_PN0_  (.D(_0029_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\aligned_a_mant[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[14]$_DFF_PN0_  (.D(_0030_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_a_mant[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[15]$_DFF_PN0_  (.D(_0031_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\aligned_a_mant[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[16]$_DFF_PN0_  (.D(_0032_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_a_mant[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[17]$_DFF_PN0_  (.D(_0033_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[18]$_DFF_PN0_  (.D(_0034_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[19]$_DFF_PN0_  (.D(_0035_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[1]$_DFF_PN0_  (.D(_0036_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[20]$_DFF_PN0_  (.D(_0037_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[21]$_DFF_PN0_  (.D(_0038_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[22]$_DFF_PN0_  (.D(_0039_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_a_mant[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[23]$_DFF_PN0_  (.D(_0040_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_a_mant[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[24]$_DFF_PN0_  (.D(_0041_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_a_mant[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[25]$_DFF_PN0_  (.D(_0042_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\aligned_a_mant[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[2]$_DFF_PN0_  (.D(_0043_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[3]$_DFF_PN0_  (.D(_0044_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[4]$_DFF_PN0_  (.D(_0045_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[5]$_DFF_PN0_  (.D(_0046_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[6]$_DFF_PN0_  (.D(_0047_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[7]$_DFF_PN0_  (.D(_0048_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[8]$_DFF_PN0_  (.D(_0049_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_a_mant[9]$_DFF_PN0_  (.D(_0050_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[0]$_DFF_PN0_  (.D(_0051_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_b_mant[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[10]$_DFF_PN0_  (.D(_0052_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[11]$_DFF_PN0_  (.D(_0053_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[12]$_DFF_PN0_  (.D(_0054_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_b_mant[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[13]$_DFF_PN0_  (.D(_0055_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[14]$_DFF_PN0_  (.D(_0056_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_b_mant[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[15]$_DFF_PN0_  (.D(_0057_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[16]$_DFF_PN0_  (.D(_0058_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\aligned_b_mant[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[17]$_DFF_PN0_  (.D(_0059_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\aligned_b_mant[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[18]$_DFF_PN0_  (.D(_0060_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[19]$_DFF_PN0_  (.D(_0061_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[1]$_DFF_PN0_  (.D(_0062_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[20]$_DFF_PN0_  (.D(_0063_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[21]$_DFF_PN0_  (.D(_0064_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[22]$_DFF_PN0_  (.D(_0065_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[23]$_DFF_PN0_  (.D(_0066_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[24]$_DFF_PN0_  (.D(_0067_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[25]$_DFF_PN0_  (.D(_0068_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[2]$_DFF_PN0_  (.D(_0069_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[3]$_DFF_PN0_  (.D(_0070_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[4]$_DFF_PN0_  (.D(_0071_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[5]$_DFF_PN0_  (.D(_0072_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[6]$_DFF_PN0_  (.D(_0073_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[7]$_DFF_PN0_  (.D(_0074_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[8]$_DFF_PN0_  (.D(_0075_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\aligned_b_mant[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \aligned_b_mant[9]$_DFF_PN0_  (.D(_0076_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \b_sign_stage1$_DFF_PN0_  (.D(net58),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(b_sign_stage1));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[0]$_DFFE_PP_  (.D(_0090_),
    .CLK(clknet_4_1_0_clk),
    .Q(\final_exp[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[1]$_DFFE_PP_  (.D(_0091_),
    .CLK(clknet_4_1_0_clk),
    .Q(\final_exp[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[2]$_DFFE_PP_  (.D(_0092_),
    .CLK(clknet_4_1_0_clk),
    .Q(\final_exp[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[3]$_DFFE_PP_  (.D(_0093_),
    .CLK(clknet_4_1_0_clk),
    .Q(\final_exp[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[4]$_DFFE_PP_  (.D(_0094_),
    .CLK(clknet_4_0_0_clk),
    .Q(\final_exp[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[5]$_DFFE_PP_  (.D(_0095_),
    .CLK(clknet_4_0_0_clk),
    .Q(\final_exp[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[6]$_DFFE_PP_  (.D(_0096_),
    .CLK(clknet_4_0_0_clk),
    .Q(\final_exp[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_exp[7]$_DFFE_PP_  (.D(_0097_),
    .CLK(clknet_4_1_0_clk),
    .Q(\final_exp[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[0]$_DFFE_PP_  (.D(_0098_),
    .CLK(clknet_4_4_0_clk),
    .Q(\final_mant[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[10]$_DFFE_PP_  (.D(_0099_),
    .CLK(clknet_4_4_0_clk),
    .Q(\final_mant[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[11]$_DFFE_PP_  (.D(_0100_),
    .CLK(clknet_4_12_0_clk),
    .Q(\final_mant[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[12]$_DFFE_PP_  (.D(_0101_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[13]$_DFFE_PP_  (.D(_0102_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[14]$_DFFE_PP_  (.D(_0103_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[15]$_DFFE_PP_  (.D(_0104_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[16]$_DFFE_PP_  (.D(_0105_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[17]$_DFFE_PP_  (.D(_0106_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[18]$_DFFE_PP_  (.D(_0107_),
    .CLK(clknet_4_6_0_clk),
    .Q(\final_mant[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[19]$_DFFE_PP_  (.D(_0108_),
    .CLK(clknet_4_6_0_clk),
    .Q(\final_mant[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[1]$_DFFE_PP_  (.D(_0109_),
    .CLK(clknet_4_5_0_clk),
    .Q(\final_mant[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[20]$_DFFE_PP_  (.D(_0110_),
    .CLK(clknet_4_7_0_clk),
    .Q(\final_mant[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[21]$_DFFE_PP_  (.D(_0111_),
    .CLK(clknet_4_6_0_clk),
    .Q(\final_mant[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[22]$_DFFE_PP_  (.D(_0112_),
    .CLK(clknet_4_6_0_clk),
    .Q(\final_mant[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[2]$_DFFE_PP_  (.D(_0113_),
    .CLK(clknet_4_5_0_clk),
    .Q(\final_mant[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[3]$_DFFE_PP_  (.D(_0114_),
    .CLK(clknet_4_4_0_clk),
    .Q(\final_mant[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[4]$_DFFE_PP_  (.D(_0115_),
    .CLK(clknet_4_4_0_clk),
    .Q(\final_mant[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[5]$_DFFE_PP_  (.D(_0116_),
    .CLK(clknet_4_5_0_clk),
    .Q(\final_mant[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[6]$_DFFE_PP_  (.D(_0117_),
    .CLK(clknet_4_5_0_clk),
    .Q(\final_mant[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[7]$_DFFE_PP_  (.D(_0118_),
    .CLK(clknet_4_5_0_clk),
    .Q(\final_mant[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[8]$_DFFE_PP_  (.D(_0119_),
    .CLK(clknet_4_13_0_clk),
    .Q(\final_mant[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \final_mant[9]$_DFFE_PP_  (.D(_0120_),
    .CLK(clknet_4_6_0_clk),
    .Q(\final_mant[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \inexact$_DFF_PN0_  (.D(_0077_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \inexact_stage2$_DFF_PN0_  (.D(_0078_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(inexact_stage2));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \invalid_op$_DFF_PN0_  (.D(invalid_op_stage2),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \invalid_op_stage2$_DFFE_PN0P_  (.D(_0121_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(invalid_op_stage2));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \is_a_larger_stage1$_DFF_PN0_  (.D(a_exp_larger),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(is_a_larger_stage1));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[0]$_DFF_PN0_  (.D(net164),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[1]$_DFF_PN0_  (.D(net162),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\larger_exp_stage1[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[2]$_DFF_PN0_  (.D(net159),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\larger_exp_stage1[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[3]$_DFF_PN0_  (.D(net154),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\larger_exp_stage1[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[4]$_DFF_PN0_  (.D(net140),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[5]$_DFF_PN0_  (.D(net156),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[6]$_DFF_PN0_  (.D(net136),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \larger_exp_stage1[7]$_DFF_PN0_  (.D(net145),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \overflow$_DFF_PN0_  (.D(_0087_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[0]$_DFF_PN0_  (.D(\final_mant[0] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[10]$_DFF_PN0_  (.D(\final_mant[10] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[11]$_DFF_PN0_  (.D(\final_mant[11] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[12]$_DFF_PN0_  (.D(\final_mant[12] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[13]$_DFF_PN0_  (.D(\final_mant[13] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[14]$_DFF_PN0_  (.D(\final_mant[14] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net76));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[15]$_DFF_PN0_  (.D(\final_mant[15] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net77));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[16]$_DFF_PN0_  (.D(\final_mant[16] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net78));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[17]$_DFF_PN0_  (.D(\final_mant[17] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net79));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[18]$_DFF_PN0_  (.D(\final_mant[18] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net80));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[19]$_DFF_PN0_  (.D(\final_mant[19] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(net81));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[1]$_DFF_PN0_  (.D(\final_mant[1] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net82));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[20]$_DFF_PN0_  (.D(\final_mant[20] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net83));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[21]$_DFF_PN0_  (.D(\final_mant[21] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net84));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[22]$_DFF_PN0_  (.D(\final_mant[22] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net85));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[23]$_DFF_PN0_  (.D(\final_exp[0] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net86));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[24]$_DFF_PN0_  (.D(\final_exp[1] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net87));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[25]$_DFF_PN0_  (.D(\final_exp[2] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net88));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[26]$_DFF_PN0_  (.D(\final_exp[3] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net89));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[27]$_DFF_PN0_  (.D(\final_exp[4] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net90));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[28]$_DFF_PN0_  (.D(\final_exp[5] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(net91));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[29]$_DFF_PN0_  (.D(\final_exp[6] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(net92));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[2]$_DFF_PN0_  (.D(\final_mant[2] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net93));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[30]$_DFF_PN0_  (.D(\final_exp[7] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net94));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[31]$_DFF_PN0_  (.D(result_sign_stage2),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(net95));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[3]$_DFF_PN0_  (.D(\final_mant[3] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net96));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[4]$_DFF_PN0_  (.D(\final_mant[4] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net97));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[5]$_DFF_PN0_  (.D(\final_mant[5] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net98));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[6]$_DFF_PN0_  (.D(\final_mant[6] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net99));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[7]$_DFF_PN0_  (.D(\final_mant[7] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[8]$_DFF_PN0_  (.D(\final_mant[8] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result[9]$_DFF_PN0_  (.D(\final_mant[9] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[0]$_DFF_PN0_  (.D(\larger_exp_stage1[0] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \result_exp_stage2[1]$_DFF_PN0_  (.D(\larger_exp_stage1[1] ),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\result_exp_stage2[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[2]$_DFF_PN0_  (.D(\larger_exp_stage1[2] ),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\result_exp_stage2[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[3]$_DFF_PN0_  (.D(\larger_exp_stage1[3] ),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\result_exp_stage2[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[4]$_DFF_PN0_  (.D(\larger_exp_stage1[4] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[5]$_DFF_PN0_  (.D(\larger_exp_stage1[5] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[6]$_DFF_PN0_  (.D(\larger_exp_stage1[6] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_exp_stage2[7]$_DFF_PN0_  (.D(\larger_exp_stage1[7] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \result_sign_stage2$_DFF_PN0_  (.D(_0088_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(result_sign_stage2));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \underflow$_DFF_PN0_  (.D(_0089_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \valid_out$_DFF_PN0_  (.D(valid_stage2),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \valid_stage1$_DFF_PN0_  (.D(net67),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(valid_stage1));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \valid_stage2$_DFF_PN0_  (.D(valid_stage1),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(valid_stage2));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net66),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_359 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net125),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(net113),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input3 (.I(net119),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input4 (.I(a[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(a[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input6 (.I(net127),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(net108),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(net109),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input9 (.I(net118),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input10 (.I(net147),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input11 (.I(net130),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(net116),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input13 (.I(net120),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input14 (.I(net117),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input15 (.I(net112),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input16 (.I(a[23]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input17 (.I(net161),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input18 (.I(a[25]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(net153),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(net139),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input21 (.I(a[28]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(net135),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input23 (.I(net114),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input24 (.I(a[30]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input25 (.I(net106),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input26 (.I(net142),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input27 (.I(net115),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input28 (.I(net133),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input29 (.I(net111),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(a[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input31 (.I(net124),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(a[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(net128),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input34 (.I(net131),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input35 (.I(net157),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input36 (.I(net151),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input37 (.I(net149),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input38 (.I(net129),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input39 (.I(net160),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input40 (.I(net134),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input41 (.I(net148),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input42 (.I(net137),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input43 (.I(net121),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(net132),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input45 (.I(net146),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input46 (.I(net123),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input47 (.I(net152),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input48 (.I(net163),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input49 (.I(b[24]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input50 (.I(net158),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input51 (.I(b[26]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input52 (.I(b[27]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input53 (.I(net155),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input54 (.I(b[29]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input55 (.I(net143),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input56 (.I(net144),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input57 (.I(net105),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input58 (.I(net138),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input59 (.I(net126),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(b[5]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input61 (.I(net150),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input62 (.I(net141),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(net110),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input64 (.I(net122),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input65 (.I(net107),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input66 (.I(valid_in),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net68),
    .Z(inexact));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net69),
    .Z(invalid_op));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(overflow));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(result[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net72),
    .Z(result[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net73),
    .Z(result[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net74),
    .Z(result[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net75),
    .Z(result[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net76),
    .Z(result[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net77),
    .Z(result[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net78),
    .Z(result[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net79),
    .Z(result[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net80),
    .Z(result[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net81),
    .Z(result[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net82),
    .Z(result[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net83),
    .Z(result[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net84),
    .Z(result[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net85),
    .Z(result[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net86),
    .Z(result[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net87),
    .Z(result[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net88),
    .Z(result[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net89),
    .Z(result[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net90),
    .Z(result[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net91),
    .Z(result[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net92),
    .Z(result[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net93),
    .Z(result[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net94),
    .Z(result[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net95),
    .Z(result[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net96),
    .Z(result[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net97),
    .Z(result[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net98),
    .Z(result[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net99),
    .Z(result[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net100),
    .Z(result[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net101),
    .Z(result[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net102),
    .Z(result[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net103),
    .Z(underflow));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net104),
    .Z(valid_out));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload0 (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload1 (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload2 (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload3 (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload4 (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload5 (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload6 (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload7 (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload8 (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload9 (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload10 (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload11 (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload12 (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload13 (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload14 (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(b[31]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(a[31]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold4 (.I(rst_n),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold5 (.I(a[15]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold6 (.I(a[16]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold7 (.I(b[8]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold8 (.I(a[6]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold9 (.I(a[22]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold10 (.I(a[10]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold11 (.I(a[2]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold12 (.I(a[4]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold13 (.I(a[1]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold14 (.I(a[21]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold15 (.I(a[17]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold16 (.I(a[11]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold17 (.I(a[20]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold18 (.I(b[19]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold19 (.I(b[9]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold20 (.I(b[21]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold21 (.I(a[8]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold22 (.I(a[0]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold23 (.I(b[4]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold24 (.I(a[14]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold25 (.I(b[0]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold26 (.I(b[14]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold27 (.I(a[19]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold28 (.I(b[10]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold29 (.I(b[1]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold30 (.I(a[5]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold31 (.I(b[16]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold32 (.I(a[29]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold33 (.I(_0085_),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold34 (.I(b[18]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold35 (.I(b[3]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold36 (.I(a[27]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold37 (.I(_0083_),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold38 (.I(b[7]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold39 (.I(a[3]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold40 (.I(b[2]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold41 (.I(b[30]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold42 (.I(_0086_),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold43 (.I(b[20]),
    .Z(net146));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold44 (.I(a[18]),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold45 (.I(b[17]),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold46 (.I(b[13]),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold47 (.I(b[6]),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold48 (.I(b[12]),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold49 (.I(b[22]),
    .Z(net152));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold50 (.I(a[26]),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold51 (.I(_0082_),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold52 (.I(b[28]),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold53 (.I(_0084_),
    .Z(net156));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold54 (.I(b[11]),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold55 (.I(b[25]),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold56 (.I(_0081_),
    .Z(net159));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold57 (.I(b[15]),
    .Z(net160));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold58 (.I(a[24]),
    .Z(net161));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold59 (.I(_0080_),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold60 (.I(b[23]),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold61 (.I(_0079_),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_802 ();
endmodule
