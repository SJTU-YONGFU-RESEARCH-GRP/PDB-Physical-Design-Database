module fwft_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    data_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 output [4:0] data_count;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire output_valid;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net30;

 sky130_fd_sc_hd__inv_1 _168_ (.A(_151_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _169_ (.A(_156_),
    .B(_153_),
    .Y(_044_));
 sky130_fd_sc_hd__a21oi_1 _170_ (.A1(_156_),
    .A2(_152_),
    .B1(_155_),
    .Y(_045_));
 sky130_fd_sc_hd__o21ai_1 _171_ (.A1(_166_),
    .A2(_044_),
    .B1(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__xnor2_1 _172_ (.A(_043_),
    .B(_046_),
    .Y(net18));
 sky130_fd_sc_hd__xor2_2 _173_ (.A(_156_),
    .B(_148_),
    .X(net17));
 sky130_fd_sc_hd__a21o_1 _174_ (.A1(_156_),
    .A2(_148_),
    .B1(_155_),
    .X(_047_));
 sky130_fd_sc_hd__a21oi_2 _175_ (.A1(_151_),
    .A2(_047_),
    .B1(_150_),
    .Y(_048_));
 sky130_fd_sc_hd__xnor2_2 _176_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Y(_049_));
 sky130_fd_sc_hd__xor2_4 _177_ (.A(_048_),
    .B(_049_),
    .X(_050_));
 sky130_fd_sc_hd__clkinv_4 _178_ (.A(_050_),
    .Y(net19));
 sky130_fd_sc_hd__inv_1 _179_ (.A(_167_),
    .Y(net15));
 sky130_fd_sc_hd__nor4_1 _180_ (.A(_151_),
    .B(net15),
    .C(net16),
    .D(net17),
    .Y(_051_));
 sky130_fd_sc_hd__nor4_1 _181_ (.A(_043_),
    .B(net15),
    .C(net16),
    .D(net17),
    .Y(_052_));
 sky130_fd_sc_hd__mux2_1 _182_ (.A0(_051_),
    .A1(_052_),
    .S(_046_),
    .X(_053_));
 sky130_fd_sc_hd__buf_6 _183_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__and2_0 _184_ (.A(_050_),
    .B(_054_),
    .X(_055_));
 sky130_fd_sc_hd__nor3b_4 _185_ (.A(output_valid),
    .B(_055_),
    .C_N(net3),
    .Y(_000_));
 sky130_fd_sc_hd__and2_0 _186_ (.A(net19),
    .B(_054_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 _187_ (.A(\rd_ptr[0] ),
    .X(_056_));
 sky130_fd_sc_hd__buf_4 _188_ (.A(_056_),
    .X(_057_));
 sky130_fd_sc_hd__inv_1 _189_ (.A(_057_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_1 _190_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .Y(_058_));
 sky130_fd_sc_hd__a21boi_2 _191_ (.A1(net19),
    .A2(_053_),
    .B1_N(net12),
    .Y(_059_));
 sky130_fd_sc_hd__and3_4 _192_ (.A(_158_),
    .B(_058_),
    .C(_059_),
    .X(_001_));
 sky130_fd_sc_hd__and3_4 _193_ (.A(_161_),
    .B(_058_),
    .C(_059_),
    .X(_008_));
 sky130_fd_sc_hd__and3_4 _194_ (.A(_159_),
    .B(_058_),
    .C(_059_),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _195_ (.A(net12),
    .B(_163_),
    .Y(_060_));
 sky130_fd_sc_hd__a21oi_2 _196_ (.A1(net19),
    .A2(_054_),
    .B1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__and2_4 _197_ (.A(_058_),
    .B(_061_),
    .X(_010_));
 sky130_fd_sc_hd__buf_6 _198_ (.A(_059_),
    .X(_062_));
 sky130_fd_sc_hd__nor2b_1 _199_ (.A(\wr_ptr[3] ),
    .B_N(\wr_ptr[2] ),
    .Y(_063_));
 sky130_fd_sc_hd__and3_4 _200_ (.A(_158_),
    .B(_062_),
    .C(_063_),
    .X(_011_));
 sky130_fd_sc_hd__and3_4 _201_ (.A(_161_),
    .B(_062_),
    .C(_063_),
    .X(_012_));
 sky130_fd_sc_hd__and3_4 _202_ (.A(_159_),
    .B(_062_),
    .C(_063_),
    .X(_013_));
 sky130_fd_sc_hd__and2_4 _203_ (.A(_061_),
    .B(_063_),
    .X(_014_));
 sky130_fd_sc_hd__nor2b_2 _204_ (.A(\wr_ptr[2] ),
    .B_N(\wr_ptr[3] ),
    .Y(_064_));
 sky130_fd_sc_hd__and3_4 _205_ (.A(_158_),
    .B(_062_),
    .C(_064_),
    .X(_015_));
 sky130_fd_sc_hd__and3_4 _206_ (.A(_161_),
    .B(_062_),
    .C(_064_),
    .X(_016_));
 sky130_fd_sc_hd__and3_4 _207_ (.A(_159_),
    .B(_062_),
    .C(_064_),
    .X(_002_));
 sky130_fd_sc_hd__and2_4 _208_ (.A(_061_),
    .B(_064_),
    .X(_003_));
 sky130_fd_sc_hd__and2_1 _209_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .X(_065_));
 sky130_fd_sc_hd__and3_4 _210_ (.A(_158_),
    .B(_062_),
    .C(_065_),
    .X(_004_));
 sky130_fd_sc_hd__and3_4 _211_ (.A(_161_),
    .B(_062_),
    .C(_065_),
    .X(_005_));
 sky130_fd_sc_hd__and3_4 _212_ (.A(_159_),
    .B(_062_),
    .C(_065_),
    .X(_006_));
 sky130_fd_sc_hd__nand3_1 _213_ (.A(net12),
    .B(_163_),
    .C(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__a21oi_4 _214_ (.A1(net19),
    .A2(_054_),
    .B1(_066_),
    .Y(_007_));
 sky130_fd_sc_hd__buf_4 _215_ (.A(\rd_ptr[2] ),
    .X(_067_));
 sky130_fd_sc_hd__clkbuf_4 _216_ (.A(_067_),
    .X(_068_));
 sky130_fd_sc_hd__xor2_1 _217_ (.A(_068_),
    .B(_165_),
    .X(_019_));
 sky130_fd_sc_hd__nand3_1 _218_ (.A(_057_),
    .B(\rd_ptr[1] ),
    .C(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__xnor2_1 _219_ (.A(\rd_ptr[3] ),
    .B(_069_),
    .Y(_020_));
 sky130_fd_sc_hd__nand3_1 _220_ (.A(_068_),
    .B(\rd_ptr[3] ),
    .C(_165_),
    .Y(_070_));
 sky130_fd_sc_hd__xnor2_1 _221_ (.A(\rd_ptr[4] ),
    .B(_070_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _222_ (.A(\rd_ptr[3] ),
    .Y(_149_));
 sky130_fd_sc_hd__clkinv_4 _223_ (.A(\rd_ptr[1] ),
    .Y(_146_));
 sky130_fd_sc_hd__inv_1 _224_ (.A(_068_),
    .Y(_154_));
 sky130_fd_sc_hd__inv_1 _225_ (.A(\wr_ptr[0] ),
    .Y(_022_));
 sky130_fd_sc_hd__inv_1 _226_ (.A(_166_),
    .Y(_147_));
 sky130_fd_sc_hd__inv_1 _227_ (.A(\wr_ptr[1] ),
    .Y(_157_));
 sky130_fd_sc_hd__buf_6 _228_ (.A(_056_),
    .X(_071_));
 sky130_fd_sc_hd__buf_4 _229_ (.A(\rd_ptr[2] ),
    .X(_072_));
 sky130_fd_sc_hd__mux4_1 _230_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[4][0] ),
    .A3(\mem[5][0] ),
    .S0(_071_),
    .S1(_072_),
    .X(_073_));
 sky130_fd_sc_hd__nor2_4 _231_ (.A(\rd_ptr[1] ),
    .B(\rd_ptr[3] ),
    .Y(_074_));
 sky130_fd_sc_hd__nor2_4 _232_ (.A(\rd_ptr[1] ),
    .B(_149_),
    .Y(_075_));
 sky130_fd_sc_hd__mux4_1 _233_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[12][0] ),
    .A3(\mem[13][0] ),
    .S0(_071_),
    .S1(_072_),
    .X(_076_));
 sky130_fd_sc_hd__a22oi_1 _234_ (.A1(_073_),
    .A2(_074_),
    .B1(_075_),
    .B2(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__buf_4 _235_ (.A(_056_),
    .X(_078_));
 sky130_fd_sc_hd__mux4_1 _236_ (.A0(\mem[2][0] ),
    .A1(\mem[3][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(_078_),
    .S1(_072_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_8 _237_ (.A(_146_),
    .B(\rd_ptr[3] ),
    .Y(_080_));
 sky130_fd_sc_hd__nor2_8 _238_ (.A(_146_),
    .B(_149_),
    .Y(_081_));
 sky130_fd_sc_hd__mux4_1 _239_ (.A0(\mem[10][0] ),
    .A1(\mem[11][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(_071_),
    .S1(_072_),
    .X(_082_));
 sky130_fd_sc_hd__a22oi_1 _240_ (.A1(_079_),
    .A2(_080_),
    .B1(_081_),
    .B2(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__nand2_1 _241_ (.A(_077_),
    .B(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__inv_1 _242_ (.A(output_valid),
    .Y(net20));
 sky130_fd_sc_hd__o2bb2ai_4 _243_ (.A1_N(_050_),
    .A2_N(_054_),
    .B1(net2),
    .B2(net20),
    .Y(_085_));
 sky130_fd_sc_hd__mux2_1 _244_ (.A0(_084_),
    .A1(net22),
    .S(_085_),
    .X(_024_));
 sky130_fd_sc_hd__mux4_1 _245_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[12][1] ),
    .A3(\mem[13][1] ),
    .S0(_078_),
    .S1(_072_),
    .X(_086_));
 sky130_fd_sc_hd__mux4_1 _246_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[4][1] ),
    .A3(\mem[5][1] ),
    .S0(_057_),
    .S1(_068_),
    .X(_087_));
 sky130_fd_sc_hd__a22oi_1 _247_ (.A1(_075_),
    .A2(_086_),
    .B1(_087_),
    .B2(_074_),
    .Y(_088_));
 sky130_fd_sc_hd__mux4_1 _248_ (.A0(\mem[10][1] ),
    .A1(\mem[11][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(_078_),
    .S1(_067_),
    .X(_089_));
 sky130_fd_sc_hd__buf_4 _249_ (.A(_067_),
    .X(_090_));
 sky130_fd_sc_hd__mux4_1 _250_ (.A0(\mem[2][1] ),
    .A1(\mem[3][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(_071_),
    .S1(_090_),
    .X(_091_));
 sky130_fd_sc_hd__a22oi_2 _251_ (.A1(_081_),
    .A2(_089_),
    .B1(_091_),
    .B2(_080_),
    .Y(_092_));
 sky130_fd_sc_hd__nand2_1 _252_ (.A(_088_),
    .B(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__mux2_1 _253_ (.A0(_093_),
    .A1(net23),
    .S(_085_),
    .X(_025_));
 sky130_fd_sc_hd__mux4_1 _254_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[12][2] ),
    .A3(\mem[13][2] ),
    .S0(_078_),
    .S1(_072_),
    .X(_094_));
 sky130_fd_sc_hd__mux4_1 _255_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[4][2] ),
    .A3(\mem[5][2] ),
    .S0(_057_),
    .S1(_068_),
    .X(_095_));
 sky130_fd_sc_hd__a22oi_1 _256_ (.A1(_075_),
    .A2(_094_),
    .B1(_095_),
    .B2(_074_),
    .Y(_096_));
 sky130_fd_sc_hd__mux4_1 _257_ (.A0(\mem[10][2] ),
    .A1(\mem[11][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(_078_),
    .S1(_067_),
    .X(_097_));
 sky130_fd_sc_hd__mux4_1 _258_ (.A0(\mem[2][2] ),
    .A1(\mem[3][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(_071_),
    .S1(_090_),
    .X(_098_));
 sky130_fd_sc_hd__a22oi_2 _259_ (.A1(_081_),
    .A2(_097_),
    .B1(_098_),
    .B2(_080_),
    .Y(_099_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(_096_),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(_100_),
    .A1(net24),
    .S(_085_),
    .X(_026_));
 sky130_fd_sc_hd__mux4_1 _262_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[12][3] ),
    .A3(\mem[13][3] ),
    .S0(_078_),
    .S1(_072_),
    .X(_101_));
 sky130_fd_sc_hd__mux4_1 _263_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[4][3] ),
    .A3(\mem[5][3] ),
    .S0(_057_),
    .S1(_068_),
    .X(_102_));
 sky130_fd_sc_hd__a22oi_1 _264_ (.A1(_075_),
    .A2(_101_),
    .B1(_102_),
    .B2(_074_),
    .Y(_103_));
 sky130_fd_sc_hd__mux4_1 _265_ (.A0(\mem[10][3] ),
    .A1(\mem[11][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(_056_),
    .S1(_067_),
    .X(_104_));
 sky130_fd_sc_hd__mux4_4 _266_ (.A0(\mem[2][3] ),
    .A1(\mem[3][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(_071_),
    .S1(_090_),
    .X(_105_));
 sky130_fd_sc_hd__a22oi_4 _267_ (.A1(_081_),
    .A2(_104_),
    .B1(_105_),
    .B2(_080_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_1 _268_ (.A(_103_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(_107_),
    .A1(net25),
    .S(_085_),
    .X(_027_));
 sky130_fd_sc_hd__mux4_1 _270_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[12][4] ),
    .A3(\mem[13][4] ),
    .S0(_078_),
    .S1(_072_),
    .X(_108_));
 sky130_fd_sc_hd__mux4_1 _271_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[4][4] ),
    .A3(\mem[5][4] ),
    .S0(_057_),
    .S1(_068_),
    .X(_109_));
 sky130_fd_sc_hd__a22oi_1 _272_ (.A1(_075_),
    .A2(_108_),
    .B1(_109_),
    .B2(_074_),
    .Y(_110_));
 sky130_fd_sc_hd__mux4_1 _273_ (.A0(\mem[10][4] ),
    .A1(\mem[11][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(_056_),
    .S1(_067_),
    .X(_111_));
 sky130_fd_sc_hd__mux4_1 _274_ (.A0(\mem[2][4] ),
    .A1(\mem[3][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(_071_),
    .S1(_090_),
    .X(_112_));
 sky130_fd_sc_hd__a22oi_2 _275_ (.A1(_081_),
    .A2(_111_),
    .B1(_112_),
    .B2(_080_),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _276_ (.A(_110_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(_114_),
    .A1(net26),
    .S(_085_),
    .X(_028_));
 sky130_fd_sc_hd__mux4_1 _278_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[12][5] ),
    .A3(\mem[13][5] ),
    .S0(_078_),
    .S1(_072_),
    .X(_115_));
 sky130_fd_sc_hd__mux4_1 _279_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[4][5] ),
    .A3(\mem[5][5] ),
    .S0(_057_),
    .S1(_090_),
    .X(_116_));
 sky130_fd_sc_hd__a22oi_1 _280_ (.A1(_075_),
    .A2(_115_),
    .B1(_116_),
    .B2(_074_),
    .Y(_117_));
 sky130_fd_sc_hd__mux4_1 _281_ (.A0(\mem[10][5] ),
    .A1(\mem[11][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(_056_),
    .S1(_067_),
    .X(_118_));
 sky130_fd_sc_hd__mux4_1 _282_ (.A0(\mem[2][5] ),
    .A1(\mem[3][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(_071_),
    .S1(_090_),
    .X(_119_));
 sky130_fd_sc_hd__a22oi_2 _283_ (.A1(_081_),
    .A2(_118_),
    .B1(_119_),
    .B2(_080_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _284_ (.A(_117_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(_121_),
    .A1(net27),
    .S(_085_),
    .X(_029_));
 sky130_fd_sc_hd__mux4_1 _286_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[12][6] ),
    .A3(\mem[13][6] ),
    .S0(_078_),
    .S1(_072_),
    .X(_122_));
 sky130_fd_sc_hd__mux4_1 _287_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[4][6] ),
    .A3(\mem[5][6] ),
    .S0(_057_),
    .S1(_090_),
    .X(_123_));
 sky130_fd_sc_hd__a22oi_1 _288_ (.A1(_075_),
    .A2(_122_),
    .B1(_123_),
    .B2(_074_),
    .Y(_124_));
 sky130_fd_sc_hd__mux4_1 _289_ (.A0(\mem[10][6] ),
    .A1(\mem[11][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(_056_),
    .S1(_067_),
    .X(_125_));
 sky130_fd_sc_hd__mux4_1 _290_ (.A0(\mem[2][6] ),
    .A1(\mem[3][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(_071_),
    .S1(_090_),
    .X(_126_));
 sky130_fd_sc_hd__a22oi_2 _291_ (.A1(_081_),
    .A2(_125_),
    .B1(_126_),
    .B2(_080_),
    .Y(_127_));
 sky130_fd_sc_hd__nand2_1 _292_ (.A(_124_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(_128_),
    .A1(net28),
    .S(_085_),
    .X(_030_));
 sky130_fd_sc_hd__mux4_1 _294_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[12][7] ),
    .A3(\mem[13][7] ),
    .S0(_078_),
    .S1(_067_),
    .X(_129_));
 sky130_fd_sc_hd__mux4_1 _295_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[4][7] ),
    .A3(\mem[5][7] ),
    .S0(_057_),
    .S1(_090_),
    .X(_130_));
 sky130_fd_sc_hd__a22oi_1 _296_ (.A1(_075_),
    .A2(_129_),
    .B1(_130_),
    .B2(_074_),
    .Y(_131_));
 sky130_fd_sc_hd__mux4_1 _297_ (.A0(\mem[10][7] ),
    .A1(\mem[11][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(_056_),
    .S1(_067_),
    .X(_132_));
 sky130_fd_sc_hd__mux4_1 _298_ (.A0(\mem[2][7] ),
    .A1(\mem[3][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(_071_),
    .S1(_090_),
    .X(_133_));
 sky130_fd_sc_hd__a22oi_2 _299_ (.A1(_081_),
    .A2(_132_),
    .B1(_133_),
    .B2(_080_),
    .Y(_134_));
 sky130_fd_sc_hd__nand2_1 _300_ (.A(_131_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__mux2_1 _301_ (.A0(_135_),
    .A1(net29),
    .S(_085_),
    .X(_031_));
 sky130_fd_sc_hd__o21ai_0 _302_ (.A1(net2),
    .A2(net20),
    .B1(_055_),
    .Y(_032_));
 sky130_fd_sc_hd__a21boi_1 _303_ (.A1(_050_),
    .A2(_054_),
    .B1_N(net2),
    .Y(_136_));
 sky130_fd_sc_hd__xnor2_1 _304_ (.A(_017_),
    .B(_136_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(\rd_ptr[1] ),
    .A1(_018_),
    .S(_136_),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _306_ (.A(net2),
    .B(_165_),
    .Y(_137_));
 sky130_fd_sc_hd__a21oi_1 _307_ (.A1(_050_),
    .A2(_054_),
    .B1(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__xnor2_1 _308_ (.A(_154_),
    .B(_138_),
    .Y(_035_));
 sky130_fd_sc_hd__nand4_1 _309_ (.A(net2),
    .B(_057_),
    .C(\rd_ptr[1] ),
    .D(_068_),
    .Y(_139_));
 sky130_fd_sc_hd__a21oi_1 _310_ (.A1(_050_),
    .A2(_054_),
    .B1(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__xnor2_1 _311_ (.A(_149_),
    .B(_140_),
    .Y(_036_));
 sky130_fd_sc_hd__nand4_1 _312_ (.A(net2),
    .B(_068_),
    .C(\rd_ptr[3] ),
    .D(_165_),
    .Y(_141_));
 sky130_fd_sc_hd__a21oi_1 _313_ (.A1(_050_),
    .A2(_054_),
    .B1(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__xor2_1 _314_ (.A(\rd_ptr[4] ),
    .B(_142_),
    .X(_037_));
 sky130_fd_sc_hd__xnor2_1 _315_ (.A(_022_),
    .B(_062_),
    .Y(_038_));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(\wr_ptr[1] ),
    .A1(_023_),
    .S(_059_),
    .X(_039_));
 sky130_fd_sc_hd__xor2_1 _317_ (.A(\wr_ptr[2] ),
    .B(_061_),
    .X(_040_));
 sky130_fd_sc_hd__nand4_1 _318_ (.A(net12),
    .B(\wr_ptr[2] ),
    .C(\wr_ptr[1] ),
    .D(\wr_ptr[0] ),
    .Y(_143_));
 sky130_fd_sc_hd__a21oi_1 _319_ (.A1(net19),
    .A2(_054_),
    .B1(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__xor2_1 _320_ (.A(\wr_ptr[3] ),
    .B(_144_),
    .X(_041_));
 sky130_fd_sc_hd__xor2_1 _321_ (.A(\wr_ptr[4] ),
    .B(_007_),
    .X(_042_));
 sky130_fd_sc_hd__xor2_1 _322_ (.A(_167_),
    .B(net16),
    .X(_145_));
 sky130_fd_sc_hd__nor4_1 _323_ (.A(net18),
    .B(net17),
    .C(net19),
    .D(_145_),
    .Y(net13));
 sky130_fd_sc_hd__a31o_1 _324_ (.A1(net16),
    .A2(net18),
    .A3(net17),
    .B1(net19),
    .X(net14));
 sky130_fd_sc_hd__fa_2 _325_ (.A(_146_),
    .B(\wr_ptr[1] ),
    .CIN(_147_),
    .COUT(_148_),
    .SUM(net16));
 sky130_fd_sc_hd__ha_1 _326_ (.A(_149_),
    .B(\wr_ptr[3] ),
    .COUT(_150_),
    .SUM(_151_));
 sky130_fd_sc_hd__ha_1 _327_ (.A(_146_),
    .B(\wr_ptr[1] ),
    .COUT(_152_),
    .SUM(_153_));
 sky130_fd_sc_hd__ha_1 _328_ (.A(_154_),
    .B(\wr_ptr[2] ),
    .COUT(_155_),
    .SUM(_156_));
 sky130_fd_sc_hd__ha_1 _329_ (.A(_022_),
    .B(_157_),
    .COUT(_158_),
    .SUM(_023_));
 sky130_fd_sc_hd__ha_1 _330_ (.A(_022_),
    .B(\wr_ptr[1] ),
    .COUT(_159_),
    .SUM(_160_));
 sky130_fd_sc_hd__ha_1 _331_ (.A(\wr_ptr[0] ),
    .B(_157_),
    .COUT(_161_),
    .SUM(_162_));
 sky130_fd_sc_hd__ha_1 _332_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_163_),
    .SUM(_164_));
 sky130_fd_sc_hd__ha_1 _333_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_165_),
    .SUM(_018_));
 sky130_fd_sc_hd__ha_1 _334_ (.A(\rd_ptr[0] ),
    .B(_022_),
    .COUT(_166_),
    .SUM(_167_));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\mem[0][0] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\mem[0][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\mem[0][2] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\mem[0][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\mem[0][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\mem[0][5] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net10),
    .DE(_001_),
    .Q(\mem[0][6] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net11),
    .DE(_001_),
    .Q(\mem[0][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\mem[10][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\mem[10][1] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\mem[10][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\mem[10][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\mem[10][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\mem[10][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net10),
    .DE(_002_),
    .Q(\mem[10][6] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net11),
    .DE(_002_),
    .Q(\mem[10][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\mem[11][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\mem[11][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\mem[11][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\mem[11][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\mem[11][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\mem[11][5] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net10),
    .DE(_003_),
    .Q(\mem[11][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net11),
    .DE(_003_),
    .Q(\mem[11][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\mem[12][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\mem[12][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\mem[12][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\mem[12][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\mem[12][4] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\mem[12][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net10),
    .DE(_004_),
    .Q(\mem[12][6] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net11),
    .DE(_004_),
    .Q(\mem[12][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\mem[13][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\mem[13][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\mem[13][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\mem[13][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\mem[13][4] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\mem[13][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net10),
    .DE(_005_),
    .Q(\mem[13][6] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net11),
    .DE(_005_),
    .Q(\mem[13][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\mem[14][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\mem[14][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\mem[14][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\mem[14][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\mem[14][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\mem[14][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net10),
    .DE(_006_),
    .Q(\mem[14][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net11),
    .DE(_006_),
    .Q(\mem[14][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\mem[15][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\mem[15][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\mem[15][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\mem[15][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\mem[15][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\mem[15][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net10),
    .DE(_007_),
    .Q(\mem[15][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net11),
    .DE(_007_),
    .Q(\mem[15][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\mem[1][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\mem[1][1] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\mem[1][2] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\mem[1][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\mem[1][4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\mem[1][5] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net10),
    .DE(_008_),
    .Q(\mem[1][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net11),
    .DE(_008_),
    .Q(\mem[1][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\mem[2][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\mem[2][1] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\mem[2][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\mem[2][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[2][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[2][5] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\mem[2][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net11),
    .DE(_009_),
    .Q(\mem[2][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\mem[3][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\mem[3][1] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\mem[3][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\mem[3][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[3][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[3][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\mem[3][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net11),
    .DE(_010_),
    .Q(\mem[3][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\mem[4][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[4][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[4][2] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[4][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[4][4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[4][5] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[4][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net11),
    .DE(_011_),
    .Q(\mem[4][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\mem[5][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[5][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[5][2] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[5][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[5][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[5][5] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[5][6] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net11),
    .DE(_012_),
    .Q(\mem[5][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\mem[6][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[6][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[6][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[6][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[6][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[6][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[6][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net11),
    .DE(_013_),
    .Q(\mem[6][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\mem[7][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[7][1] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[7][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[7][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[7][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[7][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[7][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net11),
    .DE(_014_),
    .Q(\mem[7][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\mem[8][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[8][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[8][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[8][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[8][4] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[8][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[8][6] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net11),
    .DE(_015_),
    .Q(\mem[8][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net4),
    .DE(_016_),
    .Q(\mem[9][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net5),
    .DE(_016_),
    .Q(\mem[9][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net6),
    .DE(_016_),
    .Q(\mem[9][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net7),
    .DE(_016_),
    .Q(\mem[9][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net8),
    .DE(_016_),
    .Q(\mem[9][4] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net9),
    .DE(_016_),
    .Q(\mem[9][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net10),
    .DE(_016_),
    .Q(\mem[9][6] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net11),
    .DE(_016_),
    .Q(\mem[9][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[0]$_DFFE_PN0P_  (.D(_024_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[1]$_DFFE_PN0P_  (.D(_025_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[2]$_DFFE_PN0P_  (.D(_026_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[3]$_DFFE_PN0P_  (.D(_027_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[4]$_DFFE_PN0P_  (.D(_028_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[5]$_DFFE_PN0P_  (.D(_029_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[6]$_DFFE_PN0P_  (.D(_030_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_reg[7]$_DFFE_PN0P_  (.D(_031_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \output_valid$_DFFE_PN0P_  (.D(_032_),
    .Q(output_valid),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0P_  (.D(_033_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \rd_ptr[0]$_DFFE_PP_  (.D(_017_),
    .DE(_000_),
    .Q(\rd_ptr[0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr[1]$_DFFE_PN0P_  (.D(_034_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \rd_ptr[1]$_DFFE_PP_  (.D(_018_),
    .DE(_000_),
    .Q(\rd_ptr[1] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_035_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \rd_ptr[2]$_DFFE_PP_  (.D(_019_),
    .DE(_000_),
    .Q(\rd_ptr[2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr[3]$_DFFE_PN0P_  (.D(_036_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \rd_ptr[3]$_DFFE_PP_  (.D(_020_),
    .DE(_000_),
    .Q(\rd_ptr[3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr[4]$_DFFE_PN0P_  (.D(_037_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \rd_ptr[4]$_DFFE_PP_  (.D(_021_),
    .DE(_000_),
    .Q(\rd_ptr[4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_038_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_039_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[2]$_DFFE_PN0P_  (.D(_040_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[3]$_DFFE_PN0P_  (.D(_041_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_042_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__buf_8 hold1 (.A(net3),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_139 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net30),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(wr_data[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input4 (.A(wr_data[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(wr_data[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input6 (.A(wr_data[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input8 (.A(wr_data[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input9 (.A(wr_data[6]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input10 (.A(wr_data[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wr_en),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(data_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(data_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(data_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(data_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(data_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload10 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload11 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload13 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net30));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_229 ();
endmodule
