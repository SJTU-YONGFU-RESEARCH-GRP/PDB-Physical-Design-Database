module radix4_booth_multiplier (clk,
    done,
    rst_n,
    start,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst_n;
 input start;
 input [7:0] multiplicand;
 input [7:0] multiplier;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire \a_reg[0] ;
 wire \a_reg[1] ;
 wire \a_reg[2] ;
 wire \a_reg[3] ;
 wire \a_reg[4] ;
 wire \a_reg[5] ;
 wire \a_reg[6] ;
 wire \a_reg[7] ;
 wire \b_reg[0] ;
 wire \b_reg[1] ;
 wire \b_reg[2] ;
 wire \b_reg[3] ;
 wire \b_reg[4] ;
 wire \b_reg[5] ;
 wire \b_reg[6] ;
 wire \b_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net36;
 wire net37;
 wire net38;

 INV_X1 _494_ (.A(\state[1] ),
    .ZN(_036_));
 BUF_X2 _495_ (.A(net17),
    .Z(_037_));
 BUF_X2 _496_ (.A(_037_),
    .Z(_038_));
 INV_X1 _497_ (.A(net18),
    .ZN(_039_));
 NAND2_X1 _498_ (.A1(_039_),
    .A2(\state[0] ),
    .ZN(_040_));
 NAND3_X1 _499_ (.A1(_036_),
    .A2(_038_),
    .A3(_040_),
    .ZN(_002_));
 BUF_X2 _500_ (.A(\b_reg[0] ),
    .Z(_041_));
 BUF_X2 _501_ (.A(\a_reg[6] ),
    .Z(_042_));
 NAND2_X1 _502_ (.A1(_041_),
    .A2(_042_),
    .ZN(_211_));
 BUF_X2 _503_ (.A(\b_reg[1] ),
    .Z(_043_));
 BUF_X2 _504_ (.A(\a_reg[5] ),
    .Z(_044_));
 NAND2_X1 _505_ (.A1(_043_),
    .A2(_044_),
    .ZN(_210_));
 BUF_X2 _506_ (.A(\b_reg[2] ),
    .Z(_045_));
 BUF_X2 _507_ (.A(\a_reg[4] ),
    .Z(_046_));
 NAND2_X1 _508_ (.A1(_045_),
    .A2(_046_),
    .ZN(_209_));
 AND2_X1 _509_ (.A1(_043_),
    .A2(_046_),
    .ZN(_223_));
 BUF_X2 _510_ (.A(\a_reg[3] ),
    .Z(_047_));
 AND2_X1 _511_ (.A1(_045_),
    .A2(_047_),
    .ZN(_222_));
 BUF_X2 _512_ (.A(\b_reg[3] ),
    .Z(_048_));
 AND2_X1 _513_ (.A1(_047_),
    .A2(_048_),
    .ZN(_216_));
 BUF_X2 _514_ (.A(\b_reg[4] ),
    .Z(_049_));
 BUF_X2 _515_ (.A(\a_reg[2] ),
    .Z(_050_));
 AND2_X1 _516_ (.A1(_049_),
    .A2(_050_),
    .ZN(_215_));
 BUF_X2 _517_ (.A(\b_reg[5] ),
    .Z(_051_));
 BUF_X2 _518_ (.A(\a_reg[1] ),
    .Z(_052_));
 AND2_X1 _519_ (.A1(_051_),
    .A2(_052_),
    .ZN(_214_));
 AND2_X1 _520_ (.A1(_043_),
    .A2(_047_),
    .ZN(_241_));
 AND2_X1 _521_ (.A1(_045_),
    .A2(_050_),
    .ZN(_240_));
 BUF_X2 _522_ (.A(\a_reg[0] ),
    .Z(_053_));
 BUF_X2 _523_ (.A(\b_reg[6] ),
    .Z(_054_));
 AND2_X1 _524_ (.A1(_053_),
    .A2(_054_),
    .ZN(_406_));
 NAND2_X1 _525_ (.A1(_041_),
    .A2(_047_),
    .ZN(_256_));
 AND2_X1 _526_ (.A1(_048_),
    .A2(_052_),
    .ZN(_409_));
 AND2_X1 _527_ (.A1(_049_),
    .A2(_053_),
    .ZN(_408_));
 NAND2_X1 _528_ (.A1(_041_),
    .A2(_050_),
    .ZN(_265_));
 AND2_X1 _529_ (.A1(_048_),
    .A2(_053_),
    .ZN(_258_));
 AND2_X1 _530_ (.A1(_041_),
    .A2(_052_),
    .ZN(_485_));
 AND2_X1 _531_ (.A1(_043_),
    .A2(_053_),
    .ZN(_484_));
 NAND2_X1 _532_ (.A1(_042_),
    .A2(_043_),
    .ZN(_274_));
 NAND2_X1 _533_ (.A1(_044_),
    .A2(_045_),
    .ZN(_280_));
 NAND2_X1 _534_ (.A1(_046_),
    .A2(_048_),
    .ZN(_279_));
 NAND2_X1 _535_ (.A1(_047_),
    .A2(_049_),
    .ZN(_278_));
 INV_X2 _536_ (.A(\b_reg[7] ),
    .ZN(_055_));
 OR2_X1 _537_ (.A1(_053_),
    .A2(_055_),
    .ZN(_285_));
 AND2_X1 _538_ (.A1(_042_),
    .A2(_045_),
    .ZN(_427_));
 NAND2_X1 _539_ (.A1(_044_),
    .A2(_048_),
    .ZN(_298_));
 NAND2_X1 _540_ (.A1(_046_),
    .A2(_049_),
    .ZN(_297_));
 NAND2_X1 _541_ (.A1(_047_),
    .A2(_051_),
    .ZN(_299_));
 AND2_X1 _542_ (.A1(_050_),
    .A2(_054_),
    .ZN(_432_));
 NOR2_X1 _543_ (.A1(_052_),
    .A2(_055_),
    .ZN(_431_));
 INV_X1 _544_ (.A(_313_),
    .ZN(_310_));
 BUF_X2 _545_ (.A(\a_reg[7] ),
    .Z(_056_));
 AND2_X1 _546_ (.A1(_045_),
    .A2(_056_),
    .ZN(_437_));
 AND3_X1 _547_ (.A1(_041_),
    .A2(_043_),
    .A3(_056_),
    .ZN(_057_));
 NOR2_X1 _548_ (.A1(_429_),
    .A2(_057_),
    .ZN(_319_));
 NAND2_X1 _549_ (.A1(_042_),
    .A2(_048_),
    .ZN(_316_));
 NAND2_X1 _550_ (.A1(_044_),
    .A2(_049_),
    .ZN(_315_));
 NAND2_X1 _551_ (.A1(_046_),
    .A2(_051_),
    .ZN(_314_));
 AND2_X1 _552_ (.A1(_047_),
    .A2(_054_),
    .ZN(_441_));
 NOR2_X1 _553_ (.A1(_050_),
    .A2(_055_),
    .ZN(_440_));
 NOR2_X2 _554_ (.A1(_438_),
    .A2(_057_),
    .ZN(_338_));
 AND2_X2 _555_ (.A1(_048_),
    .A2(_056_),
    .ZN(_333_));
 AND2_X1 _556_ (.A1(_042_),
    .A2(_049_),
    .ZN(_334_));
 AND2_X1 _557_ (.A1(_044_),
    .A2(_051_),
    .ZN(_335_));
 AND2_X1 _558_ (.A1(_046_),
    .A2(_054_),
    .ZN(_447_));
 NOR2_X1 _559_ (.A1(_047_),
    .A2(_055_),
    .ZN(_446_));
 INV_X1 _560_ (.A(_422_),
    .ZN(_268_));
 AND2_X1 _561_ (.A1(_049_),
    .A2(_056_),
    .ZN(_354_));
 AND2_X1 _562_ (.A1(_042_),
    .A2(_051_),
    .ZN(_353_));
 AND2_X1 _563_ (.A1(_044_),
    .A2(_054_),
    .ZN(_453_));
 NOR2_X1 _564_ (.A1(_046_),
    .A2(_055_),
    .ZN(_452_));
 AND2_X1 _565_ (.A1(_051_),
    .A2(_056_),
    .ZN(_370_));
 AND2_X1 _566_ (.A1(_042_),
    .A2(_054_),
    .ZN(_459_));
 NOR2_X1 _567_ (.A1(_044_),
    .A2(_055_),
    .ZN(_460_));
 AND2_X1 _568_ (.A1(_054_),
    .A2(_056_),
    .ZN(_468_));
 NOR2_X1 _569_ (.A1(_042_),
    .A2(_055_),
    .ZN(_469_));
 CLKBUF_X2 _570_ (.A(\state[2] ),
    .Z(_058_));
 NAND2_X1 _571_ (.A1(net17),
    .A2(_058_),
    .ZN(_059_));
 INV_X1 _572_ (.A(_059_),
    .ZN(_000_));
 INV_X1 _573_ (.A(net17),
    .ZN(_060_));
 CLKBUF_X3 _574_ (.A(_060_),
    .Z(_061_));
 NAND2_X4 _575_ (.A1(net18),
    .A2(\state[0] ),
    .ZN(_062_));
 BUF_X4 _576_ (.A(_062_),
    .Z(_063_));
 NOR2_X1 _577_ (.A1(_061_),
    .A2(_063_),
    .ZN(_001_));
 NAND2_X1 _578_ (.A1(_049_),
    .A2(_052_),
    .ZN(_227_));
 INV_X1 _579_ (.A(_410_),
    .ZN(_244_));
 NAND2_X1 _580_ (.A1(_045_),
    .A2(_052_),
    .ZN(_254_));
 NAND2_X1 _581_ (.A1(_045_),
    .A2(_053_),
    .ZN(_263_));
 NAND2_X1 _582_ (.A1(_048_),
    .A2(_050_),
    .ZN(_228_));
 NAND2_X1 _583_ (.A1(_043_),
    .A2(_050_),
    .ZN(_255_));
 NAND2_X1 _584_ (.A1(_043_),
    .A2(_052_),
    .ZN(_264_));
 NAND2_X1 _585_ (.A1(_052_),
    .A2(_054_),
    .ZN(_286_));
 NAND2_X1 _586_ (.A1(_051_),
    .A2(_053_),
    .ZN(_229_));
 NAND2_X1 _587_ (.A1(_041_),
    .A2(_056_),
    .ZN(_275_));
 NAND2_X1 _588_ (.A1(_050_),
    .A2(_051_),
    .ZN(_287_));
 INV_X1 _589_ (.A(_226_),
    .ZN(_238_));
 INV_X1 _590_ (.A(_236_),
    .ZN(_412_));
 INV_X1 _591_ (.A(_243_),
    .ZN(_250_));
 INV_X1 _592_ (.A(_327_),
    .ZN(_328_));
 INV_X1 _593_ (.A(_337_),
    .ZN(_339_));
 INV_X1 _594_ (.A(_346_),
    .ZN(_347_));
 INV_X1 _595_ (.A(_356_),
    .ZN(_357_));
 INV_X1 _596_ (.A(_363_),
    .ZN(_364_));
 INV_X1 _597_ (.A(_372_),
    .ZN(_373_));
 INV_X1 _598_ (.A(_379_),
    .ZN(_380_));
 INV_X1 _599_ (.A(_389_),
    .ZN(_390_));
 INV_X1 _600_ (.A(_399_),
    .ZN(_400_));
 INV_X1 _601_ (.A(_225_),
    .ZN(_219_));
 INV_X1 _602_ (.A(_251_),
    .ZN(_245_));
 INV_X1 _603_ (.A(_326_),
    .ZN(_350_));
 INV_X1 _604_ (.A(_345_),
    .ZN(_367_));
 INV_X1 _605_ (.A(_362_),
    .ZN(_383_));
 INV_X1 _606_ (.A(_378_),
    .ZN(_393_));
 INV_X1 _607_ (.A(_388_),
    .ZN(_403_));
 INV_X1 _608_ (.A(_221_),
    .ZN(_232_));
 INV_X1 _609_ (.A(_253_),
    .ZN(_249_));
 INV_X1 _610_ (.A(_246_),
    .ZN(_411_));
 INV_X1 _611_ (.A(_266_),
    .ZN(_259_));
 XOR2_X1 _612_ (.A(\b_reg[0] ),
    .B(_043_),
    .Z(_064_));
 AND2_X2 _613_ (.A1(_056_),
    .A2(_064_),
    .ZN(_428_));
 INV_X1 _614_ (.A(_311_),
    .ZN(_442_));
 INV_X1 _615_ (.A(_352_),
    .ZN(_448_));
 INV_X1 _616_ (.A(_351_),
    .ZN(_454_));
 INV_X1 _617_ (.A(net38),
    .ZN(_458_));
 INV_X1 _618_ (.A(_385_),
    .ZN(_461_));
 INV_X1 _619_ (.A(_395_),
    .ZN(_470_));
 INV_X1 _620_ (.A(_405_),
    .ZN(_478_));
 AND2_X1 _621_ (.A1(_041_),
    .A2(_044_),
    .ZN(_224_));
 AND2_X1 _622_ (.A1(_041_),
    .A2(_046_),
    .ZN(_242_));
 INV_X1 _623_ (.A(_230_),
    .ZN(_407_));
 INV_X1 _624_ (.A(_257_),
    .ZN(_260_));
 INV_X1 _625_ (.A(_247_),
    .ZN(_419_));
 INV_X1 _626_ (.A(_289_),
    .ZN(_423_));
 INV_X1 _627_ (.A(_292_),
    .ZN(_293_));
 INV_X1 _628_ (.A(_312_),
    .ZN(_434_));
 INV_X1 _629_ (.A(_300_),
    .ZN(_324_));
 INV_X1 _630_ (.A(_332_),
    .ZN(_443_));
 INV_X1 _631_ (.A(_317_),
    .ZN(_344_));
 INV_X1 _632_ (.A(_331_),
    .ZN(_449_));
 INV_X1 _633_ (.A(_369_),
    .ZN(_455_));
 INV_X1 _634_ (.A(_368_),
    .ZN(_462_));
 INV_X1 _635_ (.A(_374_),
    .ZN(_465_));
 INV_X1 _636_ (.A(_384_),
    .ZN(_471_));
 NOR2_X1 _637_ (.A1(_056_),
    .A2(_055_),
    .ZN(_474_));
 INV_X1 _638_ (.A(_394_),
    .ZN(_479_));
 INV_X1 _639_ (.A(_267_),
    .ZN(_488_));
 INV_X1 _640_ (.A(_414_),
    .ZN(_270_));
 INV_X1 _641_ (.A(_424_),
    .ZN(_290_));
 INV_X1 _642_ (.A(_430_),
    .ZN(_302_));
 INV_X2 _643_ (.A(_439_),
    .ZN(_320_));
 INV_X1 _644_ (.A(_433_),
    .ZN(_305_));
 INV_X1 _645_ (.A(_415_),
    .ZN(_269_));
 MUX2_X1 _646_ (.A(net1),
    .B(_053_),
    .S(_063_),
    .Z(_065_));
 AND2_X1 _647_ (.A1(_038_),
    .A2(_065_),
    .ZN(_003_));
 MUX2_X1 _648_ (.A(net2),
    .B(_052_),
    .S(_063_),
    .Z(_066_));
 AND2_X1 _649_ (.A1(_038_),
    .A2(_066_),
    .ZN(_004_));
 MUX2_X1 _650_ (.A(net3),
    .B(_050_),
    .S(_063_),
    .Z(_067_));
 AND2_X1 _651_ (.A1(_038_),
    .A2(_067_),
    .ZN(_005_));
 MUX2_X1 _652_ (.A(net4),
    .B(_047_),
    .S(_063_),
    .Z(_068_));
 AND2_X1 _653_ (.A1(_038_),
    .A2(_068_),
    .ZN(_006_));
 MUX2_X1 _654_ (.A(net5),
    .B(_046_),
    .S(_063_),
    .Z(_069_));
 AND2_X1 _655_ (.A1(_038_),
    .A2(_069_),
    .ZN(_007_));
 MUX2_X1 _656_ (.A(net6),
    .B(_044_),
    .S(_063_),
    .Z(_070_));
 AND2_X1 _657_ (.A1(_038_),
    .A2(_070_),
    .ZN(_008_));
 MUX2_X1 _658_ (.A(net7),
    .B(_042_),
    .S(_063_),
    .Z(_071_));
 AND2_X1 _659_ (.A1(_038_),
    .A2(_071_),
    .ZN(_009_));
 MUX2_X1 _660_ (.A(net8),
    .B(_056_),
    .S(_063_),
    .Z(_072_));
 AND2_X1 _661_ (.A1(_038_),
    .A2(_072_),
    .ZN(_010_));
 MUX2_X1 _662_ (.A(net9),
    .B(_041_),
    .S(_062_),
    .Z(_073_));
 AND2_X1 _663_ (.A1(_038_),
    .A2(_073_),
    .ZN(_011_));
 MUX2_X1 _664_ (.A(net10),
    .B(_043_),
    .S(_062_),
    .Z(_074_));
 AND2_X1 _665_ (.A1(_037_),
    .A2(_074_),
    .ZN(_012_));
 MUX2_X1 _666_ (.A(net11),
    .B(_045_),
    .S(_062_),
    .Z(_075_));
 AND2_X1 _667_ (.A1(_037_),
    .A2(_075_),
    .ZN(_013_));
 MUX2_X1 _668_ (.A(net12),
    .B(_048_),
    .S(_062_),
    .Z(_076_));
 AND2_X1 _669_ (.A1(_037_),
    .A2(_076_),
    .ZN(_014_));
 MUX2_X1 _670_ (.A(net13),
    .B(_049_),
    .S(_062_),
    .Z(_077_));
 AND2_X1 _671_ (.A1(_037_),
    .A2(_077_),
    .ZN(_015_));
 MUX2_X1 _672_ (.A(net14),
    .B(_051_),
    .S(_062_),
    .Z(_078_));
 AND2_X1 _673_ (.A1(_037_),
    .A2(_078_),
    .ZN(_016_));
 MUX2_X1 _674_ (.A(net15),
    .B(_054_),
    .S(_062_),
    .Z(_079_));
 AND2_X1 _675_ (.A1(_037_),
    .A2(_079_),
    .ZN(_017_));
 MUX2_X1 _676_ (.A(net16),
    .B(\b_reg[7] ),
    .S(_062_),
    .Z(_080_));
 AND2_X1 _677_ (.A1(_037_),
    .A2(_080_),
    .ZN(_018_));
 OAI21_X1 _678_ (.A(_037_),
    .B1(net19),
    .B2(_040_),
    .ZN(_081_));
 AOI21_X1 _679_ (.A(\state[1] ),
    .B1(net19),
    .B2(_063_),
    .ZN(_082_));
 NOR2_X1 _680_ (.A1(_081_),
    .A2(_082_),
    .ZN(_019_));
 INV_X2 _681_ (.A(_058_),
    .ZN(_083_));
 CLKBUF_X3 _682_ (.A(_083_),
    .Z(_084_));
 NAND2_X1 _683_ (.A1(_084_),
    .A2(net20),
    .ZN(_085_));
 CLKBUF_X3 _684_ (.A(_058_),
    .Z(_086_));
 NAND3_X1 _685_ (.A1(_041_),
    .A2(_053_),
    .A3(_086_),
    .ZN(_087_));
 AOI21_X1 _686_ (.A(_061_),
    .B1(_085_),
    .B2(_087_),
    .ZN(_020_));
 NOR2_X1 _687_ (.A1(_060_),
    .A2(_058_),
    .ZN(_088_));
 NAND2_X1 _688_ (.A1(net21),
    .A2(_088_),
    .ZN(_089_));
 INV_X1 _689_ (.A(_444_),
    .ZN(_090_));
 BUF_X4 _690_ (.A(_436_),
    .Z(_091_));
 AOI21_X1 _691_ (.A(_435_),
    .B1(_425_),
    .B2(_091_),
    .ZN(_092_));
 BUF_X4 _692_ (.A(_445_),
    .Z(_093_));
 INV_X1 _693_ (.A(_093_),
    .ZN(_094_));
 OAI21_X1 _694_ (.A(_090_),
    .B1(_092_),
    .B2(_094_),
    .ZN(_095_));
 INV_X1 _695_ (.A(_426_),
    .ZN(_096_));
 NAND2_X1 _696_ (.A1(_091_),
    .A2(_093_),
    .ZN(_097_));
 AOI21_X1 _697_ (.A(_416_),
    .B1(_422_),
    .B2(_417_),
    .ZN(_098_));
 NOR3_X1 _698_ (.A1(_096_),
    .A2(_097_),
    .A3(_098_),
    .ZN(_099_));
 NOR2_X1 _699_ (.A1(_095_),
    .A2(_099_),
    .ZN(_100_));
 XOR2_X1 _700_ (.A(net36),
    .B(_100_),
    .Z(_101_));
 OAI21_X1 _701_ (.A(_089_),
    .B1(_101_),
    .B2(_059_),
    .ZN(_021_));
 NAND2_X1 _702_ (.A1(_084_),
    .A2(net22),
    .ZN(_102_));
 BUF_X2 _703_ (.A(_457_),
    .Z(_103_));
 INV_X1 _704_ (.A(_425_),
    .ZN(_104_));
 OAI21_X2 _705_ (.A(_104_),
    .B1(_271_),
    .B2(_096_),
    .ZN(_105_));
 AND3_X1 _706_ (.A1(_091_),
    .A2(_093_),
    .A3(_451_),
    .ZN(_106_));
 AOI21_X1 _707_ (.A(_444_),
    .B1(_435_),
    .B2(_093_),
    .ZN(_107_));
 INV_X1 _708_ (.A(_107_),
    .ZN(_108_));
 AOI221_X2 _709_ (.A(_450_),
    .B1(_105_),
    .B2(_106_),
    .C1(_108_),
    .C2(_451_),
    .ZN(_109_));
 XNOR2_X1 _710_ (.A(_103_),
    .B(_109_),
    .ZN(_110_));
 NAND2_X1 _711_ (.A1(_086_),
    .A2(_110_),
    .ZN(_111_));
 AOI21_X1 _712_ (.A(_061_),
    .B1(_102_),
    .B2(_111_),
    .ZN(_022_));
 NAND2_X1 _713_ (.A1(_084_),
    .A2(net23),
    .ZN(_112_));
 BUF_X2 _714_ (.A(_464_),
    .Z(_113_));
 AOI21_X2 _715_ (.A(_456_),
    .B1(_450_),
    .B2(_103_),
    .ZN(_114_));
 AND2_X1 _716_ (.A1(_451_),
    .A2(_103_),
    .ZN(_115_));
 OAI21_X1 _717_ (.A(_115_),
    .B1(_099_),
    .B2(_095_),
    .ZN(_116_));
 AOI21_X1 _718_ (.A(_113_),
    .B1(_114_),
    .B2(_116_),
    .ZN(_117_));
 AND3_X1 _719_ (.A1(_113_),
    .A2(_114_),
    .A3(_116_),
    .ZN(_118_));
 OAI21_X1 _720_ (.A(_086_),
    .B1(_117_),
    .B2(_118_),
    .ZN(_119_));
 AOI21_X1 _721_ (.A(_061_),
    .B1(_112_),
    .B2(_119_),
    .ZN(_023_));
 BUF_X2 _722_ (.A(_473_),
    .Z(_120_));
 AOI21_X2 _723_ (.A(_463_),
    .B1(_456_),
    .B2(_113_),
    .ZN(_121_));
 NAND3_X1 _724_ (.A1(_058_),
    .A2(_120_),
    .A3(_121_),
    .ZN(_122_));
 OR2_X1 _725_ (.A1(_083_),
    .A2(_120_),
    .ZN(_123_));
 NAND2_X1 _726_ (.A1(_103_),
    .A2(_113_),
    .ZN(_124_));
 NOR2_X1 _727_ (.A1(_109_),
    .A2(_124_),
    .ZN(_125_));
 MUX2_X1 _728_ (.A(_122_),
    .B(_123_),
    .S(_125_),
    .Z(_126_));
 NOR2_X1 _729_ (.A1(_121_),
    .A2(_123_),
    .ZN(_127_));
 AOI21_X1 _730_ (.A(_127_),
    .B1(net24),
    .B2(_083_),
    .ZN(_128_));
 AOI21_X1 _731_ (.A(_061_),
    .B1(_126_),
    .B2(_128_),
    .ZN(_024_));
 NAND2_X1 _732_ (.A1(net25),
    .A2(_088_),
    .ZN(_129_));
 AOI21_X1 _733_ (.A(_472_),
    .B1(_463_),
    .B2(_120_),
    .ZN(_130_));
 NAND2_X1 _734_ (.A1(_113_),
    .A2(_120_),
    .ZN(_131_));
 NAND3_X1 _735_ (.A1(_113_),
    .A2(_120_),
    .A3(_115_),
    .ZN(_132_));
 OAI221_X2 _736_ (.A(_130_),
    .B1(_131_),
    .B2(_114_),
    .C1(_100_),
    .C2(_132_),
    .ZN(_133_));
 XNOR2_X1 _737_ (.A(_481_),
    .B(_133_),
    .ZN(_134_));
 OAI21_X1 _738_ (.A(_129_),
    .B1(_134_),
    .B2(_059_),
    .ZN(_025_));
 XOR2_X1 _739_ (.A(_398_),
    .B(_477_),
    .Z(_135_));
 XNOR2_X1 _740_ (.A(_401_),
    .B(_404_),
    .ZN(_136_));
 XNOR2_X1 _741_ (.A(_135_),
    .B(_136_),
    .ZN(_137_));
 XNOR2_X1 _742_ (.A(_475_),
    .B(_467_),
    .ZN(_138_));
 XNOR2_X1 _743_ (.A(_137_),
    .B(_138_),
    .ZN(_139_));
 OAI21_X1 _744_ (.A(_113_),
    .B1(_456_),
    .B2(_103_),
    .ZN(_140_));
 OR2_X1 _745_ (.A1(_472_),
    .A2(_480_),
    .ZN(_141_));
 NOR2_X1 _746_ (.A1(_463_),
    .A2(_141_),
    .ZN(_142_));
 NAND2_X1 _747_ (.A1(_140_),
    .A2(_142_),
    .ZN(_143_));
 OAI221_X2 _748_ (.A(_143_),
    .B1(_480_),
    .B2(_481_),
    .C1(_120_),
    .C2(_141_),
    .ZN(_144_));
 INV_X1 _749_ (.A(_121_),
    .ZN(_145_));
 AOI21_X1 _750_ (.A(_141_),
    .B1(_145_),
    .B2(_120_),
    .ZN(_146_));
 AND2_X1 _751_ (.A1(_109_),
    .A2(_146_),
    .ZN(_147_));
 OAI211_X2 _752_ (.A(_000_),
    .B(_139_),
    .C1(_144_),
    .C2(_147_),
    .ZN(_148_));
 OR4_X1 _753_ (.A1(_059_),
    .A2(_139_),
    .A3(_144_),
    .A4(_147_),
    .ZN(_149_));
 NAND2_X1 _754_ (.A1(net26),
    .A2(_088_),
    .ZN(_150_));
 NAND3_X1 _755_ (.A1(_148_),
    .A2(_149_),
    .A3(_150_),
    .ZN(_026_));
 NAND2_X1 _756_ (.A1(_086_),
    .A2(_487_),
    .ZN(_151_));
 NAND2_X1 _757_ (.A1(_084_),
    .A2(net27),
    .ZN(_152_));
 AOI21_X1 _758_ (.A(_061_),
    .B1(_151_),
    .B2(_152_),
    .ZN(_027_));
 NAND2_X1 _759_ (.A1(_086_),
    .A2(_490_),
    .ZN(_153_));
 NAND2_X1 _760_ (.A1(_084_),
    .A2(net28),
    .ZN(_154_));
 AOI21_X1 _761_ (.A(_061_),
    .B1(_153_),
    .B2(_154_),
    .ZN(_028_));
 NAND2_X1 _762_ (.A1(_086_),
    .A2(_492_),
    .ZN(_155_));
 NAND2_X1 _763_ (.A1(_084_),
    .A2(net29),
    .ZN(_156_));
 AOI21_X1 _764_ (.A(_061_),
    .B1(_155_),
    .B2(_156_),
    .ZN(_029_));
 NAND2_X1 _765_ (.A1(_086_),
    .A2(_493_),
    .ZN(_157_));
 NAND2_X1 _766_ (.A1(_084_),
    .A2(net30),
    .ZN(_158_));
 AOI21_X1 _767_ (.A(_061_),
    .B1(_157_),
    .B2(_158_),
    .ZN(_030_));
 NAND2_X1 _768_ (.A1(_086_),
    .A2(_483_),
    .ZN(_159_));
 NAND2_X1 _769_ (.A1(_084_),
    .A2(net31),
    .ZN(_160_));
 AOI21_X1 _770_ (.A(_060_),
    .B1(_159_),
    .B2(_160_),
    .ZN(_031_));
 NOR2_X1 _771_ (.A1(_083_),
    .A2(_272_),
    .ZN(_161_));
 AOI21_X1 _772_ (.A(_161_),
    .B1(net32),
    .B2(_083_),
    .ZN(_162_));
 NOR2_X1 _773_ (.A1(_061_),
    .A2(_162_),
    .ZN(_032_));
 NAND2_X1 _774_ (.A1(_084_),
    .A2(net33),
    .ZN(_163_));
 XNOR2_X1 _775_ (.A(_426_),
    .B(_271_),
    .ZN(_164_));
 NAND2_X1 _776_ (.A1(_086_),
    .A2(_164_),
    .ZN(_165_));
 AOI21_X1 _777_ (.A(_060_),
    .B1(_163_),
    .B2(_165_),
    .ZN(_033_));
 NAND2_X1 _778_ (.A1(_083_),
    .A2(net34),
    .ZN(_166_));
 OAI21_X1 _779_ (.A(_104_),
    .B1(_098_),
    .B2(_096_),
    .ZN(_167_));
 XNOR2_X1 _780_ (.A(_091_),
    .B(_167_),
    .ZN(_168_));
 OAI21_X1 _781_ (.A(_166_),
    .B1(_168_),
    .B2(_083_),
    .ZN(_169_));
 AND2_X1 _782_ (.A1(_037_),
    .A2(_169_),
    .ZN(_034_));
 NAND2_X1 _783_ (.A1(_084_),
    .A2(net35),
    .ZN(_170_));
 AOI21_X1 _784_ (.A(_435_),
    .B1(_105_),
    .B2(_091_),
    .ZN(_171_));
 XNOR2_X1 _785_ (.A(_093_),
    .B(_171_),
    .ZN(_172_));
 NAND2_X1 _786_ (.A1(_086_),
    .A2(_172_),
    .ZN(_173_));
 AOI21_X1 _787_ (.A(_060_),
    .B1(_170_),
    .B2(_173_),
    .ZN(_035_));
 FA_X1 _788_ (.A(_209_),
    .B(_210_),
    .CI(_211_),
    .CO(_212_),
    .S(_213_));
 FA_X1 _789_ (.A(_214_),
    .B(_215_),
    .CI(_216_),
    .CO(_217_),
    .S(_218_));
 FA_X1 _790_ (.A(_218_),
    .B(_219_),
    .CI(_213_),
    .CO(_220_),
    .S(_221_));
 FA_X1 _791_ (.A(_222_),
    .B(_223_),
    .CI(_224_),
    .CO(_225_),
    .S(_226_));
 FA_X1 _792_ (.A(_227_),
    .B(_228_),
    .CI(_229_),
    .CO(_230_),
    .S(_231_));
 FA_X1 _793_ (.A(_232_),
    .B(_233_),
    .CI(_234_),
    .CO(_235_),
    .S(_236_));
 FA_X1 _794_ (.A(_237_),
    .B(_238_),
    .CI(_231_),
    .CO(_234_),
    .S(_239_));
 FA_X1 _795_ (.A(_240_),
    .B(_241_),
    .CI(_242_),
    .CO(_237_),
    .S(_243_));
 FA_X1 _796_ (.A(_244_),
    .B(_245_),
    .CI(_239_),
    .CO(_246_),
    .S(_247_));
 FA_X1 _797_ (.A(_248_),
    .B(_249_),
    .CI(_250_),
    .CO(_251_),
    .S(_252_));
 FA_X1 _798_ (.A(_254_),
    .B(_255_),
    .CI(_256_),
    .CO(_253_),
    .S(_257_));
 FA_X1 _799_ (.A(_258_),
    .B(_259_),
    .CI(_260_),
    .CO(_261_),
    .S(_262_));
 FA_X1 _800_ (.A(_263_),
    .B(_264_),
    .CI(_265_),
    .CO(_266_),
    .S(_267_));
 FA_X1 _801_ (.A(_268_),
    .B(_269_),
    .CI(_270_),
    .CO(_271_),
    .S(_272_));
 FA_X1 _802_ (.A(_273_),
    .B(_274_),
    .CI(_275_),
    .CO(_276_),
    .S(_277_));
 FA_X1 _803_ (.A(_278_),
    .B(_279_),
    .CI(_280_),
    .CO(_281_),
    .S(_282_));
 FA_X1 _804_ (.A(_277_),
    .B(_282_),
    .CI(_212_),
    .CO(_283_),
    .S(_284_));
 FA_X1 _805_ (.A(_285_),
    .B(_286_),
    .CI(_287_),
    .CO(_288_),
    .S(_289_));
 FA_X1 _806_ (.A(_284_),
    .B(_220_),
    .CI(_290_),
    .CO(_291_),
    .S(_292_));
 FA_X1 _807_ (.A(_235_),
    .B(_293_),
    .CI(_294_),
    .CO(_295_),
    .S(_296_));
 FA_X1 _808_ (.A(_297_),
    .B(_298_),
    .CI(_299_),
    .CO(_300_),
    .S(_301_));
 FA_X1 _809_ (.A(_276_),
    .B(_301_),
    .CI(_302_),
    .CO(_303_),
    .S(_304_));
 FA_X1 _810_ (.A(_305_),
    .B(_281_),
    .CI(_288_),
    .CO(_306_),
    .S(_307_));
 FA_X1 _811_ (.A(_304_),
    .B(_283_),
    .CI(_307_),
    .CO(_308_),
    .S(_309_));
 FA_X1 _812_ (.A(_310_),
    .B(_291_),
    .CI(_309_),
    .CO(_311_),
    .S(_312_));
 FA_X1 _813_ (.A(_314_),
    .B(_315_),
    .CI(_316_),
    .CO(_317_),
    .S(_318_));
 FA_X1 _814_ (.A(_318_),
    .B(_319_),
    .CI(_320_),
    .CO(_321_),
    .S(_322_));
 FA_X1 _815_ (.A(_323_),
    .B(_324_),
    .CI(_325_),
    .CO(_326_),
    .S(_327_));
 FA_X1 _816_ (.A(_322_),
    .B(_328_),
    .CI(_303_),
    .CO(_329_),
    .S(_330_));
 FA_X1 _817_ (.A(_330_),
    .B(_308_),
    .CI(_306_),
    .CO(_331_),
    .S(_332_));
 FA_X1 _818_ (.A(_333_),
    .B(_334_),
    .CI(_335_),
    .CO(_336_),
    .S(_337_));
 FA_X1 _819_ (.A(_338_),
    .B(_339_),
    .CI(_320_),
    .CO(_340_),
    .S(_341_));
 FA_X1 _820_ (.A(_342_),
    .B(_343_),
    .CI(_344_),
    .CO(_345_),
    .S(_346_));
 FA_X1 _821_ (.A(_321_),
    .B(_347_),
    .CI(_341_),
    .CO(_348_),
    .S(_349_));
 FA_X1 _822_ (.A(_349_),
    .B(_350_),
    .CI(_329_),
    .CO(_351_),
    .S(_352_));
 FA_X1 _823_ (.A(_333_),
    .B(_353_),
    .CI(_354_),
    .CO(_355_),
    .S(_356_));
 FA_X1 _824_ (.A(_338_),
    .B(_357_),
    .CI(_320_),
    .CO(_358_),
    .S(_359_));
 FA_X1 _825_ (.A(_336_),
    .B(_360_),
    .CI(_361_),
    .CO(_362_),
    .S(_363_));
 FA_X1 _826_ (.A(_340_),
    .B(_359_),
    .CI(_364_),
    .CO(_365_),
    .S(_366_));
 FA_X1 _827_ (.A(_348_),
    .B(_366_),
    .CI(_367_),
    .CO(_368_),
    .S(_369_));
 FA_X1 _828_ (.A(_333_),
    .B(_354_),
    .CI(_370_),
    .CO(_371_),
    .S(_372_));
 FA_X1 _829_ (.A(_338_),
    .B(_320_),
    .CI(_373_),
    .CO(_374_),
    .S(_375_));
 FA_X1 _830_ (.A(_355_),
    .B(_376_),
    .CI(_377_),
    .CO(_378_),
    .S(_379_));
 FA_X1 _831_ (.A(_375_),
    .B(_358_),
    .CI(_380_),
    .CO(_381_),
    .S(_382_));
 FA_X1 _832_ (.A(_382_),
    .B(_365_),
    .CI(_383_),
    .CO(_384_),
    .S(_385_));
 FA_X1 _833_ (.A(_371_),
    .B(_386_),
    .CI(_387_),
    .CO(_388_),
    .S(_389_));
 FA_X1 _834_ (.A(net37),
    .B(_374_),
    .CI(_390_),
    .CO(_391_),
    .S(_392_));
 FA_X1 _835_ (.A(_392_),
    .B(_381_),
    .CI(_393_),
    .CO(_394_),
    .S(_395_));
 FA_X1 _836_ (.A(_371_),
    .B(_396_),
    .CI(_397_),
    .CO(_398_),
    .S(_399_));
 FA_X1 _837_ (.A(net37),
    .B(_374_),
    .CI(_400_),
    .CO(_401_),
    .S(_402_));
 FA_X1 _838_ (.A(_403_),
    .B(_402_),
    .CI(_391_),
    .CO(_404_),
    .S(_405_));
 HA_X1 _839_ (.A(_406_),
    .B(_407_),
    .CO(_294_),
    .S(_233_));
 HA_X1 _840_ (.A(_408_),
    .B(_409_),
    .CO(_410_),
    .S(_248_));
 HA_X1 _841_ (.A(_411_),
    .B(_412_),
    .CO(_413_),
    .S(_414_));
 HA_X1 _842_ (.A(_415_),
    .B(_414_),
    .CO(_416_),
    .S(_417_));
 HA_X1 _843_ (.A(_418_),
    .B(_419_),
    .CO(_415_),
    .S(_420_));
 HA_X1 _844_ (.A(_261_),
    .B(_252_),
    .CO(_418_),
    .S(_421_));
 HA_X1 _845_ (.A(_217_),
    .B(_423_),
    .CO(_313_),
    .S(_424_));
 HA_X1 _846_ (.A(_296_),
    .B(_413_),
    .CO(_425_),
    .S(_426_));
 HA_X1 _847_ (.A(_427_),
    .B(_428_),
    .CO(_429_),
    .S(_430_));
 HA_X1 _848_ (.A(_431_),
    .B(_432_),
    .CO(_325_),
    .S(_433_));
 HA_X1 _849_ (.A(_295_),
    .B(_434_),
    .CO(_435_),
    .S(_436_));
 HA_X1 _850_ (.A(_428_),
    .B(_437_),
    .CO(_438_),
    .S(_439_));
 HA_X1 _851_ (.A(_440_),
    .B(_441_),
    .CO(_342_),
    .S(_323_));
 HA_X1 _852_ (.A(_442_),
    .B(_443_),
    .CO(_444_),
    .S(_445_));
 HA_X1 _853_ (.A(_446_),
    .B(_447_),
    .CO(_360_),
    .S(_343_));
 HA_X1 _854_ (.A(_449_),
    .B(_448_),
    .CO(_450_),
    .S(_451_));
 HA_X1 _855_ (.A(_452_),
    .B(_453_),
    .CO(_377_),
    .S(_361_));
 HA_X1 _856_ (.A(_454_),
    .B(_455_),
    .CO(_456_),
    .S(_457_));
 HA_X1 _857_ (.A(_459_),
    .B(_460_),
    .CO(_386_),
    .S(_376_));
 HA_X1 _858_ (.A(_461_),
    .B(_462_),
    .CO(_463_),
    .S(_464_));
 HA_X1 _859_ (.A(_458_),
    .B(_465_),
    .CO(_466_),
    .S(_467_));
 HA_X1 _860_ (.A(_468_),
    .B(_469_),
    .CO(_396_),
    .S(_387_));
 HA_X1 _861_ (.A(_470_),
    .B(_471_),
    .CO(_472_),
    .S(_473_));
 HA_X1 _862_ (.A(_468_),
    .B(_474_),
    .CO(_475_),
    .S(_397_));
 HA_X1 _863_ (.A(_371_),
    .B(_397_),
    .CO(_476_),
    .S(_477_));
 HA_X1 _864_ (.A(_478_),
    .B(_479_),
    .CO(_480_),
    .S(_481_));
 HA_X1 _865_ (.A(_482_),
    .B(_420_),
    .CO(_422_),
    .S(_483_));
 HA_X1 _866_ (.A(_484_),
    .B(_485_),
    .CO(_486_),
    .S(_487_));
 HA_X1 _867_ (.A(_486_),
    .B(_488_),
    .CO(_489_),
    .S(_490_));
 HA_X1 _868_ (.A(_489_),
    .B(_262_),
    .CO(_491_),
    .S(_492_));
 HA_X1 _869_ (.A(_491_),
    .B(_421_),
    .CO(_482_),
    .S(_493_));
 DFF_X1 \a_reg[0]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\a_reg[0] ),
    .QN(_205_));
 DFF_X1 \a_reg[1]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\a_reg[1] ),
    .QN(_204_));
 DFF_X1 \a_reg[2]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\a_reg[2] ),
    .QN(_203_));
 DFF_X1 \a_reg[3]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\a_reg[3] ),
    .QN(_202_));
 DFF_X1 \a_reg[4]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\a_reg[4] ),
    .QN(_201_));
 DFF_X1 \a_reg[5]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\a_reg[5] ),
    .QN(_200_));
 DFF_X1 \a_reg[6]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\a_reg[6] ),
    .QN(_199_));
 DFF_X1 \a_reg[7]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\a_reg[7] ),
    .QN(_198_));
 DFF_X1 \b_reg[0]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\b_reg[0] ),
    .QN(_197_));
 DFF_X1 \b_reg[1]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\b_reg[1] ),
    .QN(_196_));
 DFF_X1 \b_reg[2]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\b_reg[2] ),
    .QN(_195_));
 DFF_X1 \b_reg[3]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\b_reg[3] ),
    .QN(_194_));
 DFF_X1 \b_reg[4]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\b_reg[4] ),
    .QN(_193_));
 DFF_X1 \b_reg[5]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\b_reg[5] ),
    .QN(_192_));
 DFF_X1 \b_reg[6]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\b_reg[6] ),
    .QN(_191_));
 DFF_X1 \b_reg[7]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\b_reg[7] ),
    .QN(_273_));
 DFF_X1 \done$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net19),
    .QN(_190_));
 DFF_X1 \product[0]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net20),
    .QN(_189_));
 DFF_X1 \product[10]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net21),
    .QN(_188_));
 DFF_X1 \product[11]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net22),
    .QN(_187_));
 DFF_X1 \product[12]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net23),
    .QN(_186_));
 DFF_X1 \product[13]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net24),
    .QN(_185_));
 DFF_X1 \product[14]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net25),
    .QN(_184_));
 DFF_X1 \product[15]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net26),
    .QN(_183_));
 DFF_X1 \product[1]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net27),
    .QN(_182_));
 DFF_X1 \product[2]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net28),
    .QN(_181_));
 DFF_X1 \product[3]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net29),
    .QN(_180_));
 DFF_X1 \product[4]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net30),
    .QN(_179_));
 DFF_X1 \product[5]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net31),
    .QN(_178_));
 DFF_X1 \product[6]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net32),
    .QN(_177_));
 DFF_X1 \product[7]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net33),
    .QN(_176_));
 DFF_X1 \product[8]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net34),
    .QN(_175_));
 DFF_X1 \product[9]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net35),
    .QN(_206_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[0] ),
    .QN(_207_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\state[1] ),
    .QN(_208_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\state[2] ),
    .QN(_174_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_53 ();
 BUF_X1 input1 (.A(multiplicand[0]),
    .Z(net1));
 BUF_X1 input2 (.A(multiplicand[1]),
    .Z(net2));
 BUF_X1 input3 (.A(multiplicand[2]),
    .Z(net3));
 BUF_X1 input4 (.A(multiplicand[3]),
    .Z(net4));
 BUF_X1 input5 (.A(multiplicand[4]),
    .Z(net5));
 BUF_X1 input6 (.A(multiplicand[5]),
    .Z(net6));
 BUF_X1 input7 (.A(multiplicand[6]),
    .Z(net7));
 BUF_X1 input8 (.A(multiplicand[7]),
    .Z(net8));
 BUF_X1 input9 (.A(multiplier[0]),
    .Z(net9));
 BUF_X1 input10 (.A(multiplier[1]),
    .Z(net10));
 BUF_X1 input11 (.A(multiplier[2]),
    .Z(net11));
 BUF_X1 input12 (.A(multiplier[3]),
    .Z(net12));
 BUF_X1 input13 (.A(multiplier[4]),
    .Z(net13));
 BUF_X1 input14 (.A(multiplier[5]),
    .Z(net14));
 BUF_X1 input15 (.A(multiplier[6]),
    .Z(net15));
 BUF_X1 input16 (.A(multiplier[7]),
    .Z(net16));
 BUF_X1 input17 (.A(rst_n),
    .Z(net17));
 BUF_X1 input18 (.A(start),
    .Z(net18));
 BUF_X1 output19 (.A(net19),
    .Z(done));
 BUF_X1 output20 (.A(net20),
    .Z(product[0]));
 BUF_X1 output21 (.A(net21),
    .Z(product[10]));
 BUF_X1 output22 (.A(net22),
    .Z(product[11]));
 BUF_X1 output23 (.A(net23),
    .Z(product[12]));
 BUF_X1 output24 (.A(net24),
    .Z(product[13]));
 BUF_X1 output25 (.A(net25),
    .Z(product[14]));
 BUF_X1 output26 (.A(net26),
    .Z(product[15]));
 BUF_X1 output27 (.A(net27),
    .Z(product[1]));
 BUF_X1 output28 (.A(net28),
    .Z(product[2]));
 BUF_X1 output29 (.A(net29),
    .Z(product[3]));
 BUF_X1 output30 (.A(net30),
    .Z(product[4]));
 BUF_X1 output31 (.A(net31),
    .Z(product[5]));
 BUF_X1 output32 (.A(net32),
    .Z(product[6]));
 BUF_X1 output33 (.A(net33),
    .Z(product[7]));
 BUF_X1 output34 (.A(net34),
    .Z(product[8]));
 BUF_X1 output35 (.A(net35),
    .Z(product[9]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X1 clkload0 (.A(clknet_2_1__leaf_clk));
 INV_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 BUF_X1 rebuffer1 (.A(_451_),
    .Z(net36));
 BUF_X4 rebuffer2 (.A(_375_),
    .Z(net37));
 BUF_X1 rebuffer3 (.A(net37),
    .Z(net38));
 FILLCELL_X8 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_9 ();
 FILLCELL_X2 FILLER_0_13 ();
 FILLCELL_X4 FILLER_0_39 ();
 FILLCELL_X1 FILLER_0_43 ();
 FILLCELL_X1 FILLER_0_47 ();
 FILLCELL_X2 FILLER_0_51 ();
 FILLCELL_X1 FILLER_0_53 ();
 FILLCELL_X4 FILLER_0_60 ();
 FILLCELL_X2 FILLER_0_64 ();
 FILLCELL_X4 FILLER_0_69 ();
 FILLCELL_X4 FILLER_0_76 ();
 FILLCELL_X4 FILLER_0_90 ();
 FILLCELL_X2 FILLER_0_131 ();
 FILLCELL_X1 FILLER_0_133 ();
 FILLCELL_X16 FILLER_0_137 ();
 FILLCELL_X2 FILLER_0_153 ();
 FILLCELL_X1 FILLER_0_155 ();
 FILLCELL_X4 FILLER_0_159 ();
 FILLCELL_X32 FILLER_0_166 ();
 FILLCELL_X4 FILLER_0_198 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_19 ();
 FILLCELL_X2 FILLER_1_24 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X1 FILLER_1_80 ();
 FILLCELL_X8 FILLER_1_109 ();
 FILLCELL_X4 FILLER_1_117 ();
 FILLCELL_X2 FILLER_1_121 ();
 FILLCELL_X1 FILLER_1_123 ();
 FILLCELL_X4 FILLER_1_132 ();
 FILLCELL_X4 FILLER_1_147 ();
 FILLCELL_X2 FILLER_1_151 ();
 FILLCELL_X1 FILLER_1_153 ();
 FILLCELL_X16 FILLER_1_186 ();
 FILLCELL_X4 FILLER_2_4 ();
 FILLCELL_X16 FILLER_2_12 ();
 FILLCELL_X8 FILLER_2_28 ();
 FILLCELL_X4 FILLER_2_36 ();
 FILLCELL_X2 FILLER_2_40 ();
 FILLCELL_X4 FILLER_2_63 ();
 FILLCELL_X8 FILLER_2_89 ();
 FILLCELL_X4 FILLER_2_101 ();
 FILLCELL_X8 FILLER_2_122 ();
 FILLCELL_X4 FILLER_2_139 ();
 FILLCELL_X1 FILLER_2_164 ();
 FILLCELL_X16 FILLER_2_176 ();
 FILLCELL_X8 FILLER_2_192 ();
 FILLCELL_X2 FILLER_2_200 ();
 FILLCELL_X1 FILLER_3_1 ();
 FILLCELL_X4 FILLER_3_30 ();
 FILLCELL_X1 FILLER_3_34 ();
 FILLCELL_X2 FILLER_3_39 ();
 FILLCELL_X4 FILLER_3_62 ();
 FILLCELL_X2 FILLER_3_66 ();
 FILLCELL_X1 FILLER_3_68 ();
 FILLCELL_X8 FILLER_3_73 ();
 FILLCELL_X4 FILLER_3_81 ();
 FILLCELL_X2 FILLER_3_85 ();
 FILLCELL_X4 FILLER_3_94 ();
 FILLCELL_X2 FILLER_3_98 ();
 FILLCELL_X1 FILLER_3_100 ();
 FILLCELL_X16 FILLER_3_108 ();
 FILLCELL_X8 FILLER_3_140 ();
 FILLCELL_X4 FILLER_3_148 ();
 FILLCELL_X1 FILLER_3_152 ();
 FILLCELL_X8 FILLER_3_159 ();
 FILLCELL_X4 FILLER_3_167 ();
 FILLCELL_X1 FILLER_3_171 ();
 FILLCELL_X8 FILLER_3_193 ();
 FILLCELL_X1 FILLER_3_201 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_25 ();
 FILLCELL_X1 FILLER_4_29 ();
 FILLCELL_X4 FILLER_4_47 ();
 FILLCELL_X2 FILLER_4_51 ();
 FILLCELL_X4 FILLER_4_61 ();
 FILLCELL_X4 FILLER_4_86 ();
 FILLCELL_X1 FILLER_4_90 ();
 FILLCELL_X16 FILLER_4_119 ();
 FILLCELL_X2 FILLER_4_135 ();
 FILLCELL_X4 FILLER_4_140 ();
 FILLCELL_X2 FILLER_4_144 ();
 FILLCELL_X8 FILLER_4_162 ();
 FILLCELL_X2 FILLER_4_170 ();
 FILLCELL_X1 FILLER_4_172 ();
 FILLCELL_X8 FILLER_4_190 ();
 FILLCELL_X4 FILLER_4_198 ();
 FILLCELL_X8 FILLER_5_41 ();
 FILLCELL_X2 FILLER_5_49 ();
 FILLCELL_X8 FILLER_5_72 ();
 FILLCELL_X1 FILLER_5_80 ();
 FILLCELL_X4 FILLER_5_98 ();
 FILLCELL_X2 FILLER_5_102 ();
 FILLCELL_X4 FILLER_5_123 ();
 FILLCELL_X1 FILLER_5_127 ();
 FILLCELL_X4 FILLER_5_159 ();
 FILLCELL_X1 FILLER_5_163 ();
 FILLCELL_X1 FILLER_5_171 ();
 FILLCELL_X8 FILLER_5_176 ();
 FILLCELL_X2 FILLER_5_184 ();
 FILLCELL_X4 FILLER_5_190 ();
 FILLCELL_X1 FILLER_5_194 ();
 FILLCELL_X4 FILLER_5_198 ();
 FILLCELL_X2 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_28 ();
 FILLCELL_X1 FILLER_6_32 ();
 FILLCELL_X32 FILLER_6_36 ();
 FILLCELL_X8 FILLER_6_68 ();
 FILLCELL_X1 FILLER_6_81 ();
 FILLCELL_X4 FILLER_6_88 ();
 FILLCELL_X2 FILLER_6_92 ();
 FILLCELL_X1 FILLER_6_94 ();
 FILLCELL_X4 FILLER_6_108 ();
 FILLCELL_X4 FILLER_6_141 ();
 FILLCELL_X4 FILLER_6_161 ();
 FILLCELL_X2 FILLER_6_171 ();
 FILLCELL_X1 FILLER_6_177 ();
 FILLCELL_X16 FILLER_6_182 ();
 FILLCELL_X4 FILLER_6_198 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_17 ();
 FILLCELL_X1 FILLER_7_23 ();
 FILLCELL_X16 FILLER_7_27 ();
 FILLCELL_X8 FILLER_7_43 ();
 FILLCELL_X2 FILLER_7_51 ();
 FILLCELL_X4 FILLER_7_57 ();
 FILLCELL_X1 FILLER_7_61 ();
 FILLCELL_X4 FILLER_7_66 ();
 FILLCELL_X2 FILLER_7_70 ();
 FILLCELL_X1 FILLER_7_72 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X1 FILLER_7_93 ();
 FILLCELL_X16 FILLER_7_110 ();
 FILLCELL_X2 FILLER_7_126 ();
 FILLCELL_X4 FILLER_7_132 ();
 FILLCELL_X1 FILLER_7_136 ();
 FILLCELL_X16 FILLER_7_183 ();
 FILLCELL_X2 FILLER_7_199 ();
 FILLCELL_X1 FILLER_7_201 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_17 ();
 FILLCELL_X1 FILLER_8_44 ();
 FILLCELL_X4 FILLER_8_49 ();
 FILLCELL_X1 FILLER_8_53 ();
 FILLCELL_X4 FILLER_8_64 ();
 FILLCELL_X4 FILLER_8_71 ();
 FILLCELL_X1 FILLER_8_77 ();
 FILLCELL_X8 FILLER_8_81 ();
 FILLCELL_X4 FILLER_8_89 ();
 FILLCELL_X2 FILLER_8_93 ();
 FILLCELL_X2 FILLER_8_117 ();
 FILLCELL_X1 FILLER_8_135 ();
 FILLCELL_X8 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_162 ();
 FILLCELL_X2 FILLER_8_166 ();
 FILLCELL_X1 FILLER_8_168 ();
 FILLCELL_X16 FILLER_8_179 ();
 FILLCELL_X4 FILLER_8_195 ();
 FILLCELL_X2 FILLER_8_199 ();
 FILLCELL_X1 FILLER_8_201 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_17 ();
 FILLCELL_X1 FILLER_9_22 ();
 FILLCELL_X4 FILLER_9_26 ();
 FILLCELL_X2 FILLER_9_30 ();
 FILLCELL_X8 FILLER_9_79 ();
 FILLCELL_X4 FILLER_9_87 ();
 FILLCELL_X1 FILLER_9_96 ();
 FILLCELL_X4 FILLER_9_101 ();
 FILLCELL_X4 FILLER_9_107 ();
 FILLCELL_X2 FILLER_9_111 ();
 FILLCELL_X1 FILLER_9_113 ();
 FILLCELL_X32 FILLER_9_130 ();
 FILLCELL_X1 FILLER_9_162 ();
 FILLCELL_X2 FILLER_9_165 ();
 FILLCELL_X16 FILLER_9_183 ();
 FILLCELL_X2 FILLER_9_199 ();
 FILLCELL_X1 FILLER_9_201 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_33 ();
 FILLCELL_X1 FILLER_10_37 ();
 FILLCELL_X4 FILLER_10_42 ();
 FILLCELL_X2 FILLER_10_50 ();
 FILLCELL_X4 FILLER_10_54 ();
 FILLCELL_X2 FILLER_10_74 ();
 FILLCELL_X2 FILLER_10_86 ();
 FILLCELL_X1 FILLER_10_88 ();
 FILLCELL_X2 FILLER_10_92 ();
 FILLCELL_X1 FILLER_10_94 ();
 FILLCELL_X16 FILLER_10_107 ();
 FILLCELL_X4 FILLER_10_123 ();
 FILLCELL_X1 FILLER_10_127 ();
 FILLCELL_X4 FILLER_10_144 ();
 FILLCELL_X16 FILLER_10_154 ();
 FILLCELL_X1 FILLER_10_170 ();
 FILLCELL_X1 FILLER_10_175 ();
 FILLCELL_X1 FILLER_10_178 ();
 FILLCELL_X2 FILLER_10_182 ();
 FILLCELL_X8 FILLER_10_194 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_5 ();
 FILLCELL_X1 FILLER_11_32 ();
 FILLCELL_X16 FILLER_11_49 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X2 FILLER_11_73 ();
 FILLCELL_X1 FILLER_11_75 ();
 FILLCELL_X8 FILLER_11_78 ();
 FILLCELL_X2 FILLER_11_86 ();
 FILLCELL_X2 FILLER_11_102 ();
 FILLCELL_X2 FILLER_11_109 ();
 FILLCELL_X1 FILLER_11_111 ();
 FILLCELL_X2 FILLER_11_116 ();
 FILLCELL_X1 FILLER_11_118 ();
 FILLCELL_X2 FILLER_11_122 ();
 FILLCELL_X4 FILLER_11_126 ();
 FILLCELL_X1 FILLER_11_130 ();
 FILLCELL_X8 FILLER_11_134 ();
 FILLCELL_X2 FILLER_11_142 ();
 FILLCELL_X1 FILLER_11_182 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_5 ();
 FILLCELL_X4 FILLER_12_12 ();
 FILLCELL_X1 FILLER_12_16 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X4 FILLER_12_49 ();
 FILLCELL_X4 FILLER_12_55 ();
 FILLCELL_X2 FILLER_12_59 ();
 FILLCELL_X1 FILLER_12_61 ();
 FILLCELL_X4 FILLER_12_64 ();
 FILLCELL_X1 FILLER_12_68 ();
 FILLCELL_X4 FILLER_12_85 ();
 FILLCELL_X1 FILLER_12_89 ();
 FILLCELL_X2 FILLER_12_93 ();
 FILLCELL_X1 FILLER_12_95 ();
 FILLCELL_X2 FILLER_12_101 ();
 FILLCELL_X2 FILLER_12_111 ();
 FILLCELL_X1 FILLER_12_113 ();
 FILLCELL_X2 FILLER_12_144 ();
 FILLCELL_X1 FILLER_12_146 ();
 FILLCELL_X4 FILLER_12_149 ();
 FILLCELL_X2 FILLER_12_156 ();
 FILLCELL_X8 FILLER_12_162 ();
 FILLCELL_X4 FILLER_12_170 ();
 FILLCELL_X1 FILLER_12_174 ();
 FILLCELL_X8 FILLER_12_191 ();
 FILLCELL_X2 FILLER_12_199 ();
 FILLCELL_X1 FILLER_12_201 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_9 ();
 FILLCELL_X2 FILLER_13_13 ();
 FILLCELL_X16 FILLER_13_19 ();
 FILLCELL_X4 FILLER_13_35 ();
 FILLCELL_X2 FILLER_13_39 ();
 FILLCELL_X2 FILLER_13_43 ();
 FILLCELL_X1 FILLER_13_45 ();
 FILLCELL_X4 FILLER_13_62 ();
 FILLCELL_X2 FILLER_13_66 ();
 FILLCELL_X1 FILLER_13_68 ();
 FILLCELL_X8 FILLER_13_71 ();
 FILLCELL_X2 FILLER_13_79 ();
 FILLCELL_X4 FILLER_13_99 ();
 FILLCELL_X16 FILLER_13_119 ();
 FILLCELL_X2 FILLER_13_135 ();
 FILLCELL_X8 FILLER_13_147 ();
 FILLCELL_X4 FILLER_13_155 ();
 FILLCELL_X2 FILLER_13_159 ();
 FILLCELL_X4 FILLER_13_171 ();
 FILLCELL_X8 FILLER_13_177 ();
 FILLCELL_X4 FILLER_13_185 ();
 FILLCELL_X8 FILLER_13_191 ();
 FILLCELL_X2 FILLER_13_199 ();
 FILLCELL_X1 FILLER_13_201 ();
 FILLCELL_X2 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_9 ();
 FILLCELL_X1 FILLER_14_11 ();
 FILLCELL_X2 FILLER_14_30 ();
 FILLCELL_X4 FILLER_14_48 ();
 FILLCELL_X2 FILLER_14_52 ();
 FILLCELL_X1 FILLER_14_54 ();
 FILLCELL_X2 FILLER_14_71 ();
 FILLCELL_X1 FILLER_14_73 ();
 FILLCELL_X4 FILLER_14_90 ();
 FILLCELL_X1 FILLER_14_94 ();
 FILLCELL_X8 FILLER_14_115 ();
 FILLCELL_X2 FILLER_14_123 ();
 FILLCELL_X1 FILLER_14_125 ();
 FILLCELL_X4 FILLER_14_128 ();
 FILLCELL_X2 FILLER_14_132 ();
 FILLCELL_X1 FILLER_14_134 ();
 FILLCELL_X4 FILLER_14_183 ();
 FILLCELL_X8 FILLER_14_189 ();
 FILLCELL_X4 FILLER_14_197 ();
 FILLCELL_X1 FILLER_14_201 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_37 ();
 FILLCELL_X2 FILLER_15_41 ();
 FILLCELL_X1 FILLER_15_43 ();
 FILLCELL_X16 FILLER_15_51 ();
 FILLCELL_X8 FILLER_15_67 ();
 FILLCELL_X8 FILLER_15_91 ();
 FILLCELL_X4 FILLER_15_99 ();
 FILLCELL_X2 FILLER_15_103 ();
 FILLCELL_X1 FILLER_15_105 ();
 FILLCELL_X8 FILLER_15_124 ();
 FILLCELL_X4 FILLER_15_132 ();
 FILLCELL_X2 FILLER_15_136 ();
 FILLCELL_X1 FILLER_15_138 ();
 FILLCELL_X16 FILLER_15_141 ();
 FILLCELL_X2 FILLER_15_157 ();
 FILLCELL_X1 FILLER_15_159 ();
 FILLCELL_X4 FILLER_15_164 ();
 FILLCELL_X2 FILLER_15_172 ();
 FILLCELL_X4 FILLER_15_198 ();
 FILLCELL_X2 FILLER_16_1 ();
 FILLCELL_X1 FILLER_16_3 ();
 FILLCELL_X4 FILLER_16_10 ();
 FILLCELL_X2 FILLER_16_14 ();
 FILLCELL_X1 FILLER_16_16 ();
 FILLCELL_X1 FILLER_16_21 ();
 FILLCELL_X4 FILLER_16_25 ();
 FILLCELL_X1 FILLER_16_29 ();
 FILLCELL_X1 FILLER_16_62 ();
 FILLCELL_X2 FILLER_16_81 ();
 FILLCELL_X1 FILLER_16_83 ();
 FILLCELL_X2 FILLER_16_102 ();
 FILLCELL_X8 FILLER_16_106 ();
 FILLCELL_X4 FILLER_16_114 ();
 FILLCELL_X1 FILLER_16_118 ();
 FILLCELL_X1 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_140 ();
 FILLCELL_X4 FILLER_16_148 ();
 FILLCELL_X2 FILLER_16_152 ();
 FILLCELL_X1 FILLER_16_154 ();
 FILLCELL_X8 FILLER_16_175 ();
 FILLCELL_X2 FILLER_16_183 ();
 FILLCELL_X4 FILLER_16_197 ();
 FILLCELL_X1 FILLER_16_201 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_9 ();
 FILLCELL_X16 FILLER_17_43 ();
 FILLCELL_X2 FILLER_17_59 ();
 FILLCELL_X8 FILLER_17_65 ();
 FILLCELL_X4 FILLER_17_73 ();
 FILLCELL_X1 FILLER_17_77 ();
 FILLCELL_X8 FILLER_17_88 ();
 FILLCELL_X4 FILLER_17_96 ();
 FILLCELL_X1 FILLER_17_100 ();
 FILLCELL_X8 FILLER_17_103 ();
 FILLCELL_X4 FILLER_17_111 ();
 FILLCELL_X2 FILLER_17_115 ();
 FILLCELL_X1 FILLER_17_117 ();
 FILLCELL_X1 FILLER_17_125 ();
 FILLCELL_X16 FILLER_17_135 ();
 FILLCELL_X2 FILLER_17_151 ();
 FILLCELL_X8 FILLER_17_163 ();
 FILLCELL_X1 FILLER_17_171 ();
 FILLCELL_X4 FILLER_17_174 ();
 FILLCELL_X1 FILLER_17_178 ();
 FILLCELL_X2 FILLER_17_199 ();
 FILLCELL_X1 FILLER_17_201 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_9 ();
 FILLCELL_X8 FILLER_18_16 ();
 FILLCELL_X2 FILLER_18_24 ();
 FILLCELL_X1 FILLER_18_26 ();
 FILLCELL_X4 FILLER_18_29 ();
 FILLCELL_X1 FILLER_18_33 ();
 FILLCELL_X4 FILLER_18_36 ();
 FILLCELL_X2 FILLER_18_40 ();
 FILLCELL_X2 FILLER_18_44 ();
 FILLCELL_X8 FILLER_18_48 ();
 FILLCELL_X4 FILLER_18_56 ();
 FILLCELL_X2 FILLER_18_60 ();
 FILLCELL_X1 FILLER_18_62 ();
 FILLCELL_X4 FILLER_18_73 ();
 FILLCELL_X2 FILLER_18_77 ();
 FILLCELL_X8 FILLER_18_83 ();
 FILLCELL_X8 FILLER_18_108 ();
 FILLCELL_X1 FILLER_18_128 ();
 FILLCELL_X2 FILLER_18_135 ();
 FILLCELL_X1 FILLER_18_137 ();
 FILLCELL_X1 FILLER_18_148 ();
 FILLCELL_X8 FILLER_18_151 ();
 FILLCELL_X1 FILLER_18_159 ();
 FILLCELL_X4 FILLER_18_164 ();
 FILLCELL_X2 FILLER_18_168 ();
 FILLCELL_X8 FILLER_18_180 ();
 FILLCELL_X1 FILLER_18_188 ();
 FILLCELL_X2 FILLER_18_199 ();
 FILLCELL_X1 FILLER_18_201 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_43 ();
 FILLCELL_X4 FILLER_19_62 ();
 FILLCELL_X2 FILLER_19_70 ();
 FILLCELL_X1 FILLER_19_72 ();
 FILLCELL_X1 FILLER_19_77 ();
 FILLCELL_X1 FILLER_19_82 ();
 FILLCELL_X2 FILLER_19_102 ();
 FILLCELL_X1 FILLER_19_150 ();
 FILLCELL_X8 FILLER_19_191 ();
 FILLCELL_X2 FILLER_19_199 ();
 FILLCELL_X1 FILLER_19_201 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_33 ();
 FILLCELL_X2 FILLER_20_41 ();
 FILLCELL_X2 FILLER_20_77 ();
 FILLCELL_X1 FILLER_20_90 ();
 FILLCELL_X8 FILLER_20_108 ();
 FILLCELL_X4 FILLER_20_116 ();
 FILLCELL_X2 FILLER_20_139 ();
 FILLCELL_X1 FILLER_20_141 ();
 FILLCELL_X1 FILLER_20_158 ();
 FILLCELL_X8 FILLER_20_164 ();
 FILLCELL_X2 FILLER_20_172 ();
 FILLCELL_X1 FILLER_20_174 ();
 FILLCELL_X4 FILLER_20_178 ();
 FILLCELL_X2 FILLER_20_185 ();
 FILLCELL_X8 FILLER_20_191 ();
 FILLCELL_X2 FILLER_20_199 ();
 FILLCELL_X1 FILLER_20_201 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_17 ();
 FILLCELL_X1 FILLER_21_25 ();
 FILLCELL_X4 FILLER_21_52 ();
 FILLCELL_X2 FILLER_21_60 ();
 FILLCELL_X2 FILLER_21_75 ();
 FILLCELL_X4 FILLER_21_81 ();
 FILLCELL_X1 FILLER_21_85 ();
 FILLCELL_X1 FILLER_21_95 ();
 FILLCELL_X16 FILLER_21_100 ();
 FILLCELL_X8 FILLER_21_116 ();
 FILLCELL_X8 FILLER_21_127 ();
 FILLCELL_X4 FILLER_21_135 ();
 FILLCELL_X2 FILLER_21_139 ();
 FILLCELL_X16 FILLER_21_144 ();
 FILLCELL_X1 FILLER_21_160 ();
 FILLCELL_X8 FILLER_21_165 ();
 FILLCELL_X4 FILLER_21_173 ();
 FILLCELL_X1 FILLER_21_177 ();
 FILLCELL_X2 FILLER_21_199 ();
 FILLCELL_X1 FILLER_21_201 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_33 ();
 FILLCELL_X2 FILLER_22_41 ();
 FILLCELL_X1 FILLER_22_43 ();
 FILLCELL_X16 FILLER_22_52 ();
 FILLCELL_X2 FILLER_22_85 ();
 FILLCELL_X4 FILLER_22_90 ();
 FILLCELL_X2 FILLER_22_94 ();
 FILLCELL_X2 FILLER_22_101 ();
 FILLCELL_X4 FILLER_22_106 ();
 FILLCELL_X1 FILLER_22_110 ();
 FILLCELL_X4 FILLER_22_115 ();
 FILLCELL_X2 FILLER_22_119 ();
 FILLCELL_X1 FILLER_22_121 ();
 FILLCELL_X16 FILLER_22_126 ();
 FILLCELL_X2 FILLER_22_142 ();
 FILLCELL_X2 FILLER_22_149 ();
 FILLCELL_X2 FILLER_22_171 ();
 FILLCELL_X1 FILLER_22_173 ();
 FILLCELL_X2 FILLER_22_191 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X8 FILLER_23_33 ();
 FILLCELL_X4 FILLER_23_41 ();
 FILLCELL_X1 FILLER_23_45 ();
 FILLCELL_X8 FILLER_23_50 ();
 FILLCELL_X4 FILLER_23_58 ();
 FILLCELL_X2 FILLER_23_62 ();
 FILLCELL_X8 FILLER_23_71 ();
 FILLCELL_X4 FILLER_23_100 ();
 FILLCELL_X2 FILLER_23_104 ();
 FILLCELL_X1 FILLER_23_106 ();
 FILLCELL_X4 FILLER_23_127 ();
 FILLCELL_X32 FILLER_23_151 ();
 FILLCELL_X4 FILLER_23_183 ();
 FILLCELL_X4 FILLER_23_191 ();
 FILLCELL_X1 FILLER_23_195 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X8 FILLER_24_17 ();
 FILLCELL_X4 FILLER_24_25 ();
 FILLCELL_X2 FILLER_24_29 ();
 FILLCELL_X8 FILLER_24_51 ();
 FILLCELL_X2 FILLER_24_63 ();
 FILLCELL_X1 FILLER_24_65 ();
 FILLCELL_X2 FILLER_24_71 ();
 FILLCELL_X1 FILLER_24_73 ();
 FILLCELL_X8 FILLER_24_82 ();
 FILLCELL_X2 FILLER_24_90 ();
 FILLCELL_X8 FILLER_24_113 ();
 FILLCELL_X4 FILLER_24_121 ();
 FILLCELL_X4 FILLER_24_132 ();
 FILLCELL_X2 FILLER_24_136 ();
 FILLCELL_X4 FILLER_24_149 ();
 FILLCELL_X8 FILLER_24_161 ();
 FILLCELL_X4 FILLER_24_169 ();
 FILLCELL_X4 FILLER_24_177 ();
 FILLCELL_X1 FILLER_24_181 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_33 ();
 FILLCELL_X1 FILLER_25_52 ();
 FILLCELL_X8 FILLER_25_87 ();
 FILLCELL_X8 FILLER_25_187 ();
 FILLCELL_X4 FILLER_25_195 ();
 FILLCELL_X2 FILLER_25_199 ();
 FILLCELL_X1 FILLER_25_201 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X8 FILLER_26_33 ();
 FILLCELL_X2 FILLER_26_41 ();
 FILLCELL_X1 FILLER_26_53 ();
 FILLCELL_X4 FILLER_26_57 ();
 FILLCELL_X1 FILLER_26_67 ();
 FILLCELL_X8 FILLER_26_71 ();
 FILLCELL_X1 FILLER_26_79 ();
 FILLCELL_X16 FILLER_26_83 ();
 FILLCELL_X4 FILLER_26_99 ();
 FILLCELL_X2 FILLER_26_103 ();
 FILLCELL_X1 FILLER_26_105 ();
 FILLCELL_X1 FILLER_26_115 ();
 FILLCELL_X8 FILLER_26_119 ();
 FILLCELL_X2 FILLER_26_127 ();
 FILLCELL_X1 FILLER_26_129 ();
 FILLCELL_X8 FILLER_26_133 ();
 FILLCELL_X4 FILLER_26_150 ();
 FILLCELL_X2 FILLER_26_154 ();
 FILLCELL_X2 FILLER_26_163 ();
 FILLCELL_X2 FILLER_26_168 ();
 FILLCELL_X1 FILLER_26_170 ();
 FILLCELL_X16 FILLER_26_177 ();
 FILLCELL_X8 FILLER_26_193 ();
 FILLCELL_X1 FILLER_26_201 ();
endmodule
