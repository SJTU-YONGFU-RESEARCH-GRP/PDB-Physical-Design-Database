module parameterized_i2c_master (ack_error,
    busy,
    clk,
    done,
    read,
    rst_n,
    scl,
    scl_internal_debug,
    sda,
    sda_internal_debug,
    start,
    stop,
    write,
    addr,
    bit_counter_debug,
    data_in,
    data_out,
    phase,
    shift_reg_debug,
    state);
 output ack_error;
 output busy;
 input clk;
 output done;
 input read;
 input rst_n;
 output scl;
 output scl_internal_debug;
 inout sda;
 output sda_internal_debug;
 input start;
 input stop;
 input write;
 input [6:0] addr;
 output [2:0] bit_counter_debug;
 input [7:0] data_in;
 output [7:0] data_out;
 output [1:0] phase;
 output [7:0] shift_reg_debug;
 output [3:0] state;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire clknet_0_clk;
 wire cmd_read;
 wire cmd_write;
 wire \divider_counter[0] ;
 wire \divider_counter[1] ;
 wire \divider_counter[2] ;
 wire \divider_counter[3] ;
 wire \divider_counter[4] ;
 wire \divider_counter[5] ;
 wire \divider_counter[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net54;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _290_ (.I(net23),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _291_ (.I(\divider_counter[0] ),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _292_ (.A1(\divider_counter[5] ),
    .A2(\divider_counter[4] ),
    .A3(\divider_counter[3] ),
    .A4(\divider_counter[2] ),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _293_ (.A1(\divider_counter[1] ),
    .A2(\divider_counter[0] ),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _294_ (.A1(\divider_counter[6] ),
    .A2(_039_),
    .A3(_040_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _295_ (.A1(_267_),
    .A2(_041_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _296_ (.A1(\divider_counter[6] ),
    .A2(_039_),
    .A3(_040_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _297_ (.A1(_270_),
    .A2(_042_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _298_ (.A1(\divider_counter[2] ),
    .A2(_269_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _299_ (.A1(_041_),
    .A2(_043_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _300_ (.A1(\divider_counter[2] ),
    .A2(_040_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _301_ (.A1(\divider_counter[3] ),
    .A2(_044_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _302_ (.I(_269_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _303_ (.A1(\divider_counter[3] ),
    .A2(\divider_counter[2] ),
    .A3(_045_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _304_ (.A1(\divider_counter[4] ),
    .A2(_046_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _305_ (.A1(_041_),
    .A2(_047_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _306_ (.A1(\divider_counter[4] ),
    .A2(\divider_counter[3] ),
    .A3(\divider_counter[2] ),
    .A4(_040_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _307_ (.A1(\divider_counter[5] ),
    .A2(_048_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _308_ (.A1(_045_),
    .A2(_040_),
    .B(_039_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _309_ (.A1(_045_),
    .A2(_039_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _310_ (.I0(_049_),
    .I1(_050_),
    .S(\divider_counter[6] ),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _311_ (.I(net51),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _312_ (.I(_051_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _313_ (.I(_052_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _314_ (.I(_287_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _315_ (.I(net49),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _316_ (.A1(_055_),
    .A2(net48),
    .A3(net50),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _317_ (.A1(_053_),
    .A2(_054_),
    .A3(_042_),
    .A4(_056_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _318_ (.I(net36),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _319_ (.I(\divider_counter[1] ),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _320_ (.I(net24),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _321_ (.I(net37),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _322_ (.I(net50),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _323_ (.A1(net49),
    .A2(net48),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _324_ (.A1(_057_),
    .A2(_283_),
    .A3(_058_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _325_ (.I(net48),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _326_ (.I(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _327_ (.A1(_061_),
    .A2(_057_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _328_ (.I(net48),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _329_ (.A1(_063_),
    .A2(net50),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _330_ (.A1(_283_),
    .A2(_064_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _331_ (.I(_055_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _332_ (.A1(_062_),
    .A2(_065_),
    .B(_066_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _333_ (.A1(net51),
    .A2(net50),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _334_ (.I(net19),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _335_ (.A1(_055_),
    .A2(_063_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _336_ (.A1(_069_),
    .A2(_070_),
    .B1(_058_),
    .B2(_283_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _337_ (.A1(_059_),
    .A2(_067_),
    .B1(_068_),
    .B2(_071_),
    .C(_042_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _338_ (.A1(_053_),
    .A2(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _339_ (.A1(net22),
    .A2(_073_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _340_ (.I(net49),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _341_ (.I(_074_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _342_ (.I(_063_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _343_ (.A1(_075_),
    .A2(_057_),
    .B(_052_),
    .C(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _344_ (.A1(net23),
    .A2(_077_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _345_ (.I(net50),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _346_ (.A1(_061_),
    .A2(_079_),
    .B(_066_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _347_ (.A1(_061_),
    .A2(_079_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _348_ (.A1(_080_),
    .A2(_081_),
    .B(_052_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _349_ (.I(cmd_read),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _350_ (.A1(net20),
    .A2(_083_),
    .B(_058_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _351_ (.A1(_063_),
    .A2(_051_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _352_ (.A1(_055_),
    .A2(_079_),
    .B(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _353_ (.A1(net24),
    .A2(net25),
    .A3(net23),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _354_ (.A1(_051_),
    .A2(_057_),
    .A3(_084_),
    .B1(_086_),
    .B2(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _355_ (.I0(_082_),
    .I1(_088_),
    .S(_054_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _356_ (.I(cmd_write),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _357_ (.A1(_090_),
    .A2(net20),
    .B(_074_),
    .C(_079_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _358_ (.A1(_074_),
    .A2(net50),
    .A3(_287_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _359_ (.A1(_091_),
    .A2(_092_),
    .B(_060_),
    .C(_051_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _360_ (.A1(_051_),
    .A2(net50),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _361_ (.A1(_287_),
    .A2(net22),
    .A3(_058_),
    .A4(_094_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _362_ (.A1(_041_),
    .A2(_095_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _363_ (.I0(_283_),
    .I1(_287_),
    .S(net50),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _364_ (.A1(_055_),
    .A2(_060_),
    .A3(_097_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _365_ (.I(_098_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _366_ (.I(_079_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _367_ (.A1(_055_),
    .A2(_063_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _368_ (.I(_051_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _369_ (.I(_102_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _370_ (.A1(_100_),
    .A2(net19),
    .A3(_101_),
    .B(_103_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _371_ (.A1(_093_),
    .A2(_096_),
    .A3(_099_),
    .A4(_104_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _372_ (.A1(_089_),
    .A2(_105_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _373_ (.I0(net23),
    .I1(_078_),
    .S(_106_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _374_ (.A1(_274_),
    .A2(_077_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _375_ (.I0(net24),
    .I1(_107_),
    .S(_106_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _376_ (.I(net25),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _377_ (.A1(_069_),
    .A2(_056_),
    .B(_051_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _378_ (.A1(_098_),
    .A2(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _379_ (.A1(_093_),
    .A2(_096_),
    .A3(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _380_ (.A1(_273_),
    .A2(_086_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _381_ (.A1(_089_),
    .A2(_111_),
    .A3(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _382_ (.A1(net25),
    .A2(_273_),
    .A3(_077_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _383_ (.A1(_089_),
    .A2(_111_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _384_ (.A1(_108_),
    .A2(_113_),
    .B1(_114_),
    .B2(_115_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _385_ (.A1(net19),
    .A2(_042_),
    .A3(_070_),
    .A4(_094_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _386_ (.I0(cmd_read),
    .I1(net17),
    .S(_116_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _387_ (.I0(cmd_write),
    .I1(net21),
    .S(_116_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _388_ (.I(_287_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _389_ (.A1(_055_),
    .A2(_060_),
    .A3(_102_),
    .A4(_079_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _390_ (.I(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _391_ (.A1(_117_),
    .A2(_041_),
    .A3(_087_),
    .A4(_119_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _392_ (.I0(net27),
    .I1(net40),
    .S(_120_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _393_ (.I0(net28),
    .I1(net41),
    .S(_120_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _394_ (.I0(net29),
    .I1(net42),
    .S(_120_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _395_ (.I0(net30),
    .I1(net43),
    .S(_120_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _396_ (.I0(net31),
    .I1(net44),
    .S(_120_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _397_ (.I0(net32),
    .I1(net45),
    .S(_120_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _398_ (.I0(net33),
    .I1(net46),
    .S(_120_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _399_ (.I0(net34),
    .I1(net47),
    .S(_120_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _400_ (.I(net39),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _401_ (.A1(net24),
    .A2(net25),
    .A3(net23),
    .B(_287_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _402_ (.I(net20),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _403_ (.A1(_057_),
    .A2(_054_),
    .A3(_123_),
    .B(_103_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _404_ (.A1(_079_),
    .A2(net20),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _405_ (.I0(_094_),
    .I1(_125_),
    .S(_066_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _406_ (.A1(_066_),
    .A2(_124_),
    .B1(_126_),
    .B2(_061_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _407_ (.A1(_076_),
    .A2(_054_),
    .B(_066_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _408_ (.A1(_076_),
    .A2(_287_),
    .A3(_123_),
    .A4(cmd_read),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _409_ (.A1(_103_),
    .A2(_100_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _410_ (.A1(_061_),
    .A2(_054_),
    .B(_075_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _411_ (.A1(_128_),
    .A2(_129_),
    .B(_130_),
    .C(_131_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _412_ (.A1(_121_),
    .A2(_087_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _413_ (.A1(_054_),
    .A2(_070_),
    .A3(_130_),
    .A4(_133_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _414_ (.A1(cmd_read),
    .A2(net47),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _415_ (.A1(_103_),
    .A2(_058_),
    .A3(_135_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _416_ (.A1(_103_),
    .A2(_101_),
    .B(_054_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _417_ (.A1(_075_),
    .A2(_283_),
    .B(_052_),
    .C(_061_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _418_ (.A1(_051_),
    .A2(_283_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _419_ (.A1(_117_),
    .A2(_283_),
    .B1(_101_),
    .B2(_139_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _420_ (.A1(_136_),
    .A2(_137_),
    .B1(_138_),
    .B2(_140_),
    .C(_057_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _421_ (.A1(_127_),
    .A2(_132_),
    .A3(_134_),
    .A4(_141_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _422_ (.A1(_063_),
    .A2(_079_),
    .B(_051_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _423_ (.I(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _424_ (.A1(cmd_write),
    .A2(_123_),
    .Z(_145_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _425_ (.A1(_075_),
    .A2(_064_),
    .Z(_146_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _426_ (.A1(net16),
    .A2(_145_),
    .A3(_146_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _427_ (.I0(net40),
    .I1(net41),
    .I2(net44),
    .I3(net45),
    .S0(net23),
    .S1(net25),
    .Z(_148_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _428_ (.A1(net24),
    .A2(_148_),
    .Z(_149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _429_ (.I0(net46),
    .I1(net47),
    .S(net23),
    .Z(_150_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _430_ (.A1(_272_),
    .A2(_108_),
    .A3(_150_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _431_ (.I0(net42),
    .I1(net43),
    .S(net23),
    .Z(_152_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _432_ (.A1(_272_),
    .A2(net25),
    .A3(_152_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _433_ (.A1(_103_),
    .A2(_079_),
    .A3(_117_),
    .A4(_070_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _434_ (.A1(_149_),
    .A2(_151_),
    .A3(_153_),
    .A4(_154_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _435_ (.A1(_144_),
    .A2(_147_),
    .A3(_155_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _436_ (.I(_282_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _437_ (.A1(_080_),
    .A2(_081_),
    .B(_052_),
    .C(_157_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _438_ (.A1(_075_),
    .A2(_100_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _439_ (.A1(_075_),
    .A2(_100_),
    .A3(_285_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _440_ (.A1(_061_),
    .A2(_051_),
    .A3(_287_),
    .A4(_281_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _441_ (.A1(_159_),
    .A2(_160_),
    .B(_161_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _442_ (.A1(_054_),
    .A2(_087_),
    .A3(_118_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _443_ (.A1(_096_),
    .A2(_158_),
    .A3(_162_),
    .A4(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _444_ (.A1(_122_),
    .A2(_142_),
    .A3(_156_),
    .B(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _445_ (.A1(_096_),
    .A2(_158_),
    .A3(_162_),
    .A4(_163_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _446_ (.A1(_061_),
    .A2(_094_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _447_ (.A1(_054_),
    .A2(net47),
    .Z(_168_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _448_ (.A1(_066_),
    .A2(_167_),
    .A3(_168_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _449_ (.A1(_166_),
    .A2(_142_),
    .A3(_156_),
    .A4(_169_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _450_ (.A1(_121_),
    .A2(_165_),
    .B(_170_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _451_ (.A1(_055_),
    .A2(_060_),
    .A3(_283_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _452_ (.A1(_055_),
    .A2(_060_),
    .B(_079_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _453_ (.A1(net49),
    .A2(net48),
    .A3(_287_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _454_ (.A1(net22),
    .A2(_083_),
    .A3(_068_),
    .A4(_173_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _455_ (.A1(_055_),
    .A2(_060_),
    .A3(_057_),
    .A4(_122_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _456_ (.A1(_171_),
    .A2(_172_),
    .B(_174_),
    .C(_175_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _457_ (.A1(_093_),
    .A2(_096_),
    .A3(_110_),
    .A4(_176_),
    .Z(_177_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _458_ (.I(_177_),
    .Z(_178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _459_ (.I(net17),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _460_ (.A1(_066_),
    .A2(_100_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _461_ (.A1(_066_),
    .A2(_057_),
    .Z(_181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _462_ (.I0(cmd_read),
    .I1(net9),
    .S(_100_),
    .Z(_182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _463_ (.A1(net9),
    .A2(_181_),
    .B1(_182_),
    .B2(_075_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _464_ (.A1(_179_),
    .A2(_180_),
    .B1(_183_),
    .B2(_053_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _465_ (.A1(_103_),
    .A2(_101_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _466_ (.A1(_076_),
    .A2(_184_),
    .B1(_185_),
    .B2(net17),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _467_ (.A1(net25),
    .A2(_273_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _468_ (.A1(_274_),
    .A2(_087_),
    .A3(_187_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _469_ (.A1(_118_),
    .A2(_188_),
    .Z(_189_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _470_ (.A1(_189_),
    .A2(_178_),
    .B(net40),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _471_ (.A1(_178_),
    .A2(_186_),
    .B(_190_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _472_ (.I(net2),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _473_ (.A1(_075_),
    .A2(_064_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _474_ (.A1(_103_),
    .A2(_192_),
    .Z(_193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _475_ (.I0(net40),
    .I1(net10),
    .S(_076_),
    .Z(_194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _476_ (.A1(net10),
    .A2(_146_),
    .B1(_194_),
    .B2(_181_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _477_ (.A1(_275_),
    .A2(_187_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _478_ (.A1(net41),
    .A2(_118_),
    .A3(_196_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _479_ (.A1(_191_),
    .A2(_193_),
    .B1(_195_),
    .B2(_053_),
    .C(_197_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _480_ (.I0(_198_),
    .I1(net41),
    .S(_178_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _481_ (.A1(net24),
    .A2(_108_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _482_ (.I0(_199_),
    .I1(net25),
    .S(_273_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _483_ (.A1(_274_),
    .A2(_271_),
    .Z(_201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _484_ (.A1(_200_),
    .A2(_201_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _485_ (.A1(net42),
    .A2(_118_),
    .A3(_202_),
    .Z(_203_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _486_ (.I(net3),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _487_ (.I0(net41),
    .I1(net11),
    .S(_063_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _488_ (.A1(net11),
    .A2(_146_),
    .B1(_205_),
    .B2(_181_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _489_ (.A1(_204_),
    .A2(_193_),
    .B1(_206_),
    .B2(_052_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _490_ (.I0(_207_),
    .I1(net42),
    .S(_178_),
    .Z(_208_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _491_ (.A1(_203_),
    .A2(_208_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _492_ (.I(net4),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _493_ (.I0(net42),
    .I1(net12),
    .S(_076_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _494_ (.A1(net12),
    .A2(_146_),
    .B1(_210_),
    .B2(_181_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _495_ (.A1(_277_),
    .A2(_187_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _496_ (.A1(net43),
    .A2(_118_),
    .A3(_212_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _497_ (.A1(_209_),
    .A2(_193_),
    .B1(_211_),
    .B2(_053_),
    .C(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _498_ (.I0(_214_),
    .I1(net43),
    .S(_178_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _499_ (.A1(_274_),
    .A2(net23),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _500_ (.A1(_200_),
    .A2(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _501_ (.A1(net44),
    .A2(_118_),
    .A3(_216_),
    .Z(_217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _502_ (.I(net5),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _503_ (.I0(net43),
    .I1(net13),
    .S(_063_),
    .Z(_219_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _504_ (.A1(net13),
    .A2(_146_),
    .B1(_219_),
    .B2(_181_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _505_ (.A1(_218_),
    .A2(_193_),
    .B1(_220_),
    .B2(_052_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _506_ (.I0(_221_),
    .I1(net44),
    .S(_178_),
    .Z(_222_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _507_ (.A1(_217_),
    .A2(_222_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _508_ (.I(net6),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _509_ (.I0(net44),
    .I1(net14),
    .S(_063_),
    .Z(_224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _510_ (.A1(net14),
    .A2(_146_),
    .B1(_224_),
    .B2(_181_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _511_ (.I(_275_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _512_ (.A1(_226_),
    .A2(_187_),
    .B(_118_),
    .C(net45),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _513_ (.A1(_223_),
    .A2(_193_),
    .B1(_225_),
    .B2(_053_),
    .C(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _514_ (.I0(_228_),
    .I1(net45),
    .S(_178_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _515_ (.I(net7),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _516_ (.I0(net45),
    .I1(net15),
    .S(_076_),
    .Z(_230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _517_ (.A1(net15),
    .A2(_146_),
    .B1(_230_),
    .B2(_181_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _518_ (.A1(_229_),
    .A2(_193_),
    .B1(_231_),
    .B2(_053_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _519_ (.I(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _520_ (.I0(net25),
    .I1(_199_),
    .S(_273_),
    .Z(_234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _521_ (.A1(_201_),
    .A2(_234_),
    .B(_119_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _522_ (.A1(_178_),
    .A2(_235_),
    .B(net46),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _523_ (.A1(_178_),
    .A2(_233_),
    .B(_236_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _524_ (.I(net8),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _525_ (.I0(net46),
    .I1(net16),
    .S(_063_),
    .Z(_238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _526_ (.A1(net16),
    .A2(_146_),
    .B1(_238_),
    .B2(_181_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _527_ (.I(_277_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _528_ (.A1(_240_),
    .A2(_187_),
    .B(_118_),
    .C(net47),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _529_ (.A1(_237_),
    .A2(_193_),
    .B1(_239_),
    .B2(_053_),
    .C(_241_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _530_ (.I0(_242_),
    .I1(net47),
    .S(_178_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _531_ (.A1(_068_),
    .A2(_071_),
    .B1(_086_),
    .B2(_122_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _532_ (.I(_283_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _533_ (.A1(_061_),
    .A2(_100_),
    .A3(_244_),
    .B(_103_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _534_ (.A1(_101_),
    .A2(_068_),
    .B(_143_),
    .C(_117_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _535_ (.A1(_066_),
    .A2(_245_),
    .B(_246_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _536_ (.A1(_096_),
    .A2(_243_),
    .A3(_247_),
    .Z(_248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _537_ (.I0(_085_),
    .I1(_076_),
    .S(_248_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _538_ (.A1(_054_),
    .A2(cmd_read),
    .A3(_058_),
    .A4(_094_),
    .Z(_249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _539_ (.A1(_123_),
    .A2(cmd_read),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _540_ (.A1(_076_),
    .A2(_250_),
    .B(_180_),
    .C(_052_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _541_ (.A1(_075_),
    .A2(_076_),
    .A3(_094_),
    .Z(_252_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _542_ (.A1(_249_),
    .A2(_251_),
    .A3(_252_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _543_ (.A1(_167_),
    .A2(_248_),
    .B(_066_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _544_ (.A1(_248_),
    .A2(_253_),
    .B(_254_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _545_ (.A1(_100_),
    .A2(_173_),
    .Z(_255_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _546_ (.A1(_061_),
    .A2(_145_),
    .B(_100_),
    .C(_075_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _547_ (.A1(_255_),
    .A2(_256_),
    .B(_053_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _548_ (.A1(_251_),
    .A2(_257_),
    .Z(_258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _549_ (.I0(_258_),
    .I1(_100_),
    .S(_248_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _550_ (.A1(_058_),
    .A2(_130_),
    .A3(_250_),
    .Z(_259_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _551_ (.A1(_259_),
    .A2(_093_),
    .Z(_260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _552_ (.I0(_260_),
    .I1(_053_),
    .S(_248_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _553_ (.A1(_052_),
    .A2(_117_),
    .A3(_056_),
    .Z(_261_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _554_ (.A1(_109_),
    .A2(_261_),
    .Z(_262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _555_ (.I0(net26),
    .I1(_262_),
    .S(_042_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _556_ (.A1(_281_),
    .A2(_283_),
    .Z(_263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _557_ (.I0(net36),
    .I1(_263_),
    .S(_042_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _558_ (.I0(_282_),
    .I1(net37),
    .S(_041_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _559_ (.A1(_103_),
    .A2(_157_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _560_ (.A1(_052_),
    .A2(_281_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _561_ (.I0(_264_),
    .I1(_265_),
    .S(_056_),
    .Z(_266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _562_ (.I0(net38),
    .I1(_266_),
    .S(_042_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _563_ (.A(_267_),
    .B(_268_),
    .CO(_269_),
    .S(_270_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _564_ (.A(_271_),
    .B(_272_),
    .CO(_273_),
    .S(_274_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _565_ (.A(net23),
    .B(_272_),
    .CO(_275_),
    .S(_276_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _566_ (.A(net23),
    .B(net24),
    .CO(_277_),
    .S(_278_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _567_ (.A(_279_),
    .B(_280_),
    .CO(_281_),
    .S(_282_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _568_ (.A(_279_),
    .B(net37),
    .CO(_283_),
    .S(_284_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _569_ (.A(net36),
    .B(_280_),
    .CO(_285_),
    .S(_286_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _570_ (.A(net36),
    .B(net37),
    .CO(_287_),
    .S(_288_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _572_ (.I(net52),
    .Z(scl));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _573_ (.I(net53),
    .Z(sda));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ack_error$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \bit_counter_debug[0]$_DFFE_PN1P_  (.D(_009_),
    .SETN(net18),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \bit_counter_debug[1]$_DFFE_PN1P_  (.D(_010_),
    .SETN(net18),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \bit_counter_debug[2]$_DFFE_PN1P_  (.D(_011_),
    .SETN(net18),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \busy$_DFFE_PN0N_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cmd_read$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(cmd_read));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cmd_write$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(cmd_write));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[0]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[1]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[2]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[3]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[4]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[5]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[6]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[7]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net34));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \divider_counter[0]$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\divider_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \divider_counter[1]$_DFF_PN0_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\divider_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \divider_counter[2]$_DFF_PN1_  (.D(_002_),
    .SETN(net18),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\divider_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \divider_counter[3]$_DFF_PN1_  (.D(_003_),
    .SETN(net18),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\divider_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \divider_counter[4]$_DFF_PN1_  (.D(_004_),
    .SETN(net18),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \divider_counter[5]$_DFF_PN1_  (.D(_005_),
    .SETN(net18),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\divider_counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \divider_counter[6]$_DFF_PN1_  (.D(_006_),
    .SETN(net18),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\divider_counter[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \done$_DFF_PN0_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net35));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \phase[0]$_DFFE_PN0N_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net36));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \phase[1]$_DFFE_PN0N_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \scl_internal$_DFFE_PN1N_  (.D(_025_),
    .SETN(net18),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net38));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \sda_internal$_DFFE_PN1P_  (.D(_026_),
    .SETN(net18),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net39));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[0]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net40));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[1]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[2]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[3]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[4]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net44));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[5]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[6]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shift_reg_debug[7]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[0]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[2]$_DFFE_PN0P_  (.D(_037_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[3]$_DFFE_PN0P_  (.D(_038_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 hold1 (.I(net18),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_77 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_78 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_79 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_80 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_81 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_82 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_83 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_84 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_90 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(addr[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(addr[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(addr[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(addr[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(addr[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(addr[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(addr[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(data_in[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(data_in[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(data_in[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(data_in[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(data_in[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(data_in[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(data_in[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(data_in[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(read),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input17 (.I(net54),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input18 (.I(start),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input19 (.I(stop),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(write),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(ack_error));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(bit_counter_debug[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(bit_counter_debug[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(bit_counter_debug[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net26),
    .Z(busy));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output26 (.I(net27),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net28),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output28 (.I(net29),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output29 (.I(net30),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output30 (.I(net31),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output31 (.I(net32),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output32 (.I(net33),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output33 (.I(net34),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output34 (.I(net35),
    .Z(done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output35 (.I(net36),
    .Z(phase[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output36 (.I(net37),
    .Z(phase[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net38),
    .Z(scl_internal_debug));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net39),
    .Z(sda_internal_debug));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net40),
    .Z(shift_reg_debug[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net41),
    .Z(shift_reg_debug[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net42),
    .Z(shift_reg_debug[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net43),
    .Z(shift_reg_debug[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net44),
    .Z(shift_reg_debug[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net45),
    .Z(shift_reg_debug[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net46),
    .Z(shift_reg_debug[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net47),
    .Z(shift_reg_debug[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net48),
    .Z(state[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net49),
    .Z(state[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net50),
    .Z(state[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net51),
    .Z(state[3]));
 gf180mcu_fd_sc_mcu9t5v0__tiel _572__51 (.ZN(net52));
 gf180mcu_fd_sc_mcu9t5v0__tiel _573__52 (.ZN(net53));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload1 (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload2 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_15 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_332 ();
endmodule
