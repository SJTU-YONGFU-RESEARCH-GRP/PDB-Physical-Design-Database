module bidirectional_shift_register (clk,
    direction,
    enable,
    load_en,
    rst_n,
    serial_in,
    shift_en,
    parallel_in,
    parallel_out);
 input clk;
 input direction;
 input enable;
 input load_en;
 input rst_n;
 input serial_in;
 input shift_en;
 input [7:0] parallel_in;
 output [7:0] parallel_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net21;

 sky130_fd_sc_hd__buf_6 _36_ (.A(load_en),
    .X(_08_));
 sky130_fd_sc_hd__o21ai_4 _37_ (.A1(net12),
    .A2(_08_),
    .B1(net2),
    .Y(_09_));
 sky130_fd_sc_hd__buf_6 _38_ (.A(_09_),
    .X(_10_));
 sky130_fd_sc_hd__buf_6 _39_ (.A(direction),
    .X(_11_));
 sky130_fd_sc_hd__mux2_1 _40_ (.A0(net14),
    .A1(net11),
    .S(_11_),
    .X(_12_));
 sky130_fd_sc_hd__mux2i_1 _41_ (.A0(_12_),
    .A1(net3),
    .S(_08_),
    .Y(_13_));
 sky130_fd_sc_hd__nand2_1 _42_ (.A(net13),
    .B(_10_),
    .Y(_14_));
 sky130_fd_sc_hd__o21ai_0 _43_ (.A1(_10_),
    .A2(_13_),
    .B1(_14_),
    .Y(_00_));
 sky130_fd_sc_hd__mux2_1 _44_ (.A0(net15),
    .A1(net13),
    .S(_11_),
    .X(_15_));
 sky130_fd_sc_hd__mux2i_1 _45_ (.A0(_15_),
    .A1(net4),
    .S(_08_),
    .Y(_16_));
 sky130_fd_sc_hd__nand2_1 _46_ (.A(net14),
    .B(_10_),
    .Y(_17_));
 sky130_fd_sc_hd__o21ai_0 _47_ (.A1(_10_),
    .A2(_16_),
    .B1(_17_),
    .Y(_01_));
 sky130_fd_sc_hd__mux2_1 _48_ (.A0(net16),
    .A1(net14),
    .S(_11_),
    .X(_18_));
 sky130_fd_sc_hd__mux2i_1 _49_ (.A0(_18_),
    .A1(net5),
    .S(_08_),
    .Y(_19_));
 sky130_fd_sc_hd__nand2_1 _50_ (.A(net15),
    .B(_10_),
    .Y(_20_));
 sky130_fd_sc_hd__o21ai_0 _51_ (.A1(_09_),
    .A2(_19_),
    .B1(_20_),
    .Y(_02_));
 sky130_fd_sc_hd__mux2_1 _52_ (.A0(net17),
    .A1(net15),
    .S(_11_),
    .X(_21_));
 sky130_fd_sc_hd__mux2i_1 _53_ (.A0(_21_),
    .A1(net6),
    .S(_08_),
    .Y(_22_));
 sky130_fd_sc_hd__nand2_1 _54_ (.A(net16),
    .B(_10_),
    .Y(_23_));
 sky130_fd_sc_hd__o21ai_0 _55_ (.A1(_09_),
    .A2(_22_),
    .B1(_23_),
    .Y(_03_));
 sky130_fd_sc_hd__mux2_1 _56_ (.A0(net18),
    .A1(net16),
    .S(_11_),
    .X(_24_));
 sky130_fd_sc_hd__mux2i_1 _57_ (.A0(_24_),
    .A1(net7),
    .S(_08_),
    .Y(_25_));
 sky130_fd_sc_hd__nand2_1 _58_ (.A(net17),
    .B(_10_),
    .Y(_26_));
 sky130_fd_sc_hd__o21ai_0 _59_ (.A1(_09_),
    .A2(_25_),
    .B1(_26_),
    .Y(_04_));
 sky130_fd_sc_hd__mux2_1 _60_ (.A0(net19),
    .A1(net17),
    .S(_11_),
    .X(_27_));
 sky130_fd_sc_hd__mux2i_1 _61_ (.A0(_27_),
    .A1(net8),
    .S(_08_),
    .Y(_28_));
 sky130_fd_sc_hd__nand2_1 _62_ (.A(net18),
    .B(_10_),
    .Y(_29_));
 sky130_fd_sc_hd__o21ai_0 _63_ (.A1(_09_),
    .A2(_28_),
    .B1(_29_),
    .Y(_05_));
 sky130_fd_sc_hd__mux2_1 _64_ (.A0(net20),
    .A1(net18),
    .S(_11_),
    .X(_30_));
 sky130_fd_sc_hd__mux2i_1 _65_ (.A0(_30_),
    .A1(net9),
    .S(_08_),
    .Y(_31_));
 sky130_fd_sc_hd__nand2_1 _66_ (.A(net19),
    .B(_10_),
    .Y(_32_));
 sky130_fd_sc_hd__o21ai_0 _67_ (.A1(_09_),
    .A2(_31_),
    .B1(_32_),
    .Y(_06_));
 sky130_fd_sc_hd__mux2_1 _68_ (.A0(net11),
    .A1(net19),
    .S(_11_),
    .X(_33_));
 sky130_fd_sc_hd__mux2i_1 _69_ (.A0(_33_),
    .A1(net10),
    .S(_08_),
    .Y(_34_));
 sky130_fd_sc_hd__nand2_1 _70_ (.A(net20),
    .B(_10_),
    .Y(_35_));
 sky130_fd_sc_hd__o21ai_0 _71_ (.A1(_09_),
    .A2(_34_),
    .B1(_35_),
    .Y(_07_));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[0]$_DFFE_PN0P_  (.D(_00_),
    .Q(net13),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[1]$_DFFE_PN0P_  (.D(_01_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[2]$_DFFE_PN0P_  (.D(_02_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[3]$_DFFE_PN0P_  (.D(_03_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[4]$_DFFE_PN0P_  (.D(_04_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[5]$_DFFE_PN0P_  (.D(_05_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[6]$_DFFE_PN0P_  (.D(_06_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[7]$_DFFE_PN0P_  (.D(_07_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__buf_2 hold1 (.A(net21),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_66 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(enable),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(parallel_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(parallel_in[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(parallel_in[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(parallel_in[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(parallel_in[4]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(parallel_in[5]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(parallel_in[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(parallel_in[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(serial_in),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(shift_en),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(parallel_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(parallel_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(parallel_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(parallel_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(parallel_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(parallel_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(parallel_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(parallel_out[7]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net21));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_155 ();
endmodule
