module parameterized_uart_rx (clk,
    data_valid,
    frame_error,
    parity_error,
    rst_n,
    rx,
    data_out);
 input clk;
 output data_valid;
 output frame_error;
 output parity_error;
 input rst_n;
 input rx;
 output [7:0] data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire clknet_0_clk;
 wire \bit_index[0] ;
 wire \bit_index[1] ;
 wire \bit_index[2] ;
 wire \clk_counter[0] ;
 wire \clk_counter[10] ;
 wire \clk_counter[11] ;
 wire \clk_counter[12] ;
 wire \clk_counter[13] ;
 wire \clk_counter[14] ;
 wire \clk_counter[15] ;
 wire \clk_counter[16] ;
 wire \clk_counter[17] ;
 wire \clk_counter[18] ;
 wire \clk_counter[19] ;
 wire \clk_counter[1] ;
 wire \clk_counter[20] ;
 wire \clk_counter[21] ;
 wire \clk_counter[22] ;
 wire \clk_counter[23] ;
 wire \clk_counter[24] ;
 wire \clk_counter[25] ;
 wire \clk_counter[26] ;
 wire \clk_counter[27] ;
 wire \clk_counter[28] ;
 wire \clk_counter[29] ;
 wire \clk_counter[2] ;
 wire \clk_counter[30] ;
 wire \clk_counter[31] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \clk_counter[6] ;
 wire \clk_counter[7] ;
 wire \clk_counter[8] ;
 wire \clk_counter[9] ;
 wire \rx_data[0] ;
 wire \rx_data[1] ;
 wire \rx_data[2] ;
 wire \rx_data[3] ;
 wire \rx_data[4] ;
 wire \rx_data[5] ;
 wire \rx_data[6] ;
 wire \rx_data[7] ;
 wire rx_meta;
 wire rx_sync;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 BUF_X2 _392_ (.A(rst_n),
    .Z(_064_));
 INV_X2 _393_ (.A(_064_),
    .ZN(_065_));
 CLKBUF_X3 _394_ (.A(_065_),
    .Z(_066_));
 CLKBUF_X3 _395_ (.A(\state[2] ),
    .Z(_067_));
 INV_X1 _396_ (.A(_067_),
    .ZN(_068_));
 NOR2_X1 _397_ (.A1(\clk_counter[17] ),
    .A2(\clk_counter[16] ),
    .ZN(_069_));
 BUF_X2 _398_ (.A(\clk_counter[13] ),
    .Z(_070_));
 CLKBUF_X3 _399_ (.A(\clk_counter[12] ),
    .Z(_071_));
 BUF_X4 _400_ (.A(\clk_counter[14] ),
    .Z(_072_));
 NOR4_X4 _401_ (.A1(_070_),
    .A2(_071_),
    .A3(\clk_counter[15] ),
    .A4(_072_),
    .ZN(_073_));
 BUF_X2 _402_ (.A(\clk_counter[11] ),
    .Z(_074_));
 BUF_X4 _403_ (.A(\clk_counter[10] ),
    .Z(_075_));
 BUF_X4 _404_ (.A(\clk_counter[19] ),
    .Z(_076_));
 NOR4_X2 _405_ (.A1(\clk_counter[8] ),
    .A2(_074_),
    .A3(_075_),
    .A4(_076_),
    .ZN(_077_));
 CLKBUF_X3 _406_ (.A(\clk_counter[7] ),
    .Z(_078_));
 CLKBUF_X3 _407_ (.A(\clk_counter[6] ),
    .Z(_079_));
 NOR4_X4 _408_ (.A1(_078_),
    .A2(_079_),
    .A3(\clk_counter[9] ),
    .A4(\clk_counter[30] ),
    .ZN(_080_));
 NAND4_X4 _409_ (.A1(_069_),
    .A2(_073_),
    .A3(_077_),
    .A4(_080_),
    .ZN(_081_));
 BUF_X2 _410_ (.A(\clk_counter[29] ),
    .Z(_082_));
 NOR4_X4 _411_ (.A1(\clk_counter[24] ),
    .A2(_082_),
    .A3(\clk_counter[28] ),
    .A4(\clk_counter[31] ),
    .ZN(_083_));
 BUF_X2 _412_ (.A(\clk_counter[18] ),
    .Z(_084_));
 BUF_X2 _413_ (.A(\clk_counter[25] ),
    .Z(_085_));
 NOR4_X4 _414_ (.A1(_084_),
    .A2(_085_),
    .A3(\clk_counter[27] ),
    .A4(\clk_counter[26] ),
    .ZN(_086_));
 NAND2_X2 _415_ (.A1(_083_),
    .A2(_086_),
    .ZN(_087_));
 BUF_X2 _416_ (.A(\clk_counter[21] ),
    .Z(_088_));
 BUF_X2 _417_ (.A(\clk_counter[20] ),
    .Z(_089_));
 BUF_X2 _418_ (.A(\clk_counter[22] ),
    .Z(_090_));
 OR4_X2 _419_ (.A1(_088_),
    .A2(_089_),
    .A3(\clk_counter[23] ),
    .A4(_090_),
    .ZN(_091_));
 CLKBUF_X2 _420_ (.A(\clk_counter[5] ),
    .Z(_092_));
 BUF_X2 _421_ (.A(\clk_counter[4] ),
    .Z(_093_));
 BUF_X2 _422_ (.A(\clk_counter[2] ),
    .Z(_094_));
 BUF_X2 _423_ (.A(\clk_counter[3] ),
    .Z(_095_));
 NOR2_X1 _424_ (.A1(_094_),
    .A2(_095_),
    .ZN(_096_));
 NAND4_X2 _425_ (.A1(_092_),
    .A2(_093_),
    .A3(_375_),
    .A4(_096_),
    .ZN(_097_));
 NOR4_X4 _426_ (.A1(_081_),
    .A2(_087_),
    .A3(_091_),
    .A4(_097_),
    .ZN(_098_));
 CLKBUF_X3 _427_ (.A(_098_),
    .Z(_099_));
 AOI21_X1 _428_ (.A(_068_),
    .B1(_389_),
    .B2(_099_),
    .ZN(_100_));
 BUF_X2 _429_ (.A(rx_sync),
    .Z(_101_));
 INV_X2 _430_ (.A(\state[3] ),
    .ZN(_102_));
 NOR2_X2 _431_ (.A1(_101_),
    .A2(_102_),
    .ZN(_103_));
 INV_X1 _432_ (.A(_094_),
    .ZN(_104_));
 NAND4_X4 _433_ (.A1(_104_),
    .A2(_095_),
    .A3(_377_),
    .A4(_093_),
    .ZN(_105_));
 INV_X1 _434_ (.A(_092_),
    .ZN(_106_));
 NOR4_X4 _435_ (.A1(_088_),
    .A2(_089_),
    .A3(\clk_counter[23] ),
    .A4(_090_),
    .ZN(_107_));
 NAND4_X4 _436_ (.A1(_106_),
    .A2(_083_),
    .A3(_086_),
    .A4(_107_),
    .ZN(_108_));
 NOR3_X4 _437_ (.A1(_105_),
    .A2(_081_),
    .A3(_108_),
    .ZN(_109_));
 AOI21_X1 _438_ (.A(_100_),
    .B1(_103_),
    .B2(_109_),
    .ZN(_110_));
 NOR2_X1 _439_ (.A1(_066_),
    .A2(_110_),
    .ZN(_002_));
 NAND2_X1 _440_ (.A1(_094_),
    .A2(_095_),
    .ZN(_111_));
 INV_X1 _441_ (.A(_093_),
    .ZN(_112_));
 NAND2_X1 _442_ (.A1(_112_),
    .A2(_373_),
    .ZN(_113_));
 NOR4_X4 _443_ (.A1(_081_),
    .A2(_108_),
    .A3(_111_),
    .A4(_113_),
    .ZN(_114_));
 BUF_X2 _444_ (.A(\state[0] ),
    .Z(_115_));
 AOI221_X1 _445_ (.A(_065_),
    .B1(\state[4] ),
    .B2(_114_),
    .C1(_101_),
    .C2(_115_),
    .ZN(_116_));
 INV_X1 _446_ (.A(_006_),
    .ZN(_117_));
 NAND3_X1 _447_ (.A1(\state[3] ),
    .A2(_117_),
    .A3(_109_),
    .ZN(_118_));
 NAND2_X1 _448_ (.A1(_116_),
    .A2(_118_),
    .ZN(_000_));
 BUF_X2 _449_ (.A(_064_),
    .Z(_119_));
 INV_X1 _450_ (.A(_115_),
    .ZN(_120_));
 OAI22_X1 _451_ (.A1(_120_),
    .A2(_101_),
    .B1(_102_),
    .B2(_109_),
    .ZN(_121_));
 AND2_X1 _452_ (.A1(_119_),
    .A2(_121_),
    .ZN(_003_));
 INV_X1 _453_ (.A(\state[4] ),
    .ZN(_122_));
 NOR3_X1 _454_ (.A1(_065_),
    .A2(_122_),
    .A3(_114_),
    .ZN(_123_));
 BUF_X2 _455_ (.A(\state[1] ),
    .Z(_124_));
 AND3_X1 _456_ (.A1(_064_),
    .A2(_124_),
    .A3(_099_),
    .ZN(_052_));
 OR2_X1 _457_ (.A1(_123_),
    .A2(_052_),
    .ZN(_004_));
 OR4_X2 _458_ (.A1(_081_),
    .A2(_087_),
    .A3(_091_),
    .A4(_097_),
    .ZN(_125_));
 BUF_X8 _459_ (.A(_125_),
    .Z(_126_));
 NAND2_X1 _460_ (.A1(_124_),
    .A2(_126_),
    .ZN(_127_));
 BUF_X2 _461_ (.A(_067_),
    .Z(_128_));
 NAND3_X1 _462_ (.A1(_128_),
    .A2(_389_),
    .A3(_099_),
    .ZN(_129_));
 AOI21_X1 _463_ (.A(_066_),
    .B1(_127_),
    .B2(_129_),
    .ZN(_001_));
 CLKBUF_X2 _464_ (.A(\bit_index[0] ),
    .Z(_130_));
 OR4_X1 _465_ (.A1(_068_),
    .A2(_389_),
    .A3(_130_),
    .A4(_126_),
    .ZN(_131_));
 INV_X1 _466_ (.A(_130_),
    .ZN(_132_));
 NAND2_X1 _467_ (.A1(_120_),
    .A2(_068_),
    .ZN(_133_));
 AOI22_X4 _468_ (.A1(_109_),
    .A2(_103_),
    .B1(_133_),
    .B2(_102_),
    .ZN(_134_));
 MUX2_X1 _469_ (.A(_131_),
    .B(_132_),
    .S(_134_),
    .Z(_135_));
 NAND3_X1 _470_ (.A1(_128_),
    .A2(_130_),
    .A3(_126_),
    .ZN(_136_));
 AOI21_X1 _471_ (.A(_066_),
    .B1(_135_),
    .B2(_136_),
    .ZN(_009_));
 INV_X1 _472_ (.A(_384_),
    .ZN(_137_));
 OR4_X1 _473_ (.A1(_068_),
    .A2(_389_),
    .A3(_137_),
    .A4(_126_),
    .ZN(_138_));
 INV_X1 _474_ (.A(\bit_index[1] ),
    .ZN(_139_));
 MUX2_X1 _475_ (.A(_138_),
    .B(_139_),
    .S(_134_),
    .Z(_140_));
 NAND3_X1 _476_ (.A1(_128_),
    .A2(\bit_index[1] ),
    .A3(_126_),
    .ZN(_141_));
 AOI21_X1 _477_ (.A(_066_),
    .B1(_140_),
    .B2(_141_),
    .ZN(_010_));
 NAND3_X1 _478_ (.A1(_128_),
    .A2(_390_),
    .A3(_099_),
    .ZN(_142_));
 BUF_X2 _479_ (.A(\bit_index[2] ),
    .Z(_143_));
 INV_X1 _480_ (.A(_143_),
    .ZN(_144_));
 MUX2_X1 _481_ (.A(_142_),
    .B(_144_),
    .S(_134_),
    .Z(_145_));
 NAND3_X1 _482_ (.A1(_128_),
    .A2(_143_),
    .A3(_126_),
    .ZN(_146_));
 AOI21_X1 _483_ (.A(_066_),
    .B1(_145_),
    .B2(_146_),
    .ZN(_011_));
 OR4_X2 _484_ (.A1(_067_),
    .A2(\state[3] ),
    .A3(\state[4] ),
    .A4(_124_),
    .ZN(_147_));
 NOR2_X2 _485_ (.A1(_115_),
    .A2(_147_),
    .ZN(_148_));
 BUF_X4 _486_ (.A(_148_),
    .Z(_149_));
 INV_X1 _487_ (.A(_101_),
    .ZN(_150_));
 OR2_X2 _488_ (.A1(_150_),
    .A2(_005_),
    .ZN(_151_));
 NOR4_X4 _489_ (.A1(_105_),
    .A2(_081_),
    .A3(_108_),
    .A4(_151_),
    .ZN(_152_));
 BUF_X4 _490_ (.A(_152_),
    .Z(_153_));
 OAI21_X1 _491_ (.A(\clk_counter[0] ),
    .B1(_149_),
    .B2(_153_),
    .ZN(_154_));
 INV_X1 _492_ (.A(\clk_counter[0] ),
    .ZN(_155_));
 NOR2_X1 _493_ (.A1(_067_),
    .A2(_124_),
    .ZN(_156_));
 OAI222_X2 _494_ (.A1(_102_),
    .A2(_109_),
    .B1(_099_),
    .B2(_156_),
    .C1(_114_),
    .C2(_122_),
    .ZN(_157_));
 NOR4_X4 _495_ (.A1(_067_),
    .A2(\state[3] ),
    .A3(\state[4] ),
    .A4(_124_),
    .ZN(_158_));
 NOR2_X2 _496_ (.A1(_158_),
    .A2(_153_),
    .ZN(_159_));
 NAND3_X1 _497_ (.A1(_155_),
    .A2(_157_),
    .A3(_159_),
    .ZN(_160_));
 AOI21_X1 _498_ (.A(_066_),
    .B1(_154_),
    .B2(_160_),
    .ZN(_012_));
 NAND2_X1 _499_ (.A1(_115_),
    .A2(_158_),
    .ZN(_161_));
 OAI222_X2 _500_ (.A1(_102_),
    .A2(_109_),
    .B1(_098_),
    .B2(_156_),
    .C1(_114_),
    .C2(_008_),
    .ZN(_162_));
 OR2_X1 _501_ (.A1(_158_),
    .A2(_152_),
    .ZN(_163_));
 OAI221_X2 _502_ (.A(_064_),
    .B1(_152_),
    .B2(_161_),
    .C1(_162_),
    .C2(_163_),
    .ZN(_164_));
 BUF_X4 _503_ (.A(_164_),
    .Z(_165_));
 BUF_X4 _504_ (.A(_165_),
    .Z(_166_));
 OAI21_X4 _505_ (.A(_379_),
    .B1(_147_),
    .B2(_115_),
    .ZN(_167_));
 AND4_X2 _506_ (.A1(_094_),
    .A2(_095_),
    .A3(_092_),
    .A4(_093_),
    .ZN(_168_));
 AND2_X1 _507_ (.A1(\clk_counter[9] ),
    .A2(\clk_counter[8] ),
    .ZN(_169_));
 NAND4_X4 _508_ (.A1(_078_),
    .A2(_079_),
    .A3(_168_),
    .A4(_169_),
    .ZN(_170_));
 NOR3_X1 _509_ (.A1(_153_),
    .A2(_167_),
    .A3(_170_),
    .ZN(_171_));
 XNOR2_X1 _510_ (.A(_075_),
    .B(_171_),
    .ZN(_172_));
 NOR2_X1 _511_ (.A1(_166_),
    .A2(_172_),
    .ZN(_013_));
 BUF_X4 _512_ (.A(_152_),
    .Z(_173_));
 NAND2_X4 _513_ (.A1(\clk_counter[0] ),
    .A2(\clk_counter[1] ),
    .ZN(_174_));
 AND4_X2 _514_ (.A1(_078_),
    .A2(_079_),
    .A3(_168_),
    .A4(_169_),
    .ZN(_175_));
 NAND2_X1 _515_ (.A1(_075_),
    .A2(_175_),
    .ZN(_176_));
 NOR4_X1 _516_ (.A1(_149_),
    .A2(_173_),
    .A3(_174_),
    .A4(_176_),
    .ZN(_177_));
 XNOR2_X1 _517_ (.A(_074_),
    .B(_177_),
    .ZN(_178_));
 NOR2_X1 _518_ (.A1(_166_),
    .A2(_178_),
    .ZN(_014_));
 INV_X1 _519_ (.A(_074_),
    .ZN(_179_));
 NOR4_X1 _520_ (.A1(_179_),
    .A2(_173_),
    .A3(_167_),
    .A4(_176_),
    .ZN(_180_));
 XNOR2_X1 _521_ (.A(_071_),
    .B(_180_),
    .ZN(_181_));
 NOR2_X1 _522_ (.A1(_166_),
    .A2(_181_),
    .ZN(_015_));
 NAND4_X1 _523_ (.A1(_074_),
    .A2(_075_),
    .A3(_071_),
    .A4(_175_),
    .ZN(_182_));
 NOR4_X2 _524_ (.A1(_149_),
    .A2(_173_),
    .A3(_174_),
    .A4(_182_),
    .ZN(_183_));
 XNOR2_X1 _525_ (.A(_070_),
    .B(_183_),
    .ZN(_184_));
 NOR2_X1 _526_ (.A1(_166_),
    .A2(_184_),
    .ZN(_016_));
 AND4_X2 _527_ (.A1(_074_),
    .A2(_075_),
    .A3(_070_),
    .A4(_071_),
    .ZN(_185_));
 NAND2_X2 _528_ (.A1(_175_),
    .A2(_185_),
    .ZN(_186_));
 NOR3_X1 _529_ (.A1(_153_),
    .A2(_167_),
    .A3(_186_),
    .ZN(_187_));
 XNOR2_X1 _530_ (.A(_072_),
    .B(_187_),
    .ZN(_188_));
 NOR2_X1 _531_ (.A1(_166_),
    .A2(_188_),
    .ZN(_017_));
 OR4_X2 _532_ (.A1(_105_),
    .A2(_081_),
    .A3(_108_),
    .A4(_151_),
    .ZN(_189_));
 NOR2_X2 _533_ (.A1(_148_),
    .A2(_174_),
    .ZN(_190_));
 NAND4_X2 _534_ (.A1(_074_),
    .A2(_075_),
    .A3(_070_),
    .A4(_071_),
    .ZN(_191_));
 NOR2_X1 _535_ (.A1(_170_),
    .A2(_191_),
    .ZN(_192_));
 AND4_X1 _536_ (.A1(_072_),
    .A2(_189_),
    .A3(_190_),
    .A4(_192_),
    .ZN(_193_));
 XNOR2_X1 _537_ (.A(\clk_counter[15] ),
    .B(_193_),
    .ZN(_194_));
 NOR2_X1 _538_ (.A1(_166_),
    .A2(_194_),
    .ZN(_018_));
 NAND2_X1 _539_ (.A1(\clk_counter[15] ),
    .A2(_072_),
    .ZN(_195_));
 NOR4_X2 _540_ (.A1(_153_),
    .A2(_167_),
    .A3(_186_),
    .A4(_195_),
    .ZN(_196_));
 XNOR2_X1 _541_ (.A(\clk_counter[16] ),
    .B(_196_),
    .ZN(_197_));
 NOR2_X1 _542_ (.A1(_166_),
    .A2(_197_),
    .ZN(_019_));
 NAND2_X1 _543_ (.A1(\clk_counter[17] ),
    .A2(_064_),
    .ZN(_198_));
 INV_X1 _544_ (.A(\clk_counter[16] ),
    .ZN(_199_));
 NOR3_X1 _545_ (.A1(_199_),
    .A2(_174_),
    .A3(_195_),
    .ZN(_200_));
 AOI21_X1 _546_ (.A(_198_),
    .B1(_200_),
    .B2(_192_),
    .ZN(_201_));
 NAND3_X1 _547_ (.A1(_175_),
    .A2(_185_),
    .A3(_200_),
    .ZN(_202_));
 NOR3_X1 _548_ (.A1(\clk_counter[17] ),
    .A2(_065_),
    .A3(_202_),
    .ZN(_203_));
 OAI211_X2 _549_ (.A(_159_),
    .B(_162_),
    .C1(_201_),
    .C2(_203_),
    .ZN(_204_));
 NOR2_X1 _550_ (.A1(_149_),
    .A2(_153_),
    .ZN(_205_));
 OAI21_X1 _551_ (.A(_204_),
    .B1(_198_),
    .B2(_205_),
    .ZN(_020_));
 AND4_X1 _552_ (.A1(\clk_counter[15] ),
    .A2(_072_),
    .A3(\clk_counter[17] ),
    .A4(\clk_counter[16] ),
    .ZN(_206_));
 INV_X1 _553_ (.A(_206_),
    .ZN(_207_));
 NOR4_X1 _554_ (.A1(_173_),
    .A2(_167_),
    .A3(_186_),
    .A4(_207_),
    .ZN(_208_));
 XNOR2_X1 _555_ (.A(_084_),
    .B(_208_),
    .ZN(_209_));
 NOR2_X1 _556_ (.A1(_166_),
    .A2(_209_),
    .ZN(_021_));
 NAND2_X1 _557_ (.A1(_189_),
    .A2(_190_),
    .ZN(_210_));
 NAND3_X1 _558_ (.A1(_084_),
    .A2(_192_),
    .A3(_206_),
    .ZN(_211_));
 OAI21_X1 _559_ (.A(_076_),
    .B1(_210_),
    .B2(_211_),
    .ZN(_212_));
 OR3_X1 _560_ (.A1(_076_),
    .A2(_210_),
    .A3(_211_),
    .ZN(_213_));
 AOI21_X1 _561_ (.A(_165_),
    .B1(_212_),
    .B2(_213_),
    .ZN(_022_));
 OAI21_X1 _562_ (.A(\clk_counter[1] ),
    .B1(_149_),
    .B2(_153_),
    .ZN(_214_));
 NAND3_X1 _563_ (.A1(_374_),
    .A2(_159_),
    .A3(_162_),
    .ZN(_215_));
 AOI21_X1 _564_ (.A(_066_),
    .B1(_214_),
    .B2(_215_),
    .ZN(_023_));
 NAND3_X1 _565_ (.A1(_076_),
    .A2(_084_),
    .A3(_206_),
    .ZN(_216_));
 NOR4_X4 _566_ (.A1(_167_),
    .A2(_170_),
    .A3(_191_),
    .A4(_216_),
    .ZN(_217_));
 XNOR2_X1 _567_ (.A(_089_),
    .B(_217_),
    .ZN(_218_));
 NOR2_X1 _568_ (.A1(_166_),
    .A2(_218_),
    .ZN(_024_));
 AND3_X1 _569_ (.A1(_076_),
    .A2(_084_),
    .A3(_206_),
    .ZN(_219_));
 NAND4_X1 _570_ (.A1(_089_),
    .A2(_175_),
    .A3(_185_),
    .A4(_219_),
    .ZN(_220_));
 NOR4_X1 _571_ (.A1(_149_),
    .A2(_173_),
    .A3(_174_),
    .A4(_220_),
    .ZN(_221_));
 XNOR2_X1 _572_ (.A(_088_),
    .B(_221_),
    .ZN(_222_));
 NOR2_X1 _573_ (.A1(_166_),
    .A2(_222_),
    .ZN(_025_));
 CLKBUF_X3 _574_ (.A(_164_),
    .Z(_223_));
 NAND3_X1 _575_ (.A1(_088_),
    .A2(_089_),
    .A3(_217_),
    .ZN(_224_));
 XOR2_X1 _576_ (.A(_090_),
    .B(_224_),
    .Z(_225_));
 NOR2_X1 _577_ (.A1(_223_),
    .A2(_225_),
    .ZN(_026_));
 INV_X1 _578_ (.A(_075_),
    .ZN(_226_));
 NAND3_X1 _579_ (.A1(_074_),
    .A2(_070_),
    .A3(_071_),
    .ZN(_227_));
 NOR3_X2 _580_ (.A1(_226_),
    .A2(_170_),
    .A3(_227_),
    .ZN(_228_));
 NAND4_X4 _581_ (.A1(_189_),
    .A2(_190_),
    .A3(_228_),
    .A4(_219_),
    .ZN(_229_));
 NAND3_X1 _582_ (.A1(_088_),
    .A2(_089_),
    .A3(_090_),
    .ZN(_230_));
 OAI21_X1 _583_ (.A(\clk_counter[23] ),
    .B1(_229_),
    .B2(_230_),
    .ZN(_231_));
 OR3_X1 _584_ (.A1(\clk_counter[23] ),
    .A2(_229_),
    .A3(_230_),
    .ZN(_232_));
 AOI21_X1 _585_ (.A(_165_),
    .B1(_231_),
    .B2(_232_),
    .ZN(_027_));
 AND4_X1 _586_ (.A1(_088_),
    .A2(_089_),
    .A3(\clk_counter[23] ),
    .A4(_090_),
    .ZN(_233_));
 NAND2_X1 _587_ (.A1(_217_),
    .A2(_233_),
    .ZN(_234_));
 XOR2_X1 _588_ (.A(\clk_counter[24] ),
    .B(_234_),
    .Z(_235_));
 NOR2_X1 _589_ (.A1(_223_),
    .A2(_235_),
    .ZN(_028_));
 AND2_X1 _590_ (.A1(\clk_counter[24] ),
    .A2(_233_),
    .ZN(_236_));
 NAND4_X1 _591_ (.A1(_175_),
    .A2(_185_),
    .A3(_219_),
    .A4(_236_),
    .ZN(_237_));
 NOR4_X2 _592_ (.A1(_149_),
    .A2(_173_),
    .A3(_174_),
    .A4(_237_),
    .ZN(_238_));
 XNOR2_X1 _593_ (.A(_085_),
    .B(_238_),
    .ZN(_239_));
 NOR2_X1 _594_ (.A1(_223_),
    .A2(_239_),
    .ZN(_029_));
 NAND3_X1 _595_ (.A1(_085_),
    .A2(_217_),
    .A3(_236_),
    .ZN(_240_));
 XOR2_X1 _596_ (.A(\clk_counter[26] ),
    .B(_240_),
    .Z(_241_));
 NOR2_X1 _597_ (.A1(_223_),
    .A2(_241_),
    .ZN(_030_));
 NAND4_X2 _598_ (.A1(_085_),
    .A2(\clk_counter[24] ),
    .A3(\clk_counter[26] ),
    .A4(_233_),
    .ZN(_242_));
 OAI21_X1 _599_ (.A(\clk_counter[27] ),
    .B1(_229_),
    .B2(_242_),
    .ZN(_243_));
 OR3_X1 _600_ (.A1(\clk_counter[27] ),
    .A2(_229_),
    .A3(_242_),
    .ZN(_244_));
 AOI21_X1 _601_ (.A(_165_),
    .B1(_243_),
    .B2(_244_),
    .ZN(_031_));
 INV_X1 _602_ (.A(\clk_counter[28] ),
    .ZN(_245_));
 INV_X1 _603_ (.A(\clk_counter[27] ),
    .ZN(_246_));
 NOR2_X1 _604_ (.A1(_246_),
    .A2(_242_),
    .ZN(_247_));
 NAND2_X1 _605_ (.A1(_217_),
    .A2(_247_),
    .ZN(_248_));
 XNOR2_X1 _606_ (.A(_245_),
    .B(_248_),
    .ZN(_249_));
 NOR2_X1 _607_ (.A1(_223_),
    .A2(_249_),
    .ZN(_032_));
 NAND2_X1 _608_ (.A1(\clk_counter[28] ),
    .A2(_247_),
    .ZN(_250_));
 OAI21_X1 _609_ (.A(_082_),
    .B1(_229_),
    .B2(_250_),
    .ZN(_251_));
 OR3_X1 _610_ (.A1(_082_),
    .A2(_229_),
    .A3(_250_),
    .ZN(_252_));
 AOI21_X1 _611_ (.A(_165_),
    .B1(_251_),
    .B2(_252_),
    .ZN(_033_));
 NOR2_X1 _612_ (.A1(_153_),
    .A2(_167_),
    .ZN(_253_));
 XNOR2_X1 _613_ (.A(_094_),
    .B(_253_),
    .ZN(_254_));
 NOR2_X1 _614_ (.A1(_223_),
    .A2(_254_),
    .ZN(_034_));
 NOR3_X1 _615_ (.A1(_246_),
    .A2(_245_),
    .A3(_242_),
    .ZN(_255_));
 NAND3_X1 _616_ (.A1(_082_),
    .A2(_217_),
    .A3(_255_),
    .ZN(_256_));
 XOR2_X1 _617_ (.A(\clk_counter[30] ),
    .B(_256_),
    .Z(_257_));
 NOR2_X1 _618_ (.A1(_223_),
    .A2(_257_),
    .ZN(_035_));
 NAND3_X1 _619_ (.A1(_082_),
    .A2(\clk_counter[30] ),
    .A3(_255_),
    .ZN(_258_));
 OAI21_X1 _620_ (.A(\clk_counter[31] ),
    .B1(_229_),
    .B2(_258_),
    .ZN(_259_));
 OR3_X1 _621_ (.A1(\clk_counter[31] ),
    .A2(_229_),
    .A3(_258_),
    .ZN(_260_));
 AOI21_X1 _622_ (.A(_165_),
    .B1(_259_),
    .B2(_260_),
    .ZN(_036_));
 NOR4_X2 _623_ (.A1(_104_),
    .A2(_148_),
    .A3(_152_),
    .A4(_174_),
    .ZN(_261_));
 XNOR2_X1 _624_ (.A(_095_),
    .B(_261_),
    .ZN(_262_));
 NOR2_X1 _625_ (.A1(_223_),
    .A2(_262_),
    .ZN(_037_));
 NOR3_X1 _626_ (.A1(_111_),
    .A2(_153_),
    .A3(_167_),
    .ZN(_263_));
 XNOR2_X1 _627_ (.A(_093_),
    .B(_263_),
    .ZN(_264_));
 NOR2_X1 _628_ (.A1(_223_),
    .A2(_264_),
    .ZN(_038_));
 NAND3_X1 _629_ (.A1(_094_),
    .A2(_095_),
    .A3(_093_),
    .ZN(_265_));
 NOR4_X1 _630_ (.A1(_149_),
    .A2(_173_),
    .A3(_174_),
    .A4(_265_),
    .ZN(_266_));
 XNOR2_X1 _631_ (.A(_092_),
    .B(_266_),
    .ZN(_267_));
 NOR2_X1 _632_ (.A1(_223_),
    .A2(_267_),
    .ZN(_039_));
 INV_X1 _633_ (.A(_168_),
    .ZN(_268_));
 NOR3_X1 _634_ (.A1(_153_),
    .A2(_167_),
    .A3(_268_),
    .ZN(_269_));
 XNOR2_X1 _635_ (.A(_079_),
    .B(_269_),
    .ZN(_270_));
 NOR2_X1 _636_ (.A1(_165_),
    .A2(_270_),
    .ZN(_040_));
 NAND2_X1 _637_ (.A1(_079_),
    .A2(_168_),
    .ZN(_271_));
 NOR4_X1 _638_ (.A1(_149_),
    .A2(_173_),
    .A3(_271_),
    .A4(_174_),
    .ZN(_272_));
 XNOR2_X1 _639_ (.A(_078_),
    .B(_272_),
    .ZN(_273_));
 NOR2_X1 _640_ (.A1(_165_),
    .A2(_273_),
    .ZN(_041_));
 INV_X1 _641_ (.A(_078_),
    .ZN(_274_));
 NOR4_X1 _642_ (.A1(_274_),
    .A2(_173_),
    .A3(_167_),
    .A4(_271_),
    .ZN(_275_));
 XNOR2_X1 _643_ (.A(\clk_counter[8] ),
    .B(_275_),
    .ZN(_276_));
 NOR2_X1 _644_ (.A1(_165_),
    .A2(_276_),
    .ZN(_042_));
 NAND4_X1 _645_ (.A1(_078_),
    .A2(_079_),
    .A3(\clk_counter[8] ),
    .A4(_168_),
    .ZN(_277_));
 NOR4_X1 _646_ (.A1(_149_),
    .A2(_173_),
    .A3(_277_),
    .A4(_174_),
    .ZN(_278_));
 XNOR2_X1 _647_ (.A(\clk_counter[9] ),
    .B(_278_),
    .ZN(_279_));
 NOR2_X1 _648_ (.A1(_165_),
    .A2(_279_),
    .ZN(_043_));
 NOR2_X4 _649_ (.A1(_007_),
    .A2(_126_),
    .ZN(_280_));
 MUX2_X1 _650_ (.A(net2),
    .B(\rx_data[0] ),
    .S(_280_),
    .Z(_281_));
 AND2_X1 _651_ (.A1(_119_),
    .A2(_281_),
    .ZN(_044_));
 MUX2_X1 _652_ (.A(net3),
    .B(\rx_data[1] ),
    .S(_280_),
    .Z(_282_));
 AND2_X1 _653_ (.A1(_119_),
    .A2(_282_),
    .ZN(_045_));
 MUX2_X1 _654_ (.A(net4),
    .B(\rx_data[2] ),
    .S(_280_),
    .Z(_283_));
 AND2_X1 _655_ (.A1(_119_),
    .A2(_283_),
    .ZN(_046_));
 MUX2_X1 _656_ (.A(net5),
    .B(\rx_data[3] ),
    .S(_280_),
    .Z(_284_));
 AND2_X1 _657_ (.A1(_119_),
    .A2(_284_),
    .ZN(_047_));
 MUX2_X1 _658_ (.A(net6),
    .B(\rx_data[4] ),
    .S(_280_),
    .Z(_285_));
 AND2_X1 _659_ (.A1(_119_),
    .A2(_285_),
    .ZN(_048_));
 MUX2_X1 _660_ (.A(net7),
    .B(\rx_data[5] ),
    .S(_280_),
    .Z(_286_));
 AND2_X1 _661_ (.A1(_119_),
    .A2(_286_),
    .ZN(_049_));
 MUX2_X1 _662_ (.A(net8),
    .B(\rx_data[6] ),
    .S(_280_),
    .Z(_287_));
 AND2_X1 _663_ (.A1(_119_),
    .A2(_287_),
    .ZN(_050_));
 MUX2_X1 _664_ (.A(net9),
    .B(\rx_data[7] ),
    .S(_280_),
    .Z(_288_));
 AND2_X1 _665_ (.A1(_119_),
    .A2(_288_),
    .ZN(_051_));
 OAI21_X1 _666_ (.A(net11),
    .B1(_124_),
    .B2(_120_),
    .ZN(_289_));
 NAND3_X1 _667_ (.A1(_150_),
    .A2(_124_),
    .A3(_099_),
    .ZN(_290_));
 AOI21_X1 _668_ (.A(_066_),
    .B1(_289_),
    .B2(_290_),
    .ZN(_053_));
 NOR4_X1 _669_ (.A1(_130_),
    .A2(\bit_index[1] ),
    .A3(_143_),
    .A4(_384_),
    .ZN(_291_));
 XOR2_X2 _670_ (.A(_143_),
    .B(_383_),
    .Z(_292_));
 NAND4_X1 _671_ (.A1(_128_),
    .A2(_099_),
    .A3(_291_),
    .A4(_292_),
    .ZN(_293_));
 MUX2_X1 _672_ (.A(_101_),
    .B(\rx_data[0] ),
    .S(_293_),
    .Z(_294_));
 AND2_X1 _673_ (.A1(_119_),
    .A2(_294_),
    .ZN(_054_));
 INV_X1 _674_ (.A(_385_),
    .ZN(_295_));
 XNOR2_X2 _675_ (.A(_143_),
    .B(_383_),
    .ZN(_296_));
 NAND3_X2 _676_ (.A1(_067_),
    .A2(_098_),
    .A3(_296_),
    .ZN(_297_));
 OAI21_X1 _677_ (.A(\rx_data[1] ),
    .B1(_295_),
    .B2(_297_),
    .ZN(_298_));
 NAND2_X1 _678_ (.A1(_101_),
    .A2(_130_),
    .ZN(_299_));
 OR3_X1 _679_ (.A1(_137_),
    .A2(_297_),
    .A3(_299_),
    .ZN(_300_));
 AOI21_X1 _680_ (.A(_066_),
    .B1(_298_),
    .B2(_300_),
    .ZN(_055_));
 NOR2_X1 _681_ (.A1(\bit_index[1] ),
    .A2(_143_),
    .ZN(_301_));
 NOR3_X1 _682_ (.A1(_130_),
    .A2(_137_),
    .A3(_301_),
    .ZN(_302_));
 NAND4_X1 _683_ (.A1(_128_),
    .A2(_098_),
    .A3(_296_),
    .A4(_302_),
    .ZN(_303_));
 MUX2_X1 _684_ (.A(_117_),
    .B(\rx_data[2] ),
    .S(_303_),
    .Z(_304_));
 AND2_X1 _685_ (.A1(_064_),
    .A2(_304_),
    .ZN(_056_));
 INV_X1 _686_ (.A(_387_),
    .ZN(_305_));
 OAI21_X1 _687_ (.A(\rx_data[3] ),
    .B1(_305_),
    .B2(_297_),
    .ZN(_306_));
 NOR2_X1 _688_ (.A1(_384_),
    .A2(_299_),
    .ZN(_307_));
 NAND4_X1 _689_ (.A1(_128_),
    .A2(_099_),
    .A3(_296_),
    .A4(_307_),
    .ZN(_308_));
 AOI21_X1 _690_ (.A(_066_),
    .B1(_306_),
    .B2(_308_),
    .ZN(_057_));
 OR3_X1 _691_ (.A1(_130_),
    .A2(_384_),
    .A3(_301_),
    .ZN(_309_));
 OAI21_X1 _692_ (.A(\rx_data[4] ),
    .B1(_297_),
    .B2(_309_),
    .ZN(_310_));
 OR3_X1 _693_ (.A1(_006_),
    .A2(_297_),
    .A3(_309_),
    .ZN(_311_));
 AOI21_X1 _694_ (.A(_065_),
    .B1(_310_),
    .B2(_311_),
    .ZN(_058_));
 NAND3_X1 _695_ (.A1(_128_),
    .A2(_099_),
    .A3(_292_),
    .ZN(_312_));
 OAI21_X1 _696_ (.A(\rx_data[5] ),
    .B1(_295_),
    .B2(_312_),
    .ZN(_313_));
 OR3_X1 _697_ (.A1(_137_),
    .A2(_312_),
    .A3(_299_),
    .ZN(_314_));
 AOI21_X1 _698_ (.A(_065_),
    .B1(_313_),
    .B2(_314_),
    .ZN(_059_));
 NAND4_X1 _699_ (.A1(_067_),
    .A2(_098_),
    .A3(_292_),
    .A4(_302_),
    .ZN(_315_));
 MUX2_X1 _700_ (.A(_117_),
    .B(\rx_data[6] ),
    .S(_315_),
    .Z(_316_));
 AND2_X1 _701_ (.A1(_064_),
    .A2(_316_),
    .ZN(_060_));
 OAI21_X1 _702_ (.A(\rx_data[7] ),
    .B1(_305_),
    .B2(_312_),
    .ZN(_317_));
 NAND4_X1 _703_ (.A1(_128_),
    .A2(_099_),
    .A3(_292_),
    .A4(_307_),
    .ZN(_318_));
 AOI21_X1 _704_ (.A(_065_),
    .B1(_317_),
    .B2(_318_),
    .ZN(_061_));
 OR2_X1 _705_ (.A1(_065_),
    .A2(net1),
    .ZN(_062_));
 OR2_X1 _706_ (.A1(_065_),
    .A2(rx_meta),
    .ZN(_063_));
 HA_X1 _707_ (.A(_371_),
    .B(_372_),
    .CO(_373_),
    .S(_374_));
 HA_X1 _708_ (.A(_371_),
    .B(\clk_counter[1] ),
    .CO(_375_),
    .S(_376_));
 HA_X1 _709_ (.A(\clk_counter[0] ),
    .B(_372_),
    .CO(_377_),
    .S(_378_));
 HA_X1 _710_ (.A(\clk_counter[0] ),
    .B(\clk_counter[1] ),
    .CO(_379_),
    .S(_380_));
 HA_X1 _711_ (.A(_381_),
    .B(_382_),
    .CO(_383_),
    .S(_384_));
 HA_X1 _712_ (.A(\bit_index[0] ),
    .B(_382_),
    .CO(_385_),
    .S(_386_));
 HA_X1 _713_ (.A(\bit_index[0] ),
    .B(\bit_index[1] ),
    .CO(_387_),
    .S(_388_));
 HA_X1 _714_ (.A(\bit_index[2] ),
    .B(_387_),
    .CO(_389_),
    .S(_390_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X1 _716_ (.A(net12),
    .Z(parity_error));
 DFF_X1 \bit_index[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\bit_index[0] ),
    .QN(_381_));
 DFF_X2 \bit_index[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\bit_index[1] ),
    .QN(_382_));
 DFF_X1 \bit_index[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\bit_index[2] ),
    .QN(_368_));
 DFF_X2 \clk_counter[0]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[0] ),
    .QN(_371_));
 DFF_X1 \clk_counter[10]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[10] ),
    .QN(_367_));
 DFF_X1 \clk_counter[11]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[11] ),
    .QN(_366_));
 DFF_X1 \clk_counter[12]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[12] ),
    .QN(_365_));
 DFF_X1 \clk_counter[13]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[13] ),
    .QN(_364_));
 DFF_X1 \clk_counter[14]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[14] ),
    .QN(_363_));
 DFF_X2 \clk_counter[15]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[15] ),
    .QN(_362_));
 DFF_X1 \clk_counter[16]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[16] ),
    .QN(_361_));
 DFF_X1 \clk_counter[17]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[17] ),
    .QN(_360_));
 DFF_X1 \clk_counter[18]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[18] ),
    .QN(_359_));
 DFF_X1 \clk_counter[19]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[19] ),
    .QN(_358_));
 DFF_X2 \clk_counter[1]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[1] ),
    .QN(_372_));
 DFF_X1 \clk_counter[20]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[20] ),
    .QN(_357_));
 DFF_X1 \clk_counter[21]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[21] ),
    .QN(_356_));
 DFF_X1 \clk_counter[22]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[22] ),
    .QN(_355_));
 DFF_X2 \clk_counter[23]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[23] ),
    .QN(_354_));
 DFF_X2 \clk_counter[24]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[24] ),
    .QN(_353_));
 DFF_X1 \clk_counter[25]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\clk_counter[25] ),
    .QN(_352_));
 DFF_X2 \clk_counter[26]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[26] ),
    .QN(_351_));
 DFF_X2 \clk_counter[27]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[27] ),
    .QN(_350_));
 DFF_X2 \clk_counter[28]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\clk_counter[28] ),
    .QN(_349_));
 DFF_X1 \clk_counter[29]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[29] ),
    .QN(_348_));
 DFF_X1 \clk_counter[2]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[2] ),
    .QN(_347_));
 DFF_X2 \clk_counter[30]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[30] ),
    .QN(_346_));
 DFF_X2 \clk_counter[31]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[31] ),
    .QN(_345_));
 DFF_X1 \clk_counter[3]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[3] ),
    .QN(_344_));
 DFF_X1 \clk_counter[4]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[4] ),
    .QN(_343_));
 DFF_X1 \clk_counter[5]$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[5] ),
    .QN(_342_));
 DFF_X1 \clk_counter[6]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[6] ),
    .QN(_341_));
 DFF_X1 \clk_counter[7]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[7] ),
    .QN(_340_));
 DFF_X2 \clk_counter[8]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[8] ),
    .QN(_339_));
 DFF_X2 \clk_counter[9]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[9] ),
    .QN(_338_));
 DFF_X1 \data_out[0]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net2),
    .QN(_337_));
 DFF_X1 \data_out[1]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net3),
    .QN(_336_));
 DFF_X1 \data_out[2]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net4),
    .QN(_335_));
 DFF_X1 \data_out[3]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net5),
    .QN(_334_));
 DFF_X1 \data_out[4]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net6),
    .QN(_333_));
 DFF_X1 \data_out[5]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net7),
    .QN(_332_));
 DFF_X1 \data_out[6]$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net8),
    .QN(_331_));
 DFF_X1 \data_out[7]$_SDFFE_PN0P_  (.D(_051_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net9),
    .QN(_330_));
 DFF_X1 \data_valid$_SDFF_PN0_  (.D(_052_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net10),
    .QN(_329_));
 DFF_X1 \frame_error$_SDFFE_PN0P_  (.D(_053_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net11),
    .QN(_328_));
 DFF_X1 \rx_data[0]$_SDFFE_PN0P_  (.D(_054_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\rx_data[0] ),
    .QN(_327_));
 DFF_X1 \rx_data[1]$_SDFFE_PN0P_  (.D(_055_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\rx_data[1] ),
    .QN(_326_));
 DFF_X1 \rx_data[2]$_SDFFE_PN0P_  (.D(_056_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\rx_data[2] ),
    .QN(_325_));
 DFF_X1 \rx_data[3]$_SDFFE_PN0P_  (.D(_057_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\rx_data[3] ),
    .QN(_324_));
 DFF_X1 \rx_data[4]$_SDFFE_PN0P_  (.D(_058_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\rx_data[4] ),
    .QN(_323_));
 DFF_X1 \rx_data[5]$_SDFFE_PN0P_  (.D(_059_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\rx_data[5] ),
    .QN(_322_));
 DFF_X1 \rx_data[6]$_SDFFE_PN0P_  (.D(_060_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\rx_data[6] ),
    .QN(_321_));
 DFF_X1 \rx_data[7]$_SDFFE_PN0P_  (.D(_061_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\rx_data[7] ),
    .QN(_320_));
 DFF_X1 \rx_meta$_SDFF_PN1_  (.D(_062_),
    .CK(clknet_3_1__leaf_clk),
    .Q(rx_meta),
    .QN(_319_));
 DFF_X1 \rx_sync$_SDFF_PN1_  (.D(_063_),
    .CK(clknet_3_4__leaf_clk),
    .Q(rx_sync),
    .QN(_006_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_000_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\state[0] ),
    .QN(_369_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_001_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\state[1] ),
    .QN(_007_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\state[2] ),
    .QN(_370_));
 DFF_X2 \state[3]$_DFF_P_  (.D(_003_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\state[3] ),
    .QN(_005_));
 DFF_X2 \state[4]$_DFF_P_  (.D(_004_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\state[4] ),
    .QN(_008_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_73 ();
 BUF_X1 input1 (.A(rx),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(data_out[0]));
 BUF_X1 output3 (.A(net3),
    .Z(data_out[1]));
 BUF_X1 output4 (.A(net4),
    .Z(data_out[2]));
 BUF_X1 output5 (.A(net5),
    .Z(data_out[3]));
 BUF_X1 output6 (.A(net6),
    .Z(data_out[4]));
 BUF_X1 output7 (.A(net7),
    .Z(data_out[5]));
 BUF_X1 output8 (.A(net8),
    .Z(data_out[6]));
 BUF_X1 output9 (.A(net9),
    .Z(data_out[7]));
 BUF_X1 output10 (.A(net10),
    .Z(data_valid));
 BUF_X1 output11 (.A(net11),
    .Z(frame_error));
 LOGIC0_X1 _716__12 (.Z(net12));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_3_1__leaf_clk));
 INV_X1 clkload2 (.A(clknet_3_2__leaf_clk));
 INV_X4 clkload3 (.A(clknet_3_3__leaf_clk));
 INV_X1 clkload4 (.A(clknet_3_4__leaf_clk));
 INV_X1 clkload5 (.A(clknet_3_6__leaf_clk));
 INV_X4 clkload6 (.A(clknet_3_7__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_81 ();
 FILLCELL_X2 FILLER_0_85 ();
 FILLCELL_X16 FILLER_0_90 ();
 FILLCELL_X1 FILLER_0_106 ();
 FILLCELL_X8 FILLER_0_110 ();
 FILLCELL_X2 FILLER_0_118 ();
 FILLCELL_X1 FILLER_0_120 ();
 FILLCELL_X1 FILLER_0_125 ();
 FILLCELL_X32 FILLER_0_133 ();
 FILLCELL_X32 FILLER_0_165 ();
 FILLCELL_X32 FILLER_0_197 ();
 FILLCELL_X32 FILLER_0_229 ();
 FILLCELL_X8 FILLER_0_261 ();
 FILLCELL_X4 FILLER_0_269 ();
 FILLCELL_X2 FILLER_0_273 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X16 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_113 ();
 FILLCELL_X1 FILLER_1_117 ();
 FILLCELL_X32 FILLER_1_139 ();
 FILLCELL_X32 FILLER_1_171 ();
 FILLCELL_X32 FILLER_1_203 ();
 FILLCELL_X32 FILLER_1_235 ();
 FILLCELL_X8 FILLER_1_267 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_73 ();
 FILLCELL_X2 FILLER_2_77 ();
 FILLCELL_X4 FILLER_2_96 ();
 FILLCELL_X16 FILLER_2_117 ();
 FILLCELL_X1 FILLER_2_133 ();
 FILLCELL_X8 FILLER_2_151 ();
 FILLCELL_X4 FILLER_2_159 ();
 FILLCELL_X2 FILLER_2_163 ();
 FILLCELL_X1 FILLER_2_165 ();
 FILLCELL_X4 FILLER_2_185 ();
 FILLCELL_X2 FILLER_2_189 ();
 FILLCELL_X1 FILLER_2_191 ();
 FILLCELL_X4 FILLER_2_202 ();
 FILLCELL_X2 FILLER_2_206 ();
 FILLCELL_X32 FILLER_2_218 ();
 FILLCELL_X16 FILLER_2_250 ();
 FILLCELL_X8 FILLER_2_266 ();
 FILLCELL_X1 FILLER_2_274 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X4 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_37 ();
 FILLCELL_X32 FILLER_3_55 ();
 FILLCELL_X2 FILLER_3_87 ();
 FILLCELL_X8 FILLER_3_92 ();
 FILLCELL_X4 FILLER_3_100 ();
 FILLCELL_X4 FILLER_3_112 ();
 FILLCELL_X2 FILLER_3_116 ();
 FILLCELL_X16 FILLER_3_123 ();
 FILLCELL_X8 FILLER_3_139 ();
 FILLCELL_X1 FILLER_3_147 ();
 FILLCELL_X8 FILLER_3_152 ();
 FILLCELL_X2 FILLER_3_160 ();
 FILLCELL_X1 FILLER_3_162 ();
 FILLCELL_X8 FILLER_3_176 ();
 FILLCELL_X1 FILLER_3_184 ();
 FILLCELL_X16 FILLER_3_212 ();
 FILLCELL_X4 FILLER_3_230 ();
 FILLCELL_X2 FILLER_3_251 ();
 FILLCELL_X1 FILLER_3_253 ();
 FILLCELL_X16 FILLER_3_258 ();
 FILLCELL_X1 FILLER_3_274 ();
 FILLCELL_X4 FILLER_4_1 ();
 FILLCELL_X2 FILLER_4_5 ();
 FILLCELL_X4 FILLER_4_24 ();
 FILLCELL_X1 FILLER_4_28 ();
 FILLCELL_X4 FILLER_4_32 ();
 FILLCELL_X2 FILLER_4_36 ();
 FILLCELL_X1 FILLER_4_38 ();
 FILLCELL_X16 FILLER_4_48 ();
 FILLCELL_X2 FILLER_4_64 ();
 FILLCELL_X1 FILLER_4_66 ();
 FILLCELL_X2 FILLER_4_98 ();
 FILLCELL_X1 FILLER_4_104 ();
 FILLCELL_X2 FILLER_4_116 ();
 FILLCELL_X1 FILLER_4_118 ();
 FILLCELL_X4 FILLER_4_127 ();
 FILLCELL_X2 FILLER_4_135 ();
 FILLCELL_X16 FILLER_4_141 ();
 FILLCELL_X2 FILLER_4_157 ();
 FILLCELL_X1 FILLER_4_169 ();
 FILLCELL_X1 FILLER_4_179 ();
 FILLCELL_X1 FILLER_4_184 ();
 FILLCELL_X8 FILLER_4_189 ();
 FILLCELL_X4 FILLER_4_197 ();
 FILLCELL_X2 FILLER_4_201 ();
 FILLCELL_X8 FILLER_4_207 ();
 FILLCELL_X4 FILLER_4_215 ();
 FILLCELL_X16 FILLER_4_232 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_17 ();
 FILLCELL_X2 FILLER_5_21 ();
 FILLCELL_X32 FILLER_5_30 ();
 FILLCELL_X8 FILLER_5_62 ();
 FILLCELL_X4 FILLER_5_70 ();
 FILLCELL_X2 FILLER_5_74 ();
 FILLCELL_X1 FILLER_5_76 ();
 FILLCELL_X4 FILLER_5_98 ();
 FILLCELL_X2 FILLER_5_102 ();
 FILLCELL_X1 FILLER_5_104 ();
 FILLCELL_X8 FILLER_5_108 ();
 FILLCELL_X1 FILLER_5_116 ();
 FILLCELL_X16 FILLER_5_137 ();
 FILLCELL_X8 FILLER_5_153 ();
 FILLCELL_X4 FILLER_5_161 ();
 FILLCELL_X1 FILLER_5_165 ();
 FILLCELL_X32 FILLER_5_172 ();
 FILLCELL_X8 FILLER_5_209 ();
 FILLCELL_X1 FILLER_5_217 ();
 FILLCELL_X2 FILLER_5_223 ();
 FILLCELL_X16 FILLER_5_250 ();
 FILLCELL_X8 FILLER_5_266 ();
 FILLCELL_X1 FILLER_5_274 ();
 FILLCELL_X1 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_7 ();
 FILLCELL_X4 FILLER_6_23 ();
 FILLCELL_X1 FILLER_6_27 ();
 FILLCELL_X32 FILLER_6_34 ();
 FILLCELL_X16 FILLER_6_66 ();
 FILLCELL_X4 FILLER_6_82 ();
 FILLCELL_X2 FILLER_6_86 ();
 FILLCELL_X1 FILLER_6_88 ();
 FILLCELL_X2 FILLER_6_93 ();
 FILLCELL_X2 FILLER_6_98 ();
 FILLCELL_X1 FILLER_6_100 ();
 FILLCELL_X16 FILLER_6_105 ();
 FILLCELL_X2 FILLER_6_121 ();
 FILLCELL_X1 FILLER_6_123 ();
 FILLCELL_X8 FILLER_6_146 ();
 FILLCELL_X4 FILLER_6_154 ();
 FILLCELL_X2 FILLER_6_158 ();
 FILLCELL_X1 FILLER_6_160 ();
 FILLCELL_X16 FILLER_6_163 ();
 FILLCELL_X8 FILLER_6_179 ();
 FILLCELL_X2 FILLER_6_187 ();
 FILLCELL_X1 FILLER_6_189 ();
 FILLCELL_X32 FILLER_6_210 ();
 FILLCELL_X8 FILLER_6_242 ();
 FILLCELL_X4 FILLER_6_250 ();
 FILLCELL_X8 FILLER_6_265 ();
 FILLCELL_X2 FILLER_6_273 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_33 ();
 FILLCELL_X4 FILLER_7_41 ();
 FILLCELL_X1 FILLER_7_45 ();
 FILLCELL_X16 FILLER_7_49 ();
 FILLCELL_X1 FILLER_7_65 ();
 FILLCELL_X2 FILLER_7_85 ();
 FILLCELL_X1 FILLER_7_89 ();
 FILLCELL_X32 FILLER_7_114 ();
 FILLCELL_X16 FILLER_7_146 ();
 FILLCELL_X2 FILLER_7_166 ();
 FILLCELL_X16 FILLER_7_178 ();
 FILLCELL_X2 FILLER_7_194 ();
 FILLCELL_X1 FILLER_7_196 ();
 FILLCELL_X32 FILLER_7_206 ();
 FILLCELL_X16 FILLER_7_238 ();
 FILLCELL_X1 FILLER_7_254 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_56 ();
 FILLCELL_X4 FILLER_8_72 ();
 FILLCELL_X2 FILLER_8_76 ();
 FILLCELL_X4 FILLER_8_96 ();
 FILLCELL_X16 FILLER_8_117 ();
 FILLCELL_X8 FILLER_8_138 ();
 FILLCELL_X4 FILLER_8_146 ();
 FILLCELL_X2 FILLER_8_150 ();
 FILLCELL_X1 FILLER_8_152 ();
 FILLCELL_X1 FILLER_8_166 ();
 FILLCELL_X8 FILLER_8_175 ();
 FILLCELL_X2 FILLER_8_183 ();
 FILLCELL_X1 FILLER_8_196 ();
 FILLCELL_X8 FILLER_8_207 ();
 FILLCELL_X32 FILLER_8_221 ();
 FILLCELL_X16 FILLER_8_253 ();
 FILLCELL_X4 FILLER_8_269 ();
 FILLCELL_X2 FILLER_8_273 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_9 ();
 FILLCELL_X1 FILLER_9_13 ();
 FILLCELL_X8 FILLER_9_34 ();
 FILLCELL_X4 FILLER_9_42 ();
 FILLCELL_X1 FILLER_9_46 ();
 FILLCELL_X32 FILLER_9_53 ();
 FILLCELL_X4 FILLER_9_85 ();
 FILLCELL_X2 FILLER_9_89 ();
 FILLCELL_X32 FILLER_9_98 ();
 FILLCELL_X16 FILLER_9_130 ();
 FILLCELL_X2 FILLER_9_146 ();
 FILLCELL_X1 FILLER_9_148 ();
 FILLCELL_X16 FILLER_9_170 ();
 FILLCELL_X2 FILLER_9_186 ();
 FILLCELL_X1 FILLER_9_188 ();
 FILLCELL_X4 FILLER_9_199 ();
 FILLCELL_X2 FILLER_9_203 ();
 FILLCELL_X1 FILLER_9_220 ();
 FILLCELL_X1 FILLER_9_225 ();
 FILLCELL_X1 FILLER_9_230 ();
 FILLCELL_X2 FILLER_9_248 ();
 FILLCELL_X8 FILLER_9_261 ();
 FILLCELL_X4 FILLER_9_269 ();
 FILLCELL_X2 FILLER_9_273 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_17 ();
 FILLCELL_X4 FILLER_10_25 ();
 FILLCELL_X8 FILLER_10_39 ();
 FILLCELL_X4 FILLER_10_47 ();
 FILLCELL_X1 FILLER_10_51 ();
 FILLCELL_X32 FILLER_10_69 ();
 FILLCELL_X2 FILLER_10_101 ();
 FILLCELL_X1 FILLER_10_103 ();
 FILLCELL_X32 FILLER_10_112 ();
 FILLCELL_X32 FILLER_10_144 ();
 FILLCELL_X8 FILLER_10_176 ();
 FILLCELL_X2 FILLER_10_184 ();
 FILLCELL_X32 FILLER_10_188 ();
 FILLCELL_X32 FILLER_10_220 ();
 FILLCELL_X2 FILLER_10_252 ();
 FILLCELL_X1 FILLER_10_254 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_33 ();
 FILLCELL_X1 FILLER_11_38 ();
 FILLCELL_X2 FILLER_11_48 ();
 FILLCELL_X8 FILLER_11_53 ();
 FILLCELL_X1 FILLER_11_61 ();
 FILLCELL_X4 FILLER_11_78 ();
 FILLCELL_X2 FILLER_11_82 ();
 FILLCELL_X1 FILLER_11_84 ();
 FILLCELL_X16 FILLER_11_90 ();
 FILLCELL_X1 FILLER_11_106 ();
 FILLCELL_X2 FILLER_11_121 ();
 FILLCELL_X16 FILLER_11_142 ();
 FILLCELL_X4 FILLER_11_158 ();
 FILLCELL_X1 FILLER_11_162 ();
 FILLCELL_X4 FILLER_11_166 ();
 FILLCELL_X16 FILLER_11_174 ();
 FILLCELL_X2 FILLER_11_190 ();
 FILLCELL_X1 FILLER_11_192 ();
 FILLCELL_X2 FILLER_11_205 ();
 FILLCELL_X8 FILLER_11_211 ();
 FILLCELL_X2 FILLER_11_219 ();
 FILLCELL_X1 FILLER_11_221 ();
 FILLCELL_X1 FILLER_11_226 ();
 FILLCELL_X32 FILLER_11_231 ();
 FILLCELL_X8 FILLER_11_263 ();
 FILLCELL_X4 FILLER_11_271 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_5 ();
 FILLCELL_X2 FILLER_12_23 ();
 FILLCELL_X1 FILLER_12_25 ();
 FILLCELL_X8 FILLER_12_29 ();
 FILLCELL_X4 FILLER_12_37 ();
 FILLCELL_X2 FILLER_12_41 ();
 FILLCELL_X1 FILLER_12_43 ();
 FILLCELL_X4 FILLER_12_59 ();
 FILLCELL_X2 FILLER_12_63 ();
 FILLCELL_X2 FILLER_12_72 ();
 FILLCELL_X1 FILLER_12_86 ();
 FILLCELL_X32 FILLER_12_114 ();
 FILLCELL_X16 FILLER_12_146 ();
 FILLCELL_X1 FILLER_12_162 ();
 FILLCELL_X32 FILLER_12_167 ();
 FILLCELL_X4 FILLER_12_199 ();
 FILLCELL_X2 FILLER_12_203 ();
 FILLCELL_X8 FILLER_12_209 ();
 FILLCELL_X4 FILLER_12_217 ();
 FILLCELL_X2 FILLER_12_221 ();
 FILLCELL_X32 FILLER_12_240 ();
 FILLCELL_X2 FILLER_12_272 ();
 FILLCELL_X1 FILLER_12_274 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_17 ();
 FILLCELL_X16 FILLER_13_26 ();
 FILLCELL_X1 FILLER_13_42 ();
 FILLCELL_X16 FILLER_13_61 ();
 FILLCELL_X4 FILLER_13_77 ();
 FILLCELL_X2 FILLER_13_81 ();
 FILLCELL_X1 FILLER_13_83 ();
 FILLCELL_X2 FILLER_13_91 ();
 FILLCELL_X1 FILLER_13_98 ();
 FILLCELL_X1 FILLER_13_108 ();
 FILLCELL_X2 FILLER_13_117 ();
 FILLCELL_X16 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_145 ();
 FILLCELL_X4 FILLER_13_153 ();
 FILLCELL_X1 FILLER_13_157 ();
 FILLCELL_X16 FILLER_13_184 ();
 FILLCELL_X4 FILLER_13_200 ();
 FILLCELL_X1 FILLER_13_204 ();
 FILLCELL_X16 FILLER_13_222 ();
 FILLCELL_X8 FILLER_13_238 ();
 FILLCELL_X4 FILLER_13_246 ();
 FILLCELL_X8 FILLER_13_261 ();
 FILLCELL_X2 FILLER_13_272 ();
 FILLCELL_X1 FILLER_13_274 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X8 FILLER_14_17 ();
 FILLCELL_X2 FILLER_14_25 ();
 FILLCELL_X1 FILLER_14_27 ();
 FILLCELL_X16 FILLER_14_34 ();
 FILLCELL_X8 FILLER_14_50 ();
 FILLCELL_X2 FILLER_14_58 ();
 FILLCELL_X1 FILLER_14_60 ();
 FILLCELL_X8 FILLER_14_71 ();
 FILLCELL_X4 FILLER_14_79 ();
 FILLCELL_X8 FILLER_14_94 ();
 FILLCELL_X2 FILLER_14_102 ();
 FILLCELL_X1 FILLER_14_104 ();
 FILLCELL_X32 FILLER_14_144 ();
 FILLCELL_X4 FILLER_14_176 ();
 FILLCELL_X2 FILLER_14_180 ();
 FILLCELL_X16 FILLER_14_196 ();
 FILLCELL_X2 FILLER_14_212 ();
 FILLCELL_X1 FILLER_14_214 ();
 FILLCELL_X32 FILLER_14_220 ();
 FILLCELL_X4 FILLER_14_269 ();
 FILLCELL_X2 FILLER_14_273 ();
 FILLCELL_X2 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_24 ();
 FILLCELL_X1 FILLER_15_29 ();
 FILLCELL_X32 FILLER_15_37 ();
 FILLCELL_X16 FILLER_15_69 ();
 FILLCELL_X4 FILLER_15_85 ();
 FILLCELL_X2 FILLER_15_89 ();
 FILLCELL_X32 FILLER_15_98 ();
 FILLCELL_X8 FILLER_15_130 ();
 FILLCELL_X2 FILLER_15_138 ();
 FILLCELL_X1 FILLER_15_140 ();
 FILLCELL_X32 FILLER_15_145 ();
 FILLCELL_X4 FILLER_15_177 ();
 FILLCELL_X2 FILLER_15_181 ();
 FILLCELL_X16 FILLER_15_191 ();
 FILLCELL_X8 FILLER_15_207 ();
 FILLCELL_X1 FILLER_15_215 ();
 FILLCELL_X2 FILLER_15_240 ();
 FILLCELL_X1 FILLER_15_242 ();
 FILLCELL_X16 FILLER_15_246 ();
 FILLCELL_X8 FILLER_15_262 ();
 FILLCELL_X4 FILLER_15_270 ();
 FILLCELL_X1 FILLER_15_274 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X2 FILLER_16_27 ();
 FILLCELL_X2 FILLER_16_43 ();
 FILLCELL_X16 FILLER_16_50 ();
 FILLCELL_X8 FILLER_16_66 ();
 FILLCELL_X4 FILLER_16_74 ();
 FILLCELL_X2 FILLER_16_78 ();
 FILLCELL_X1 FILLER_16_80 ();
 FILLCELL_X32 FILLER_16_100 ();
 FILLCELL_X16 FILLER_16_132 ();
 FILLCELL_X4 FILLER_16_148 ();
 FILLCELL_X16 FILLER_16_165 ();
 FILLCELL_X4 FILLER_16_181 ();
 FILLCELL_X2 FILLER_16_185 ();
 FILLCELL_X16 FILLER_16_204 ();
 FILLCELL_X4 FILLER_16_220 ();
 FILLCELL_X16 FILLER_16_228 ();
 FILLCELL_X8 FILLER_16_244 ();
 FILLCELL_X4 FILLER_16_263 ();
 FILLCELL_X2 FILLER_16_267 ();
 FILLCELL_X2 FILLER_16_272 ();
 FILLCELL_X1 FILLER_16_274 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_41 ();
 FILLCELL_X1 FILLER_17_43 ();
 FILLCELL_X16 FILLER_17_51 ();
 FILLCELL_X8 FILLER_17_67 ();
 FILLCELL_X4 FILLER_17_75 ();
 FILLCELL_X1 FILLER_17_79 ();
 FILLCELL_X4 FILLER_17_87 ();
 FILLCELL_X2 FILLER_17_91 ();
 FILLCELL_X8 FILLER_17_130 ();
 FILLCELL_X2 FILLER_17_138 ();
 FILLCELL_X1 FILLER_17_140 ();
 FILLCELL_X32 FILLER_17_150 ();
 FILLCELL_X2 FILLER_17_182 ();
 FILLCELL_X1 FILLER_17_184 ();
 FILLCELL_X8 FILLER_17_202 ();
 FILLCELL_X4 FILLER_17_210 ();
 FILLCELL_X2 FILLER_17_214 ();
 FILLCELL_X16 FILLER_17_223 ();
 FILLCELL_X8 FILLER_17_239 ();
 FILLCELL_X4 FILLER_17_247 ();
 FILLCELL_X2 FILLER_17_251 ();
 FILLCELL_X1 FILLER_17_253 ();
 FILLCELL_X4 FILLER_17_271 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_33 ();
 FILLCELL_X4 FILLER_18_41 ();
 FILLCELL_X1 FILLER_18_45 ();
 FILLCELL_X8 FILLER_18_64 ();
 FILLCELL_X1 FILLER_18_72 ();
 FILLCELL_X2 FILLER_18_91 ();
 FILLCELL_X1 FILLER_18_93 ();
 FILLCELL_X4 FILLER_18_103 ();
 FILLCELL_X2 FILLER_18_107 ();
 FILLCELL_X1 FILLER_18_109 ();
 FILLCELL_X2 FILLER_18_136 ();
 FILLCELL_X32 FILLER_18_153 ();
 FILLCELL_X16 FILLER_18_185 ();
 FILLCELL_X4 FILLER_18_201 ();
 FILLCELL_X2 FILLER_18_205 ();
 FILLCELL_X8 FILLER_18_218 ();
 FILLCELL_X4 FILLER_18_226 ();
 FILLCELL_X1 FILLER_18_230 ();
 FILLCELL_X16 FILLER_18_235 ();
 FILLCELL_X2 FILLER_18_251 ();
 FILLCELL_X4 FILLER_18_260 ();
 FILLCELL_X2 FILLER_18_264 ();
 FILLCELL_X1 FILLER_18_266 ();
 FILLCELL_X2 FILLER_18_270 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_33 ();
 FILLCELL_X1 FILLER_19_48 ();
 FILLCELL_X32 FILLER_19_58 ();
 FILLCELL_X16 FILLER_19_90 ();
 FILLCELL_X8 FILLER_19_106 ();
 FILLCELL_X2 FILLER_19_114 ();
 FILLCELL_X1 FILLER_19_116 ();
 FILLCELL_X8 FILLER_19_120 ();
 FILLCELL_X4 FILLER_19_128 ();
 FILLCELL_X32 FILLER_19_150 ();
 FILLCELL_X32 FILLER_19_182 ();
 FILLCELL_X4 FILLER_19_214 ();
 FILLCELL_X4 FILLER_19_252 ();
 FILLCELL_X2 FILLER_19_256 ();
 FILLCELL_X8 FILLER_19_262 ();
 FILLCELL_X4 FILLER_19_270 ();
 FILLCELL_X1 FILLER_19_274 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_41 ();
 FILLCELL_X2 FILLER_20_45 ();
 FILLCELL_X1 FILLER_20_49 ();
 FILLCELL_X32 FILLER_20_60 ();
 FILLCELL_X16 FILLER_20_92 ();
 FILLCELL_X4 FILLER_20_108 ();
 FILLCELL_X2 FILLER_20_112 ();
 FILLCELL_X8 FILLER_20_124 ();
 FILLCELL_X1 FILLER_20_132 ();
 FILLCELL_X32 FILLER_20_157 ();
 FILLCELL_X32 FILLER_20_189 ();
 FILLCELL_X32 FILLER_20_221 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X2 FILLER_20_272 ();
 FILLCELL_X1 FILLER_20_274 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_25 ();
 FILLCELL_X1 FILLER_21_27 ();
 FILLCELL_X8 FILLER_21_31 ();
 FILLCELL_X16 FILLER_21_49 ();
 FILLCELL_X1 FILLER_21_65 ();
 FILLCELL_X1 FILLER_21_73 ();
 FILLCELL_X2 FILLER_21_92 ();
 FILLCELL_X4 FILLER_21_106 ();
 FILLCELL_X2 FILLER_21_110 ();
 FILLCELL_X8 FILLER_21_115 ();
 FILLCELL_X4 FILLER_21_132 ();
 FILLCELL_X32 FILLER_21_160 ();
 FILLCELL_X32 FILLER_21_192 ();
 FILLCELL_X32 FILLER_21_224 ();
 FILLCELL_X16 FILLER_21_256 ();
 FILLCELL_X2 FILLER_21_272 ();
 FILLCELL_X1 FILLER_21_274 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_17 ();
 FILLCELL_X4 FILLER_22_25 ();
 FILLCELL_X2 FILLER_22_35 ();
 FILLCELL_X2 FILLER_22_42 ();
 FILLCELL_X1 FILLER_22_44 ();
 FILLCELL_X8 FILLER_22_47 ();
 FILLCELL_X4 FILLER_22_55 ();
 FILLCELL_X2 FILLER_22_59 ();
 FILLCELL_X1 FILLER_22_83 ();
 FILLCELL_X16 FILLER_22_91 ();
 FILLCELL_X4 FILLER_22_107 ();
 FILLCELL_X2 FILLER_22_111 ();
 FILLCELL_X1 FILLER_22_113 ();
 FILLCELL_X32 FILLER_22_146 ();
 FILLCELL_X4 FILLER_22_178 ();
 FILLCELL_X8 FILLER_22_199 ();
 FILLCELL_X1 FILLER_22_207 ();
 FILLCELL_X32 FILLER_22_218 ();
 FILLCELL_X16 FILLER_22_250 ();
 FILLCELL_X8 FILLER_22_266 ();
 FILLCELL_X1 FILLER_22_274 ();
 FILLCELL_X8 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_9 ();
 FILLCELL_X2 FILLER_23_13 ();
 FILLCELL_X8 FILLER_23_37 ();
 FILLCELL_X2 FILLER_23_45 ();
 FILLCELL_X4 FILLER_23_65 ();
 FILLCELL_X8 FILLER_23_86 ();
 FILLCELL_X4 FILLER_23_94 ();
 FILLCELL_X2 FILLER_23_98 ();
 FILLCELL_X32 FILLER_23_105 ();
 FILLCELL_X16 FILLER_23_137 ();
 FILLCELL_X8 FILLER_23_153 ();
 FILLCELL_X1 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_184 ();
 FILLCELL_X1 FILLER_23_188 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X16 FILLER_23_257 ();
 FILLCELL_X2 FILLER_23_273 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X8 FILLER_24_17 ();
 FILLCELL_X4 FILLER_24_25 ();
 FILLCELL_X2 FILLER_24_29 ();
 FILLCELL_X32 FILLER_24_39 ();
 FILLCELL_X4 FILLER_24_71 ();
 FILLCELL_X2 FILLER_24_75 ();
 FILLCELL_X1 FILLER_24_77 ();
 FILLCELL_X1 FILLER_24_85 ();
 FILLCELL_X4 FILLER_24_95 ();
 FILLCELL_X2 FILLER_24_99 ();
 FILLCELL_X1 FILLER_24_101 ();
 FILLCELL_X16 FILLER_24_108 ();
 FILLCELL_X8 FILLER_24_124 ();
 FILLCELL_X2 FILLER_24_132 ();
 FILLCELL_X4 FILLER_24_136 ();
 FILLCELL_X2 FILLER_24_140 ();
 FILLCELL_X16 FILLER_24_147 ();
 FILLCELL_X8 FILLER_24_163 ();
 FILLCELL_X1 FILLER_24_171 ();
 FILLCELL_X32 FILLER_24_187 ();
 FILLCELL_X32 FILLER_24_219 ();
 FILLCELL_X16 FILLER_24_251 ();
 FILLCELL_X8 FILLER_24_267 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X16 FILLER_25_65 ();
 FILLCELL_X8 FILLER_25_91 ();
 FILLCELL_X2 FILLER_25_99 ();
 FILLCELL_X16 FILLER_25_118 ();
 FILLCELL_X8 FILLER_25_152 ();
 FILLCELL_X2 FILLER_25_160 ();
 FILLCELL_X32 FILLER_25_186 ();
 FILLCELL_X32 FILLER_25_218 ();
 FILLCELL_X16 FILLER_25_250 ();
 FILLCELL_X8 FILLER_25_266 ();
 FILLCELL_X1 FILLER_25_274 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_17 ();
 FILLCELL_X2 FILLER_26_21 ();
 FILLCELL_X1 FILLER_26_23 ();
 FILLCELL_X8 FILLER_26_42 ();
 FILLCELL_X16 FILLER_26_55 ();
 FILLCELL_X8 FILLER_26_71 ();
 FILLCELL_X4 FILLER_26_79 ();
 FILLCELL_X1 FILLER_26_83 ();
 FILLCELL_X8 FILLER_26_89 ();
 FILLCELL_X1 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_115 ();
 FILLCELL_X16 FILLER_26_147 ();
 FILLCELL_X2 FILLER_26_163 ();
 FILLCELL_X2 FILLER_26_174 ();
 FILLCELL_X1 FILLER_26_176 ();
 FILLCELL_X32 FILLER_26_190 ();
 FILLCELL_X32 FILLER_26_222 ();
 FILLCELL_X16 FILLER_26_254 ();
 FILLCELL_X4 FILLER_26_270 ();
 FILLCELL_X1 FILLER_26_274 ();
 FILLCELL_X8 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_9 ();
 FILLCELL_X2 FILLER_27_33 ();
 FILLCELL_X1 FILLER_27_35 ();
 FILLCELL_X16 FILLER_27_64 ();
 FILLCELL_X2 FILLER_27_80 ();
 FILLCELL_X1 FILLER_27_82 ();
 FILLCELL_X16 FILLER_27_89 ();
 FILLCELL_X2 FILLER_27_105 ();
 FILLCELL_X1 FILLER_27_107 ();
 FILLCELL_X32 FILLER_27_133 ();
 FILLCELL_X4 FILLER_27_165 ();
 FILLCELL_X2 FILLER_27_169 ();
 FILLCELL_X1 FILLER_27_171 ();
 FILLCELL_X32 FILLER_27_181 ();
 FILLCELL_X32 FILLER_27_213 ();
 FILLCELL_X16 FILLER_27_245 ();
 FILLCELL_X8 FILLER_27_261 ();
 FILLCELL_X4 FILLER_27_269 ();
 FILLCELL_X2 FILLER_27_273 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X8 FILLER_28_17 ();
 FILLCELL_X4 FILLER_28_25 ();
 FILLCELL_X2 FILLER_28_29 ();
 FILLCELL_X8 FILLER_28_37 ();
 FILLCELL_X1 FILLER_28_45 ();
 FILLCELL_X16 FILLER_28_55 ();
 FILLCELL_X8 FILLER_28_71 ();
 FILLCELL_X1 FILLER_28_79 ();
 FILLCELL_X32 FILLER_28_83 ();
 FILLCELL_X8 FILLER_28_115 ();
 FILLCELL_X2 FILLER_28_123 ();
 FILLCELL_X1 FILLER_28_125 ();
 FILLCELL_X16 FILLER_28_132 ();
 FILLCELL_X8 FILLER_28_148 ();
 FILLCELL_X2 FILLER_28_156 ();
 FILLCELL_X1 FILLER_28_158 ();
 FILLCELL_X2 FILLER_28_178 ();
 FILLCELL_X1 FILLER_28_180 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X16 FILLER_28_257 ();
 FILLCELL_X2 FILLER_28_273 ();
 FILLCELL_X16 FILLER_29_1 ();
 FILLCELL_X8 FILLER_29_17 ();
 FILLCELL_X4 FILLER_29_25 ();
 FILLCELL_X2 FILLER_29_29 ();
 FILLCELL_X4 FILLER_29_34 ();
 FILLCELL_X2 FILLER_29_38 ();
 FILLCELL_X1 FILLER_29_40 ();
 FILLCELL_X4 FILLER_29_46 ();
 FILLCELL_X2 FILLER_29_50 ();
 FILLCELL_X8 FILLER_29_70 ();
 FILLCELL_X32 FILLER_29_99 ();
 FILLCELL_X16 FILLER_29_131 ();
 FILLCELL_X2 FILLER_29_147 ();
 FILLCELL_X1 FILLER_29_149 ();
 FILLCELL_X4 FILLER_29_153 ();
 FILLCELL_X2 FILLER_29_157 ();
 FILLCELL_X8 FILLER_29_165 ();
 FILLCELL_X4 FILLER_29_173 ();
 FILLCELL_X1 FILLER_29_179 ();
 FILLCELL_X32 FILLER_29_199 ();
 FILLCELL_X32 FILLER_29_231 ();
 FILLCELL_X8 FILLER_29_263 ();
 FILLCELL_X4 FILLER_29_271 ();
 FILLCELL_X16 FILLER_30_1 ();
 FILLCELL_X8 FILLER_30_17 ();
 FILLCELL_X2 FILLER_30_25 ();
 FILLCELL_X32 FILLER_30_44 ();
 FILLCELL_X1 FILLER_30_76 ();
 FILLCELL_X16 FILLER_30_83 ();
 FILLCELL_X8 FILLER_30_99 ();
 FILLCELL_X2 FILLER_30_107 ();
 FILLCELL_X8 FILLER_30_132 ();
 FILLCELL_X2 FILLER_30_140 ();
 FILLCELL_X8 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_169 ();
 FILLCELL_X2 FILLER_30_173 ();
 FILLCELL_X32 FILLER_30_191 ();
 FILLCELL_X32 FILLER_30_223 ();
 FILLCELL_X16 FILLER_30_255 ();
 FILLCELL_X4 FILLER_30_271 ();
 FILLCELL_X16 FILLER_31_1 ();
 FILLCELL_X8 FILLER_31_17 ();
 FILLCELL_X4 FILLER_31_25 ();
 FILLCELL_X1 FILLER_31_42 ();
 FILLCELL_X1 FILLER_31_48 ();
 FILLCELL_X16 FILLER_31_55 ();
 FILLCELL_X8 FILLER_31_71 ();
 FILLCELL_X8 FILLER_31_82 ();
 FILLCELL_X2 FILLER_31_90 ();
 FILLCELL_X16 FILLER_31_96 ();
 FILLCELL_X4 FILLER_31_112 ();
 FILLCELL_X2 FILLER_31_116 ();
 FILLCELL_X1 FILLER_31_130 ();
 FILLCELL_X16 FILLER_31_136 ();
 FILLCELL_X8 FILLER_31_152 ();
 FILLCELL_X2 FILLER_31_160 ();
 FILLCELL_X1 FILLER_31_166 ();
 FILLCELL_X1 FILLER_31_185 ();
 FILLCELL_X1 FILLER_31_188 ();
 FILLCELL_X32 FILLER_31_192 ();
 FILLCELL_X32 FILLER_31_224 ();
 FILLCELL_X16 FILLER_31_256 ();
 FILLCELL_X2 FILLER_31_272 ();
 FILLCELL_X1 FILLER_31_274 ();
 FILLCELL_X16 FILLER_32_1 ();
 FILLCELL_X8 FILLER_32_17 ();
 FILLCELL_X4 FILLER_32_25 ();
 FILLCELL_X2 FILLER_32_29 ();
 FILLCELL_X8 FILLER_32_34 ();
 FILLCELL_X2 FILLER_32_42 ();
 FILLCELL_X8 FILLER_32_63 ();
 FILLCELL_X4 FILLER_32_71 ();
 FILLCELL_X2 FILLER_32_75 ();
 FILLCELL_X16 FILLER_32_94 ();
 FILLCELL_X4 FILLER_32_110 ();
 FILLCELL_X2 FILLER_32_114 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X2 FILLER_32_161 ();
 FILLCELL_X8 FILLER_32_167 ();
 FILLCELL_X2 FILLER_32_175 ();
 FILLCELL_X8 FILLER_32_180 ();
 FILLCELL_X4 FILLER_32_188 ();
 FILLCELL_X32 FILLER_32_211 ();
 FILLCELL_X32 FILLER_32_243 ();
 FILLCELL_X16 FILLER_33_1 ();
 FILLCELL_X8 FILLER_33_17 ();
 FILLCELL_X2 FILLER_33_25 ();
 FILLCELL_X1 FILLER_33_27 ();
 FILLCELL_X4 FILLER_33_45 ();
 FILLCELL_X32 FILLER_33_52 ();
 FILLCELL_X16 FILLER_33_84 ();
 FILLCELL_X8 FILLER_33_100 ();
 FILLCELL_X2 FILLER_33_108 ();
 FILLCELL_X32 FILLER_33_127 ();
 FILLCELL_X1 FILLER_33_159 ();
 FILLCELL_X1 FILLER_33_169 ();
 FILLCELL_X32 FILLER_33_179 ();
 FILLCELL_X32 FILLER_33_211 ();
 FILLCELL_X32 FILLER_33_243 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X16 FILLER_34_129 ();
 FILLCELL_X4 FILLER_34_168 ();
 FILLCELL_X2 FILLER_34_172 ();
 FILLCELL_X1 FILLER_34_174 ();
 FILLCELL_X4 FILLER_34_179 ();
 FILLCELL_X1 FILLER_34_183 ();
 FILLCELL_X32 FILLER_34_188 ();
 FILLCELL_X32 FILLER_34_220 ();
 FILLCELL_X16 FILLER_34_252 ();
 FILLCELL_X4 FILLER_34_268 ();
 FILLCELL_X2 FILLER_34_272 ();
 FILLCELL_X1 FILLER_34_274 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X8 FILLER_35_161 ();
 FILLCELL_X4 FILLER_35_169 ();
 FILLCELL_X1 FILLER_35_173 ();
 FILLCELL_X32 FILLER_35_191 ();
 FILLCELL_X32 FILLER_35_223 ();
 FILLCELL_X16 FILLER_35_255 ();
 FILLCELL_X4 FILLER_35_271 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X16 FILLER_36_257 ();
 FILLCELL_X2 FILLER_36_273 ();
endmodule
