module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire net1;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire \ctrl$a_reg_en ;
 wire \ctrl$b_reg_en ;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire \dpath.a_mux$out[0] ;
 wire \dpath.a_mux$out[10] ;
 wire \dpath.a_mux$out[11] ;
 wire \dpath.a_mux$out[12] ;
 wire \dpath.a_mux$out[13] ;
 wire \dpath.a_mux$out[14] ;
 wire \dpath.a_mux$out[15] ;
 wire \dpath.a_mux$out[1] ;
 wire \dpath.a_mux$out[2] ;
 wire \dpath.a_mux$out[3] ;
 wire \dpath.a_mux$out[4] ;
 wire \dpath.a_mux$out[5] ;
 wire \dpath.a_mux$out[6] ;
 wire \dpath.a_mux$out[7] ;
 wire \dpath.a_mux$out[8] ;
 wire \dpath.a_mux$out[9] ;
 wire \dpath.b_mux$out[0] ;
 wire \dpath.b_mux$out[10] ;
 wire \dpath.b_mux$out[11] ;
 wire \dpath.b_mux$out[12] ;
 wire \dpath.b_mux$out[13] ;
 wire \dpath.b_mux$out[14] ;
 wire \dpath.b_mux$out[15] ;
 wire \dpath.b_mux$out[1] ;
 wire \dpath.b_mux$out[2] ;
 wire \dpath.b_mux$out[3] ;
 wire \dpath.b_mux$out[4] ;
 wire \dpath.b_mux$out[5] ;
 wire \dpath.b_mux$out[6] ;
 wire \dpath.b_mux$out[7] ;
 wire \dpath.b_mux$out[8] ;
 wire \dpath.b_mux$out[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net86;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net119;
 wire net74;
 wire net75;
 wire net80;
 wire net81;
 wire net82;
 wire net134;
 wire net84;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net227;
 wire net110;
 wire net111;
 wire net112;
 wire net217;
 wire net216;
 wire net215;
 wire net116;
 wire net117;
 wire net118;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net85;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net135;
 wire net136;
 wire net137;

 sky130_fd_sc_hd__and2b_2 _243_ (.A_N(\dpath.a_lt_b$in0[0] ),
    .B(\dpath.a_lt_b$in1[0] ),
    .X(_003_));
 sky130_fd_sc_hd__or2b_1 _244_ (.A(net75),
    .B_N(net60),
    .X(_004_));
 sky130_fd_sc_hd__nand2b_1 _245_ (.A_N(_003_),
    .B(_004_),
    .Y(net38));
 sky130_fd_sc_hd__buf_4 _246_ (.A(net37),
    .X(_005_));
 sky130_fd_sc_hd__clkbuf_4 _247_ (.A(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nor4_1 _248_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(net89),
    .C(\dpath.a_lt_b$in1[4] ),
    .D(net309),
    .Y(_007_));
 sky130_fd_sc_hd__buf_4 _249_ (.A(\dpath.a_lt_b$in1[12] ),
    .X(_008_));
 sky130_fd_sc_hd__buf_2 _250_ (.A(\dpath.a_lt_b$in1[11] ),
    .X(_009_));
 sky130_fd_sc_hd__nor4_4 _251_ (.A(_008_),
    .B(_009_),
    .C(net116),
    .D(net125),
    .Y(_010_));
 sky130_fd_sc_hd__buf_6 _252_ (.A(\dpath.a_lt_b$in1[5] ),
    .X(_011_));
 sky130_fd_sc_hd__clkbuf_2 _253_ (.A(\dpath.a_lt_b$in1[3] ),
    .X(_012_));
 sky130_fd_sc_hd__nor2_2 _254_ (.A(_012_),
    .B(net135),
    .Y(_013_));
 sky130_fd_sc_hd__clkbuf_2 _255_ (.A(\dpath.a_lt_b$in1[1] ),
    .X(_014_));
 sky130_fd_sc_hd__nor2_1 _256_ (.A(_014_),
    .B(net77),
    .Y(_015_));
 sky130_fd_sc_hd__buf_6 _257_ (.A(\dpath.a_lt_b$in1[13] ),
    .X(_016_));
 sky130_fd_sc_hd__nor4_1 _258_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(net123),
    .C(net96),
    .D(net311),
    .Y(_017_));
 sky130_fd_sc_hd__and3_1 _259_ (.A(net215),
    .B(_015_),
    .C(_017_),
    .X(_018_));
 sky130_fd_sc_hd__nand3_2 _260_ (.A(_007_),
    .B(_018_),
    .C(_010_),
    .Y(_019_));
 sky130_fd_sc_hd__a22oi_1 _261_ (.A1(_006_),
    .A2(net34),
    .B1(\ctrl.state.out[2] ),
    .B2(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__nor2_1 _262_ (.A(net35),
    .B(_020_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_1 _263_ (.A(\ctrl.state.out[1] ),
    .Y(_021_));
 sky130_fd_sc_hd__or2_4 _264_ (.A(net37),
    .B(\ctrl.state.out[2] ),
    .X(\ctrl$a_reg_en ));
 sky130_fd_sc_hd__nor2_1 _265_ (.A(_021_),
    .B(\ctrl$a_reg_en ),
    .Y(net54));
 sky130_fd_sc_hd__inv_1 _266_ (.A(net34),
    .Y(_022_));
 sky130_fd_sc_hd__a221o_1 _267_ (.A1(_006_),
    .A2(_022_),
    .B1(net36),
    .B2(net54),
    .C1(net35),
    .X(_000_));
 sky130_fd_sc_hd__inv_1 _268_ (.A(net36),
    .Y(_023_));
 sky130_fd_sc_hd__o21ai_0 _269_ (.A1(_006_),
    .A2(_023_),
    .B1(\ctrl.state.out[1] ),
    .Y(_024_));
 sky130_fd_sc_hd__a21bo_1 _270_ (.A1(_021_),
    .A2(_019_),
    .B1_N(\ctrl.state.out[2] ),
    .X(_025_));
 sky130_fd_sc_hd__a21oi_1 _271_ (.A1(_024_),
    .A2(_025_),
    .B1(net35),
    .Y(_001_));
 sky130_fd_sc_hd__a21o_4 clone1 (.A1(_106_),
    .A2(\ctrl.state.out[2] ),
    .B1(_107_),
    .X(net1));
 sky130_fd_sc_hd__xnor2_4 _273_ (.A(_008_),
    .B(\dpath.a_lt_b$in0[12] ),
    .Y(_027_));
 sky130_fd_sc_hd__nand2b_2 _274_ (.A_N(\dpath.a_lt_b$in0[14] ),
    .B(\dpath.a_lt_b$in1[14] ),
    .Y(_028_));
 sky130_fd_sc_hd__nand2b_2 _275_ (.A_N(\dpath.a_lt_b$in1[14] ),
    .B(\dpath.a_lt_b$in0[14] ),
    .Y(_029_));
 sky130_fd_sc_hd__nand2b_1 _276_ (.A_N(_016_),
    .B(\dpath.a_lt_b$in0[13] ),
    .Y(_030_));
 sky130_fd_sc_hd__nand2b_4 _277_ (.A_N(\dpath.a_lt_b$in0[13] ),
    .B(_016_),
    .Y(_031_));
 sky130_fd_sc_hd__and2_4 _278_ (.A(_031_),
    .B(_030_),
    .X(_032_));
 sky130_fd_sc_hd__nand4_4 _279_ (.A(_027_),
    .B(_028_),
    .C(_029_),
    .D(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__buf_2 _280_ (.A(\dpath.a_lt_b$in0[11] ),
    .X(_034_));
 sky130_fd_sc_hd__xor2_2 _281_ (.A(_034_),
    .B(_009_),
    .X(_035_));
 sky130_fd_sc_hd__nor2_4 _282_ (.A(_035_),
    .B(_033_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2b_4 _283_ (.A(\dpath.a_lt_b$in0[8] ),
    .B_N(net312),
    .Y(_037_));
 sky130_fd_sc_hd__nor2b_1 _284_ (.A(\dpath.a_lt_b$in1[8] ),
    .B_N(\dpath.a_lt_b$in0[8] ),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_2 _285_ (.A(_038_),
    .B(_037_),
    .Y(_039_));
 sky130_fd_sc_hd__nor2b_4 _286_ (.A(\dpath.a_lt_b$in1[10] ),
    .B_N(\dpath.a_lt_b$in0[10] ),
    .Y(_040_));
 sky130_fd_sc_hd__nor2b_4 _287_ (.A(net112),
    .B_N(\dpath.a_lt_b$in1[10] ),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_2 _288_ (.A(_041_),
    .B(_040_),
    .Y(_042_));
 sky130_fd_sc_hd__inv_1 _289_ (.A(\dpath.a_lt_b$in1[9] ),
    .Y(_043_));
 sky130_fd_sc_hd__nor2_1 _290_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _291_ (.A(\dpath.a_lt_b$in0[9] ),
    .Y(_045_));
 sky130_fd_sc_hd__nor2_1 _292_ (.A(_045_),
    .B(net99),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_2 _293_ (.A(_046_),
    .B(_044_),
    .Y(_047_));
 sky130_fd_sc_hd__and3_4 _294_ (.A(_039_),
    .B(_042_),
    .C(_047_),
    .X(_048_));
 sky130_fd_sc_hd__xnor2_2 _295_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(\dpath.a_lt_b$in1[15] ),
    .Y(_049_));
 sky130_fd_sc_hd__nand3_4 _296_ (.A(net119),
    .B(_048_),
    .C(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__buf_6 _297_ (.A(\dpath.a_lt_b$in0[7] ),
    .X(_051_));
 sky130_fd_sc_hd__xor2_4 _298_ (.A(_051_),
    .B(net110),
    .X(_052_));
 sky130_fd_sc_hd__nor2b_2 _299_ (.A(net63),
    .B_N(net87),
    .Y(_053_));
 sky130_fd_sc_hd__nor2b_2 _300_ (.A(net87),
    .B_N(\dpath.a_lt_b$in0[6] ),
    .Y(_054_));
 sky130_fd_sc_hd__xor2_2 _301_ (.A(\dpath.a_lt_b$in0[5] ),
    .B(_011_),
    .X(_055_));
 sky130_fd_sc_hd__nor4_4 _302_ (.A(_055_),
    .B(_052_),
    .C(_054_),
    .D(_053_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2b_1 _303_ (.A(\dpath.a_lt_b$in0[4] ),
    .B_N(\dpath.a_lt_b$in1[4] ),
    .Y(_057_));
 sky130_fd_sc_hd__nor2b_1 _304_ (.A(\dpath.a_lt_b$in1[4] ),
    .B_N(\dpath.a_lt_b$in0[4] ),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _305_ (.A(_057_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__xnor2_1 _306_ (.A(\dpath.a_lt_b$in0[3] ),
    .B(_012_),
    .Y(_060_));
 sky130_fd_sc_hd__nand2b_1 _307_ (.A_N(\dpath.a_lt_b$in0[2] ),
    .B(net308),
    .Y(_061_));
 sky130_fd_sc_hd__nand2b_1 _308_ (.A_N(\dpath.a_lt_b$in1[2] ),
    .B(\dpath.a_lt_b$in0[2] ),
    .Y(_062_));
 sky130_fd_sc_hd__and2_0 _309_ (.A(_061_),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__nand4_1 _310_ (.A(_056_),
    .B(_059_),
    .C(_060_),
    .D(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__xnor2_1 _311_ (.A(\dpath.a_lt_b$in0[1] ),
    .B(_014_),
    .Y(_065_));
 sky130_fd_sc_hd__or4b_4 _312_ (.A(net38),
    .B(_050_),
    .C(_064_),
    .D_N(_065_),
    .X(_066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__inv_1 _314_ (.A(\dpath.a_lt_b$in0[3] ),
    .Y(_068_));
 sky130_fd_sc_hd__nor2b_2 _315_ (.A(\dpath.a_lt_b$in0[2] ),
    .B_N(net308),
    .Y(_069_));
 sky130_fd_sc_hd__maj3_2 _316_ (.A(_068_),
    .B(_012_),
    .C(_069_),
    .X(_070_));
 sky130_fd_sc_hd__inv_1 _317_ (.A(\dpath.a_lt_b$in0[5] ),
    .Y(_071_));
 sky130_fd_sc_hd__o21ai_1 _318_ (.A1(\dpath.a_lt_b$in0[3] ),
    .A2(_061_),
    .B1(_013_),
    .Y(_072_));
 sky130_fd_sc_hd__a21oi_2 _319_ (.A1(_072_),
    .A2(_071_),
    .B1(\dpath.a_lt_b$in1[4] ),
    .Y(_073_));
 sky130_fd_sc_hd__nand2b_1 _320_ (.A_N(_070_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__o31a_1 _321_ (.A1(\dpath.a_lt_b$in1[4] ),
    .A2(_068_),
    .A3(_069_),
    .B1(_071_),
    .X(_075_));
 sky130_fd_sc_hd__nand2_1 _322_ (.A(\dpath.a_lt_b$in0[5] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .Y(_076_));
 sky130_fd_sc_hd__nor3_1 _323_ (.A(_052_),
    .B(_053_),
    .C(_054_),
    .Y(_077_));
 sky130_fd_sc_hd__o221a_1 _324_ (.A1(net135),
    .A2(_075_),
    .B1(_076_),
    .B2(_070_),
    .C1(_077_),
    .X(_078_));
 sky130_fd_sc_hd__a21oi_2 _325_ (.A1(_070_),
    .A2(\dpath.a_lt_b$in1[4] ),
    .B1(net135),
    .Y(_079_));
 sky130_fd_sc_hd__o21ai_2 _326_ (.A1(_073_),
    .A2(_079_),
    .B1(\dpath.a_lt_b$in0[4] ),
    .Y(_080_));
 sky130_fd_sc_hd__a21oi_1 _327_ (.A1(net60),
    .A2(_015_),
    .B1(\dpath.a_lt_b$in0[1] ),
    .Y(_081_));
 sky130_fd_sc_hd__a21oi_1 _328_ (.A1(_014_),
    .A2(_004_),
    .B1(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__inv_1 _329_ (.A(\dpath.a_lt_b$in1[7] ),
    .Y(_083_));
 sky130_fd_sc_hd__nand2b_4 _330_ (.A_N(\dpath.a_lt_b$in0[6] ),
    .B(\dpath.a_lt_b$in1[6] ),
    .Y(_084_));
 sky130_fd_sc_hd__maj3_2 _331_ (.A(_084_),
    .B(_051_),
    .C(_083_),
    .X(_085_));
 sky130_fd_sc_hd__o21ai_2 _332_ (.A1(_082_),
    .A2(net104),
    .B1(net68),
    .Y(_086_));
 sky130_fd_sc_hd__a31oi_4 _333_ (.A1(_074_),
    .A2(_078_),
    .A3(_080_),
    .B1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__inv_1 _334_ (.A(\dpath.a_lt_b$in0[15] ),
    .Y(_088_));
 sky130_fd_sc_hd__inv_1 _335_ (.A(_008_),
    .Y(_089_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(_089_),
    .B(net105),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_1 _337_ (.A(net122),
    .B(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__inv_1 _338_ (.A(\dpath.a_lt_b$in0[13] ),
    .Y(_092_));
 sky130_fd_sc_hd__o21ai_0 _339_ (.A1(net122),
    .A2(_090_),
    .B1(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__nand3_1 _340_ (.A(_028_),
    .B(_091_),
    .C(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_1 _341_ (.A(_009_),
    .Y(_095_));
 sky130_fd_sc_hd__inv_1 _342_ (.A(_041_),
    .Y(_096_));
 sky130_fd_sc_hd__nand2_1 _343_ (.A(net102),
    .B(_037_),
    .Y(_097_));
 sky130_fd_sc_hd__o21ai_0 _344_ (.A1(net100),
    .A2(_037_),
    .B1(net128),
    .Y(_098_));
 sky130_fd_sc_hd__o2111a_1 _345_ (.A1(_034_),
    .A2(_095_),
    .B1(_096_),
    .C1(_097_),
    .D1(_098_),
    .X(_099_));
 sky130_fd_sc_hd__maj3_1 _346_ (.A(_034_),
    .B(_095_),
    .C(_040_),
    .X(_100_));
 sky130_fd_sc_hd__nor3_1 _347_ (.A(_033_),
    .B(_099_),
    .C(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__a221oi_2 _348_ (.A1(_088_),
    .A2(\dpath.a_lt_b$in1[15] ),
    .B1(_029_),
    .B2(_094_),
    .C1(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__nor2_1 _349_ (.A(_088_),
    .B(\dpath.a_lt_b$in1[15] ),
    .Y(_103_));
 sky130_fd_sc_hd__o22ai_4 _350_ (.A1(_050_),
    .A2(_087_),
    .B1(_102_),
    .B2(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__and2_4 _351_ (.A(_104_),
    .B(_066_),
    .X(_105_));
 sky130_fd_sc_hd__buf_12 _352_ (.A(_105_),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_4 _353_ (.A(_005_),
    .X(_107_));
 sky130_fd_sc_hd__a21o_4 _354_ (.A1(\ctrl.state.out[2] ),
    .A2(_106_),
    .B1(_107_),
    .X(\ctrl$b_reg_en ));
 sky130_fd_sc_hd__nand2b_2 _355_ (.A_N(_005_),
    .B(\ctrl.state.out[2] ),
    .Y(_108_));
 sky130_fd_sc_hd__clkbuf_4 _356_ (.A(_108_),
    .X(_109_));
 sky130_fd_sc_hd__a21boi_2 _357_ (.A1(_104_),
    .A2(net93),
    .B1_N(net61),
    .Y(_110_));
 sky130_fd_sc_hd__xnor2_1 _358_ (.A(_110_),
    .B(net59),
    .Y(_111_));
 sky130_fd_sc_hd__nand2_1 _359_ (.A(net9),
    .B(_109_),
    .Y(_112_));
 sky130_fd_sc_hd__o21ai_1 _360_ (.A1(_111_),
    .A2(_109_),
    .B1(_112_),
    .Y(\dpath.a_mux$out[0] ));
 sky130_fd_sc_hd__maj3_1 _361_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(_043_),
    .C(_038_),
    .X(_113_));
 sky130_fd_sc_hd__a211oi_2 _362_ (.A1(net107),
    .A2(_083_),
    .B1(_054_),
    .C1(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__inv_1 _363_ (.A(\dpath.a_lt_b$in0[1] ),
    .Y(_115_));
 sky130_fd_sc_hd__maj3_2 _364_ (.A(_115_),
    .B(_014_),
    .C(_003_),
    .X(_116_));
 sky130_fd_sc_hd__a211oi_4 _365_ (.A1(_062_),
    .A2(_116_),
    .B1(_012_),
    .C1(_069_),
    .Y(_117_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_014_),
    .B(_003_),
    .Y(_118_));
 sky130_fd_sc_hd__o21ai_1 _367_ (.A1(_014_),
    .A2(_003_),
    .B1(_115_),
    .Y(_119_));
 sky130_fd_sc_hd__a21oi_1 _368_ (.A1(_012_),
    .A2(_062_),
    .B1(_068_),
    .Y(_120_));
 sky130_fd_sc_hd__a41o_1 _369_ (.A1(\dpath.a_lt_b$in0[3] ),
    .A2(_061_),
    .A3(_118_),
    .A4(_119_),
    .B1(_120_),
    .X(_121_));
 sky130_fd_sc_hd__nor2_1 _370_ (.A(_071_),
    .B(_011_),
    .Y(_122_));
 sky130_fd_sc_hd__or2_0 _371_ (.A(_122_),
    .B(_058_),
    .X(_123_));
 sky130_fd_sc_hd__o21ai_0 _372_ (.A1(net134),
    .A2(_057_),
    .B1(_071_),
    .Y(_124_));
 sky130_fd_sc_hd__a21boi_1 _373_ (.A1(net134),
    .A2(_057_),
    .B1_N(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__o31ai_4 _374_ (.A1(_117_),
    .A2(_123_),
    .A3(_121_),
    .B1(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__inv_1 _375_ (.A(\dpath.a_lt_b$in1[8] ),
    .Y(_127_));
 sky130_fd_sc_hd__maj3_2 _376_ (.A(net69),
    .B(_127_),
    .C(_085_),
    .X(_128_));
 sky130_fd_sc_hd__o21bai_2 _377_ (.A1(_046_),
    .A2(_128_),
    .B1_N(_044_),
    .Y(_129_));
 sky130_fd_sc_hd__a21oi_2 _378_ (.A1(_126_),
    .A2(_114_),
    .B1(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__xor2_1 _379_ (.A(net124),
    .B(_130_),
    .X(net39));
 sky130_fd_sc_hd__inv_1 _380_ (.A(\dpath.a_lt_b$in1[10] ),
    .Y(_131_));
 sky130_fd_sc_hd__nand3_1 _381_ (.A(_131_),
    .B(net93),
    .C(net91),
    .Y(_132_));
 sky130_fd_sc_hd__o21ai_4 _382_ (.A1(net39),
    .A2(_106_),
    .B1(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__nand2_1 _383_ (.A(net20),
    .B(_109_),
    .Y(_134_));
 sky130_fd_sc_hd__o21ai_1 _384_ (.A1(_109_),
    .A2(_133_),
    .B1(_134_),
    .Y(\dpath.a_mux$out[10] ));
 sky130_fd_sc_hd__maj3_2 _385_ (.A(_131_),
    .B(_130_),
    .C(net111),
    .X(_135_));
 sky130_fd_sc_hd__xnor2_2 _386_ (.A(_035_),
    .B(net64),
    .Y(net40));
 sky130_fd_sc_hd__nand2_4 _387_ (.A(_066_),
    .B(net90),
    .Y(_136_));
 sky130_fd_sc_hd__mux2i_1 _388_ (.A0(_009_),
    .A1(net40),
    .S(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(net21),
    .B(_109_),
    .Y(_138_));
 sky130_fd_sc_hd__o21ai_1 _390_ (.A1(_108_),
    .A2(_137_),
    .B1(_138_),
    .Y(\dpath.a_mux$out[11] ));
 sky130_fd_sc_hd__xor2_2 _391_ (.A(_008_),
    .B(\dpath.a_lt_b$in0[12] ),
    .X(_139_));
 sky130_fd_sc_hd__nand2b_1 _392_ (.A_N(\dpath.a_lt_b$in0[4] ),
    .B(\dpath.a_lt_b$in1[4] ),
    .Y(_140_));
 sky130_fd_sc_hd__nor3_1 _393_ (.A(_012_),
    .B(_057_),
    .C(_069_),
    .Y(_141_));
 sky130_fd_sc_hd__nand2_1 _394_ (.A(_062_),
    .B(net84),
    .Y(_142_));
 sky130_fd_sc_hd__a221o_1 _395_ (.A1(_121_),
    .A2(_140_),
    .B1(_142_),
    .B2(_141_),
    .C1(_058_),
    .X(_143_));
 sky130_fd_sc_hd__inv_1 _396_ (.A(net87),
    .Y(_144_));
 sky130_fd_sc_hd__maj3_1 _397_ (.A(_144_),
    .B(\dpath.a_lt_b$in0[6] ),
    .C(_122_),
    .X(_145_));
 sky130_fd_sc_hd__maj3_1 _398_ (.A(net107),
    .B(_083_),
    .C(_145_),
    .X(_146_));
 sky130_fd_sc_hd__a21oi_4 _399_ (.A1(_143_),
    .A2(net92),
    .B1(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__nor2b_1 _400_ (.A(_009_),
    .B_N(_034_),
    .Y(_148_));
 sky130_fd_sc_hd__maj3_1 _401_ (.A(_131_),
    .B(\dpath.a_lt_b$in0[10] ),
    .C(_113_),
    .X(_149_));
 sky130_fd_sc_hd__nand2b_1 _402_ (.A_N(_034_),
    .B(_009_),
    .Y(_150_));
 sky130_fd_sc_hd__o21ai_0 _403_ (.A1(_148_),
    .A2(_149_),
    .B1(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__nor2_1 _404_ (.A(_139_),
    .B(_035_),
    .Y(_152_));
 sky130_fd_sc_hd__nand2_1 _405_ (.A(net121),
    .B(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__nor2_2 _406_ (.A(_147_),
    .B(_153_),
    .Y(_154_));
 sky130_fd_sc_hd__a21oi_1 _407_ (.A1(net101),
    .A2(_037_),
    .B1(net120),
    .Y(_155_));
 sky130_fd_sc_hd__o2bb2ai_1 _408_ (.A1_N(_098_),
    .A2_N(_155_),
    .B1(_113_),
    .B2(_139_),
    .Y(_156_));
 sky130_fd_sc_hd__nand3_1 _409_ (.A(_034_),
    .B(_042_),
    .C(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__o21ai_0 _410_ (.A1(_139_),
    .A2(_096_),
    .B1(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__nand3_1 _411_ (.A(_095_),
    .B(net127),
    .C(_156_),
    .Y(_159_));
 sky130_fd_sc_hd__o21ai_0 _412_ (.A1(_009_),
    .A2(_041_),
    .B1(net120),
    .Y(_160_));
 sky130_fd_sc_hd__a21oi_1 _413_ (.A1(_159_),
    .A2(_160_),
    .B1(_034_),
    .Y(_161_));
 sky130_fd_sc_hd__a221oi_1 _414_ (.A1(_139_),
    .A2(_100_),
    .B1(_158_),
    .B2(_009_),
    .C1(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__a311oi_2 _415_ (.A1(_139_),
    .A2(net81),
    .A3(_151_),
    .B1(_154_),
    .C1(_162_),
    .Y(net41));
 sky130_fd_sc_hd__mux2i_1 _416_ (.A0(_008_),
    .A1(net79),
    .S(_136_),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_1 _417_ (.A(net22),
    .B(_109_),
    .Y(_164_));
 sky130_fd_sc_hd__o21ai_1 _418_ (.A1(_163_),
    .A2(_108_),
    .B1(_164_),
    .Y(\dpath.a_mux$out[12] ));
 sky130_fd_sc_hd__nand2_1 _419_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(_152_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _420_ (.A(_131_),
    .B(_152_),
    .Y(_166_));
 sky130_fd_sc_hd__a221oi_4 _421_ (.A1(_114_),
    .A2(net57),
    .B1(_165_),
    .B2(_166_),
    .C1(net55),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(net105),
    .B(_148_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _423_ (.A(_008_),
    .B(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o21ai_1 _424_ (.A1(net105),
    .A2(_148_),
    .B1(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(_040_),
    .B(_152_),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _426_ (.A(_170_),
    .B(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__o21ai_1 _427_ (.A1(_167_),
    .A2(_172_),
    .B1(\dpath.a_lt_b$in0[13] ),
    .Y(_173_));
 sky130_fd_sc_hd__or3_1 _428_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(_172_),
    .C(net74),
    .X(_174_));
 sky130_fd_sc_hd__a22oi_2 _429_ (.A1(net93),
    .A2(net217),
    .B1(_174_),
    .B2(_173_),
    .Y(_175_));
 sky130_fd_sc_hd__xnor2_1 _430_ (.A(_175_),
    .B(net122),
    .Y(_176_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(net23),
    .B(_109_),
    .Y(_177_));
 sky130_fd_sc_hd__o21ai_1 _432_ (.A1(_176_),
    .A2(_108_),
    .B1(_177_),
    .Y(\dpath.a_mux$out[13] ));
 sky130_fd_sc_hd__nor2b_1 _433_ (.A(net37),
    .B_N(\ctrl.state.out[2] ),
    .Y(_178_));
 sky130_fd_sc_hd__buf_2 _434_ (.A(_178_),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_4 _435_ (.A(_179_),
    .X(_180_));
 sky130_fd_sc_hd__nor2_1 _436_ (.A(_092_),
    .B(_016_),
    .Y(_181_));
 sky130_fd_sc_hd__a2111oi_2 _437_ (.A1(_089_),
    .A2(net105),
    .B1(_181_),
    .C1(_148_),
    .D1(_149_),
    .Y(_182_));
 sky130_fd_sc_hd__a211oi_1 _438_ (.A1(_089_),
    .A2(net105),
    .B1(_181_),
    .C1(_150_),
    .Y(_183_));
 sky130_fd_sc_hd__a211oi_1 _439_ (.A1(_090_),
    .A2(_030_),
    .B1(_182_),
    .C1(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__nand3_1 _440_ (.A(_031_),
    .B(_048_),
    .C(_152_),
    .Y(_185_));
 sky130_fd_sc_hd__o2bb2ai_2 _441_ (.A1_N(net227),
    .A2_N(_184_),
    .B1(_185_),
    .B2(net80),
    .Y(_186_));
 sky130_fd_sc_hd__xor2_1 _442_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(_186_),
    .X(_187_));
 sky130_fd_sc_hd__o21ai_0 _443_ (.A1(_106_),
    .A2(_187_),
    .B1(\dpath.a_lt_b$in1[14] ),
    .Y(_188_));
 sky130_fd_sc_hd__or3_1 _444_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(_105_),
    .C(_187_),
    .X(_189_));
 sky130_fd_sc_hd__nor2_1 _445_ (.A(net25),
    .B(_180_),
    .Y(_190_));
 sky130_fd_sc_hd__a31oi_1 _446_ (.A1(_189_),
    .A2(_188_),
    .A3(_180_),
    .B1(_190_),
    .Y(\dpath.a_mux$out[14] ));
 sky130_fd_sc_hd__nand2_1 _447_ (.A(net26),
    .B(_109_),
    .Y(_191_));
 sky130_fd_sc_hd__maj3_1 _448_ (.A(_092_),
    .B(net122),
    .C(_170_),
    .X(_192_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(_029_),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__a22oi_4 _450_ (.A1(_135_),
    .A2(net95),
    .B1(_193_),
    .B2(_028_),
    .Y(_194_));
 sky130_fd_sc_hd__or3_1 _451_ (.A(_049_),
    .B(_108_),
    .C(_194_),
    .X(_195_));
 sky130_fd_sc_hd__nand3_1 _452_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(_106_),
    .C(_180_),
    .Y(_196_));
 sky130_fd_sc_hd__nand3_1 _453_ (.A(_191_),
    .B(_195_),
    .C(_196_),
    .Y(\dpath.a_mux$out[15] ));
 sky130_fd_sc_hd__nand2_1 _454_ (.A(_014_),
    .B(net137),
    .Y(_197_));
 sky130_fd_sc_hd__xnor2_1 _455_ (.A(_003_),
    .B(_065_),
    .Y(net45));
 sky130_fd_sc_hd__nand2_1 _456_ (.A(_136_),
    .B(net45),
    .Y(_198_));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(net10),
    .B(_179_),
    .Y(_199_));
 sky130_fd_sc_hd__a31oi_1 _458_ (.A1(_180_),
    .A2(_197_),
    .A3(_198_),
    .B1(_199_),
    .Y(\dpath.a_mux$out[1] ));
 sky130_fd_sc_hd__nand2_1 _459_ (.A(net307),
    .B(_106_),
    .Y(_200_));
 sky130_fd_sc_hd__xnor2_1 _460_ (.A(_063_),
    .B(net66),
    .Y(net46));
 sky130_fd_sc_hd__nand2_1 _461_ (.A(_136_),
    .B(net46),
    .Y(_201_));
 sky130_fd_sc_hd__nor2_1 _462_ (.A(net11),
    .B(_179_),
    .Y(_202_));
 sky130_fd_sc_hd__a31oi_1 _463_ (.A1(_180_),
    .A2(_201_),
    .A3(_200_),
    .B1(_202_),
    .Y(\dpath.a_mux$out[2] ));
 sky130_fd_sc_hd__nand2_1 _464_ (.A(_012_),
    .B(net137),
    .Y(_203_));
 sky130_fd_sc_hd__nand2_1 _465_ (.A(_061_),
    .B(_142_),
    .Y(_204_));
 sky130_fd_sc_hd__xnor2_1 _466_ (.A(_060_),
    .B(_204_),
    .Y(net47));
 sky130_fd_sc_hd__nand2_1 _467_ (.A(_136_),
    .B(net47),
    .Y(_205_));
 sky130_fd_sc_hd__nor2_1 _468_ (.A(net12),
    .B(_179_),
    .Y(_206_));
 sky130_fd_sc_hd__a31oi_1 _469_ (.A1(_180_),
    .A2(_203_),
    .A3(_205_),
    .B1(_206_),
    .Y(\dpath.a_mux$out[3] ));
 sky130_fd_sc_hd__nand2_1 _470_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(net137),
    .Y(_207_));
 sky130_fd_sc_hd__nor2_2 _471_ (.A(net72),
    .B(net58),
    .Y(_208_));
 sky130_fd_sc_hd__xnor2_1 _472_ (.A(_208_),
    .B(_059_),
    .Y(net48));
 sky130_fd_sc_hd__nand2_1 _473_ (.A(_136_),
    .B(net48),
    .Y(_209_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(net14),
    .B(_179_),
    .Y(_210_));
 sky130_fd_sc_hd__a31oi_1 _475_ (.A1(_180_),
    .A2(_207_),
    .A3(_209_),
    .B1(_210_),
    .Y(\dpath.a_mux$out[4] ));
 sky130_fd_sc_hd__nand2_1 _476_ (.A(_011_),
    .B(net137),
    .Y(_211_));
 sky130_fd_sc_hd__xnor2_2 _477_ (.A(_055_),
    .B(_143_),
    .Y(net49));
 sky130_fd_sc_hd__nand2_1 _478_ (.A(_136_),
    .B(net49),
    .Y(_212_));
 sky130_fd_sc_hd__nor2_1 _479_ (.A(net15),
    .B(_179_),
    .Y(_213_));
 sky130_fd_sc_hd__a31oi_1 _480_ (.A1(_180_),
    .A2(_212_),
    .A3(_211_),
    .B1(_213_),
    .Y(\dpath.a_mux$out[5] ));
 sky130_fd_sc_hd__nand2_1 _481_ (.A(net88),
    .B(net137),
    .Y(_214_));
 sky130_fd_sc_hd__nor2_1 _482_ (.A(_053_),
    .B(_054_),
    .Y(_215_));
 sky130_fd_sc_hd__xnor2_1 _483_ (.A(_215_),
    .B(_126_),
    .Y(net50));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(_136_),
    .B(net50),
    .Y(_216_));
 sky130_fd_sc_hd__nor2_1 _485_ (.A(net16),
    .B(_179_),
    .Y(_217_));
 sky130_fd_sc_hd__a31oi_1 _486_ (.A1(_180_),
    .A2(_214_),
    .A3(_216_),
    .B1(_217_),
    .Y(\dpath.a_mux$out[6] ));
 sky130_fd_sc_hd__nand2_1 _487_ (.A(_144_),
    .B(net85),
    .Y(_218_));
 sky130_fd_sc_hd__a21oi_2 _488_ (.A1(_218_),
    .A2(net56),
    .B1(_053_),
    .Y(_219_));
 sky130_fd_sc_hd__xor2_2 _489_ (.A(net108),
    .B(net67),
    .X(_220_));
 sky130_fd_sc_hd__a21oi_2 _490_ (.A1(net94),
    .A2(net91),
    .B1(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__xnor2_1 _491_ (.A(_221_),
    .B(net116),
    .Y(_222_));
 sky130_fd_sc_hd__nand2_1 _492_ (.A(net17),
    .B(_109_),
    .Y(_223_));
 sky130_fd_sc_hd__o21ai_1 _493_ (.A1(_108_),
    .A2(_222_),
    .B1(_223_),
    .Y(\dpath.a_mux$out[7] ));
 sky130_fd_sc_hd__xnor2_2 _494_ (.A(net71),
    .B(net216),
    .Y(_224_));
 sky130_fd_sc_hd__a21oi_2 _495_ (.A1(net94),
    .A2(net91),
    .B1(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_1 _496_ (.A(net313),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(net18),
    .B(_109_),
    .Y(_227_));
 sky130_fd_sc_hd__o21ai_1 _498_ (.A1(_108_),
    .A2(_226_),
    .B1(_227_),
    .Y(\dpath.a_mux$out[8] ));
 sky130_fd_sc_hd__inv_1 _499_ (.A(net70),
    .Y(_228_));
 sky130_fd_sc_hd__maj3_2 _500_ (.A(_147_),
    .B(net310),
    .C(_228_),
    .X(_229_));
 sky130_fd_sc_hd__xnor2_2 _501_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(net82),
    .Y(_230_));
 sky130_fd_sc_hd__o21ai_0 _502_ (.A1(_105_),
    .A2(_230_),
    .B1(net98),
    .Y(_231_));
 sky130_fd_sc_hd__or3_1 _503_ (.A(net97),
    .B(_105_),
    .C(_230_),
    .X(_232_));
 sky130_fd_sc_hd__nor2_1 _504_ (.A(net19),
    .B(_179_),
    .Y(_233_));
 sky130_fd_sc_hd__a31oi_1 _505_ (.A1(_232_),
    .A2(_180_),
    .A3(_231_),
    .B1(_233_),
    .Y(\dpath.a_mux$out[9] ));
 sky130_fd_sc_hd__mux2_1 _506_ (.A0(net62),
    .A1(net2),
    .S(_006_),
    .X(\dpath.b_mux$out[0] ));
 sky130_fd_sc_hd__mux2_1 _507_ (.A0(\dpath.a_lt_b$in0[10] ),
    .A1(net3),
    .S(_006_),
    .X(\dpath.b_mux$out[10] ));
 sky130_fd_sc_hd__mux2_1 _508_ (.A0(_034_),
    .A1(net4),
    .S(_005_),
    .X(\dpath.b_mux$out[11] ));
 sky130_fd_sc_hd__mux2_1 _509_ (.A0(net106),
    .A1(net5),
    .S(_005_),
    .X(\dpath.b_mux$out[12] ));
 sky130_fd_sc_hd__nand2_1 _510_ (.A(_107_),
    .B(net6),
    .Y(_234_));
 sky130_fd_sc_hd__o21ai_0 _511_ (.A1(_107_),
    .A2(_092_),
    .B1(_234_),
    .Y(\dpath.b_mux$out[13] ));
 sky130_fd_sc_hd__mux2_1 _512_ (.A0(\dpath.a_lt_b$in0[14] ),
    .A1(net7),
    .S(_005_),
    .X(\dpath.b_mux$out[14] ));
 sky130_fd_sc_hd__nand2_1 _513_ (.A(_107_),
    .B(net8),
    .Y(_235_));
 sky130_fd_sc_hd__o21ai_0 _514_ (.A1(_107_),
    .A2(_088_),
    .B1(_235_),
    .Y(\dpath.b_mux$out[15] ));
 sky130_fd_sc_hd__nand2_1 _515_ (.A(_107_),
    .B(net13),
    .Y(_236_));
 sky130_fd_sc_hd__o21ai_0 _516_ (.A1(_006_),
    .A2(_115_),
    .B1(_236_),
    .Y(\dpath.b_mux$out[1] ));
 sky130_fd_sc_hd__mux2_1 _517_ (.A0(\dpath.a_lt_b$in0[2] ),
    .A1(net24),
    .S(_005_),
    .X(\dpath.b_mux$out[2] ));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(_107_),
    .B(net27),
    .Y(_237_));
 sky130_fd_sc_hd__o21ai_0 _519_ (.A1(_006_),
    .A2(_068_),
    .B1(_237_),
    .Y(\dpath.b_mux$out[3] ));
 sky130_fd_sc_hd__mux2_1 _520_ (.A0(\dpath.a_lt_b$in0[4] ),
    .A1(net28),
    .S(_005_),
    .X(\dpath.b_mux$out[4] ));
 sky130_fd_sc_hd__nand2_1 _521_ (.A(_107_),
    .B(net29),
    .Y(_238_));
 sky130_fd_sc_hd__o21ai_0 _522_ (.A1(_006_),
    .A2(_071_),
    .B1(_238_),
    .Y(\dpath.b_mux$out[5] ));
 sky130_fd_sc_hd__mux2_1 _523_ (.A0(\dpath.a_lt_b$in0[6] ),
    .A1(net30),
    .S(_005_),
    .X(\dpath.b_mux$out[6] ));
 sky130_fd_sc_hd__mux2_1 _524_ (.A0(_051_),
    .A1(net31),
    .S(_005_),
    .X(\dpath.b_mux$out[7] ));
 sky130_fd_sc_hd__nand2_1 _525_ (.A(_107_),
    .B(net32),
    .Y(_239_));
 sky130_fd_sc_hd__o21ai_0 _526_ (.A1(_006_),
    .A2(_228_),
    .B1(_239_),
    .Y(\dpath.b_mux$out[8] ));
 sky130_fd_sc_hd__nand2_1 _527_ (.A(_107_),
    .B(net33),
    .Y(_240_));
 sky130_fd_sc_hd__o21ai_0 _528_ (.A1(_006_),
    .A2(net129),
    .B1(_240_),
    .Y(\dpath.b_mux$out[9] ));
 sky130_fd_sc_hd__nor2_2 _529_ (.A(_167_),
    .B(_172_),
    .Y(_241_));
 sky130_fd_sc_hd__xnor2_1 _530_ (.A(_241_),
    .B(net126),
    .Y(net42));
 sky130_fd_sc_hd__nand2_1 _531_ (.A(_028_),
    .B(_029_),
    .Y(_242_));
 sky130_fd_sc_hd__xnor2_1 _532_ (.A(_242_),
    .B(_186_),
    .Y(net43));
 sky130_fd_sc_hd__xnor2_2 _533_ (.A(_049_),
    .B(_194_),
    .Y(net44));
 sky130_fd_sc_hd__xnor2_1 _534_ (.A(_052_),
    .B(_219_),
    .Y(net51));
 sky130_fd_sc_hd__xnor2_1 _535_ (.A(net76),
    .B(net314),
    .Y(net52));
 sky130_fd_sc_hd__xnor2_2 _536_ (.A(_047_),
    .B(_229_),
    .Y(net53));
 sky130_fd_sc_hd__dfxtp_1 \ctrl.state.out[0]$_DFF_P_  (.D(_000_),
    .Q(net37),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \ctrl.state.out[1]$_DFF_P_  (.D(_001_),
    .Q(\ctrl.state.out[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \ctrl.state.out[2]$_DFF_P_  (.D(_002_),
    .Q(\ctrl.state.out[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[0]$_DFFE_PP_  (.D(\dpath.a_mux$out[0] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[0] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[10]$_DFFE_PP_  (.D(\dpath.a_mux$out[10] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[10] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[11]$_DFFE_PP_  (.D(\dpath.a_mux$out[11] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[11] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[12]$_DFFE_PP_  (.D(\dpath.a_mux$out[12] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[12] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[13]$_DFFE_PP_  (.D(\dpath.a_mux$out[13] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[13] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[14]$_DFFE_PP_  (.D(\dpath.a_mux$out[14] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[14] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[15]$_DFFE_PP_  (.D(\dpath.a_mux$out[15] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[15] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[1]$_DFFE_PP_  (.D(\dpath.a_mux$out[1] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[1] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[2]$_DFFE_PP_  (.D(\dpath.a_mux$out[2] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[3]$_DFFE_PP_  (.D(\dpath.a_mux$out[3] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[4]$_DFFE_PP_  (.D(\dpath.a_mux$out[4] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[4] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[5]$_DFFE_PP_  (.D(\dpath.a_mux$out[5] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[5] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[6]$_DFFE_PP_  (.D(\dpath.a_mux$out[6] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[6] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[7]$_DFFE_PP_  (.D(\dpath.a_mux$out[7] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[7] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[8]$_DFFE_PP_  (.D(\dpath.a_mux$out[8] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[8] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.a_reg.out[9]$_DFFE_PP_  (.D(\dpath.a_mux$out[9] ),
    .DE(\ctrl$a_reg_en ),
    .Q(\dpath.a_lt_b$in0[9] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[0]$_DFFE_PP_  (.D(\dpath.b_mux$out[0] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[0] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[10]$_DFFE_PP_  (.D(\dpath.b_mux$out[10] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[10] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[11]$_DFFE_PP_  (.D(\dpath.b_mux$out[11] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[11] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[12]$_DFFE_PP_  (.D(\dpath.b_mux$out[12] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[12] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[13]$_DFFE_PP_  (.D(\dpath.b_mux$out[13] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[13] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[14]$_DFFE_PP_  (.D(\dpath.b_mux$out[14] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[14] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[15]$_DFFE_PP_  (.D(\dpath.b_mux$out[15] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[15] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[1]$_DFFE_PP_  (.D(\dpath.b_mux$out[1] ),
    .DE(net1),
    .Q(\dpath.a_lt_b$in1[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[2]$_DFFE_PP_  (.D(\dpath.b_mux$out[2] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[3]$_DFFE_PP_  (.D(\dpath.b_mux$out[3] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[4]$_DFFE_PP_  (.D(\dpath.b_mux$out[4] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[4] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[5]$_DFFE_PP_  (.D(\dpath.b_mux$out[5] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[5] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[6]$_DFFE_PP_  (.D(\dpath.b_mux$out[6] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[6] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[7]$_DFFE_PP_  (.D(\dpath.b_mux$out[7] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[7] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[8]$_DFFE_PP_  (.D(\dpath.b_mux$out[8] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[8] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dpath.b_reg.out[9]$_DFFE_PP_  (.D(\dpath.b_mux$out[9] ),
    .DE(\ctrl$b_reg_en ),
    .Q(\dpath.a_lt_b$in1[9] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_95 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(req_msg[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(req_msg[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(req_msg[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(req_msg[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(req_msg[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(req_msg[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(req_msg[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(req_msg[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(req_msg[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(req_msg[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(req_msg[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(req_msg[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(req_msg[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(req_msg[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(req_msg[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(req_msg[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(req_msg[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(req_msg[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(req_msg[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(req_msg[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(req_msg[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(req_msg[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(req_msg[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(req_msg[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(req_msg[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(req_msg[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(req_msg[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(req_msg[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(req_msg[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(req_msg[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(req_msg[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(req_msg[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(req_val),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(reset),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(resp_rdy),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(req_rdy));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(resp_msg[0]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(resp_msg[10]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(resp_msg[11]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(resp_msg[12]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(resp_msg[13]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(resp_msg[14]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(resp_msg[15]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(resp_msg[1]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(resp_msg[2]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(resp_msg[3]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(resp_msg[4]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(resp_msg[5]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(resp_msg[6]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(resp_msg[7]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net52),
    .X(resp_msg[8]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net53),
    .X(resp_msg[9]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net54),
    .X(resp_val));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 rebuffer1 (.A(_129_),
    .X(net55));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(_126_),
    .X(net56));
 sky130_fd_sc_hd__buf_2 rebuffer3 (.A(_126_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 rebuffer4 (.A(_117_),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net78),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(\dpath.a_lt_b$in0[0] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(\dpath.a_lt_b$in0[0] ),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer8 (.A(net61),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(\dpath.a_lt_b$in0[6] ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 rebuffer10 (.A(_135_),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer32 (.A(_039_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(_116_),
    .X(net66));
 sky130_fd_sc_hd__buf_2 rebuffer13 (.A(_219_),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(_085_),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(\dpath.a_lt_b$in0[8] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net69),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net69),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(_121_),
    .X(net72));
 sky130_fd_sc_hd__buf_6 rebuffer65 (.A(_036_),
    .X(net119));
 sky130_fd_sc_hd__buf_1 rebuffer20 (.A(_167_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(\dpath.a_lt_b$in1[0] ),
    .X(net75));
 sky130_fd_sc_hd__buf_2 rebuffer26 (.A(_147_),
    .X(net80));
 sky130_fd_sc_hd__buf_2 rebuffer27 (.A(_147_),
    .X(net81));
 sky130_fd_sc_hd__buf_6 rebuffer28 (.A(_229_),
    .X(net82));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer80 (.A(_011_),
    .X(net134));
 sky130_fd_sc_hd__buf_1 rebuffer30 (.A(_116_),
    .X(net84));
 sky130_fd_sc_hd__buf_6 rebuffer33 (.A(\dpath.a_lt_b$in1[6] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net87),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net87),
    .X(net89));
 sky130_fd_sc_hd__buf_2 rebuffer36 (.A(_104_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 rebuffer37 (.A(_104_),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(_056_),
    .X(net92));
 sky130_fd_sc_hd__buf_6 rebuffer39 (.A(_066_),
    .X(net93));
 sky130_fd_sc_hd__buf_6 rebuffer40 (.A(_066_),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net103),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(\dpath.a_lt_b$in1[9] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net96),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net97),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 rebuffer45 (.A(\dpath.a_lt_b$in1[9] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(\dpath.a_lt_b$in1[9] ),
    .X(net100));
 sky130_fd_sc_hd__buf_1 rebuffer47 (.A(net100),
    .X(net101));
 sky130_fd_sc_hd__buf_2 rebuffer48 (.A(net101),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(_036_),
    .X(net103));
 sky130_fd_sc_hd__buf_1 rebuffer50 (.A(_064_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 rebuffer51 (.A(\dpath.a_lt_b$in0[12] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net105),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(_051_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(_051_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer173 (.A(_031_),
    .X(net227));
 sky130_fd_sc_hd__buf_6 rebuffer56 (.A(\dpath.a_lt_b$in1[7] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(\dpath.a_lt_b$in0[10] ),
    .X(net111));
 sky130_fd_sc_hd__buf_2 rebuffer58 (.A(\dpath.a_lt_b$in0[10] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer163 (.A(_104_),
    .X(net217));
 sky130_fd_sc_hd__buf_2 rebuffer162 (.A(_147_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer161 (.A(_013_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net136),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer253 (.A(\dpath.a_lt_b$in1[2] ),
    .X(net307));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer254 (.A(\dpath.a_lt_b$in1[2] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer255 (.A(net308),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer256 (.A(\dpath.a_lt_b$in1[8] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer257 (.A(net310),
    .X(net311));
 sky130_fd_sc_hd__buf_2 rebuffer258 (.A(\dpath.a_lt_b$in1[8] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer259 (.A(net312),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer260 (.A(net86),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(_147_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(\dpath.a_lt_b$in1[0] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(\dpath.a_lt_b$in1[0] ),
    .X(net78));
 sky130_fd_sc_hd__buf_2 rebuffer25 (.A(net41),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(\dpath.a_lt_b$in0[6] ),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer66 (.A(_027_),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer67 (.A(_048_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(_016_),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(_016_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(_042_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(\dpath.a_lt_b$in1[10] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer72 (.A(_032_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer73 (.A(_042_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer74 (.A(_045_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer75 (.A(_045_),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer81 (.A(net134),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer82 (.A(\dpath.a_lt_b$in1[7] ),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_16 clone83 (.A(_105_),
    .X(net137));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
endmodule
