module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire \dcnt[0] ;
 wire \dcnt[1] ;
 wire \dcnt[2] ;
 wire \dcnt[3] ;
 wire ld_r;
 wire \sa00_sr[0] ;
 wire \sa00_sr[1] ;
 wire \sa00_sr[2] ;
 wire \sa00_sr[3] ;
 wire \sa00_sr[4] ;
 wire \sa00_sr[5] ;
 wire \sa00_sr[6] ;
 wire \sa00_sr[7] ;
 wire \sa01_sr[0] ;
 wire \sa01_sr[1] ;
 wire \sa01_sr[2] ;
 wire \sa01_sr[3] ;
 wire \sa01_sr[4] ;
 wire \sa01_sr[5] ;
 wire \sa01_sr[6] ;
 wire \sa01_sr[7] ;
 wire \sa02_sr[0] ;
 wire \sa02_sr[1] ;
 wire \sa02_sr[2] ;
 wire \sa02_sr[3] ;
 wire \sa02_sr[4] ;
 wire \sa02_sr[5] ;
 wire \sa02_sr[6] ;
 wire \sa02_sr[7] ;
 wire \sa03_sr[0] ;
 wire \sa03_sr[1] ;
 wire \sa03_sr[2] ;
 wire \sa03_sr[3] ;
 wire \sa03_sr[4] ;
 wire \sa03_sr[5] ;
 wire \sa03_sr[6] ;
 wire \sa03_sr[7] ;
 wire \sa10_sr[0] ;
 wire \sa10_sr[1] ;
 wire \sa10_sr[2] ;
 wire \sa10_sr[3] ;
 wire \sa10_sr[4] ;
 wire \sa10_sr[5] ;
 wire \sa10_sr[6] ;
 wire \sa10_sr[7] ;
 wire \sa10_sub[0] ;
 wire \sa10_sub[1] ;
 wire \sa10_sub[2] ;
 wire \sa10_sub[3] ;
 wire \sa10_sub[4] ;
 wire \sa10_sub[5] ;
 wire \sa10_sub[6] ;
 wire \sa10_sub[7] ;
 wire \sa11_sr[0] ;
 wire \sa11_sr[1] ;
 wire \sa11_sr[2] ;
 wire \sa11_sr[3] ;
 wire \sa11_sr[4] ;
 wire \sa11_sr[5] ;
 wire \sa11_sr[6] ;
 wire \sa11_sr[7] ;
 wire \sa12_sr[0] ;
 wire \sa12_sr[1] ;
 wire \sa12_sr[2] ;
 wire \sa12_sr[3] ;
 wire \sa12_sr[4] ;
 wire \sa12_sr[5] ;
 wire \sa12_sr[6] ;
 wire \sa12_sr[7] ;
 wire \sa20_sr[0] ;
 wire \sa20_sr[1] ;
 wire \sa20_sr[2] ;
 wire \sa20_sr[3] ;
 wire \sa20_sr[4] ;
 wire \sa20_sr[5] ;
 wire \sa20_sr[6] ;
 wire \sa20_sr[7] ;
 wire \sa20_sub[0] ;
 wire \sa20_sub[1] ;
 wire \sa20_sub[2] ;
 wire \sa20_sub[3] ;
 wire \sa20_sub[4] ;
 wire \sa20_sub[5] ;
 wire \sa20_sub[6] ;
 wire \sa20_sub[7] ;
 wire \sa21_sr[0] ;
 wire \sa21_sr[1] ;
 wire \sa21_sr[2] ;
 wire \sa21_sr[3] ;
 wire \sa21_sr[4] ;
 wire \sa21_sr[5] ;
 wire \sa21_sr[6] ;
 wire \sa21_sr[7] ;
 wire \sa21_sub[0] ;
 wire \sa21_sub[1] ;
 wire \sa21_sub[2] ;
 wire \sa21_sub[3] ;
 wire \sa21_sub[4] ;
 wire \sa21_sub[5] ;
 wire \sa21_sub[6] ;
 wire \sa21_sub[7] ;
 wire \sa30_sr[0] ;
 wire \sa30_sr[1] ;
 wire \sa30_sr[2] ;
 wire \sa30_sr[3] ;
 wire \sa30_sr[4] ;
 wire \sa30_sr[5] ;
 wire \sa30_sr[6] ;
 wire \sa30_sr[7] ;
 wire \sa30_sub[0] ;
 wire \sa30_sub[1] ;
 wire \sa30_sub[2] ;
 wire \sa30_sub[3] ;
 wire \sa30_sub[4] ;
 wire \sa30_sub[5] ;
 wire \sa30_sub[6] ;
 wire \sa30_sub[7] ;
 wire \sa31_sub[0] ;
 wire \sa31_sub[1] ;
 wire \sa31_sub[2] ;
 wire \sa31_sub[3] ;
 wire \sa31_sub[4] ;
 wire \sa31_sub[5] ;
 wire \sa31_sub[6] ;
 wire \sa31_sub[7] ;
 wire \sa32_sub[0] ;
 wire \sa32_sub[1] ;
 wire \sa32_sub[2] ;
 wire \sa32_sub[3] ;
 wire \sa32_sub[4] ;
 wire \sa32_sub[5] ;
 wire \sa32_sub[6] ;
 wire \sa32_sub[7] ;
 wire \text_in_r[0] ;
 wire \text_in_r[100] ;
 wire \text_in_r[101] ;
 wire \text_in_r[102] ;
 wire \text_in_r[103] ;
 wire \text_in_r[104] ;
 wire \text_in_r[105] ;
 wire \text_in_r[106] ;
 wire \text_in_r[107] ;
 wire \text_in_r[108] ;
 wire \text_in_r[109] ;
 wire \text_in_r[10] ;
 wire \text_in_r[110] ;
 wire \text_in_r[111] ;
 wire \text_in_r[112] ;
 wire \text_in_r[113] ;
 wire \text_in_r[114] ;
 wire \text_in_r[115] ;
 wire \text_in_r[116] ;
 wire \text_in_r[117] ;
 wire \text_in_r[118] ;
 wire \text_in_r[119] ;
 wire \text_in_r[11] ;
 wire \text_in_r[120] ;
 wire \text_in_r[121] ;
 wire \text_in_r[122] ;
 wire \text_in_r[123] ;
 wire \text_in_r[124] ;
 wire \text_in_r[125] ;
 wire \text_in_r[126] ;
 wire \text_in_r[127] ;
 wire \text_in_r[12] ;
 wire \text_in_r[13] ;
 wire \text_in_r[14] ;
 wire \text_in_r[15] ;
 wire \text_in_r[16] ;
 wire \text_in_r[17] ;
 wire \text_in_r[18] ;
 wire \text_in_r[19] ;
 wire \text_in_r[1] ;
 wire \text_in_r[20] ;
 wire \text_in_r[21] ;
 wire \text_in_r[22] ;
 wire \text_in_r[23] ;
 wire \text_in_r[24] ;
 wire \text_in_r[25] ;
 wire \text_in_r[26] ;
 wire \text_in_r[27] ;
 wire \text_in_r[28] ;
 wire \text_in_r[29] ;
 wire \text_in_r[2] ;
 wire \text_in_r[30] ;
 wire \text_in_r[31] ;
 wire \text_in_r[32] ;
 wire \text_in_r[33] ;
 wire \text_in_r[34] ;
 wire \text_in_r[35] ;
 wire \text_in_r[36] ;
 wire \text_in_r[37] ;
 wire \text_in_r[38] ;
 wire \text_in_r[39] ;
 wire \text_in_r[3] ;
 wire \text_in_r[40] ;
 wire \text_in_r[41] ;
 wire \text_in_r[42] ;
 wire \text_in_r[43] ;
 wire \text_in_r[44] ;
 wire \text_in_r[45] ;
 wire \text_in_r[46] ;
 wire \text_in_r[47] ;
 wire \text_in_r[48] ;
 wire \text_in_r[49] ;
 wire \text_in_r[4] ;
 wire \text_in_r[50] ;
 wire \text_in_r[51] ;
 wire \text_in_r[52] ;
 wire \text_in_r[53] ;
 wire \text_in_r[54] ;
 wire \text_in_r[55] ;
 wire \text_in_r[56] ;
 wire \text_in_r[57] ;
 wire \text_in_r[58] ;
 wire \text_in_r[59] ;
 wire \text_in_r[5] ;
 wire \text_in_r[60] ;
 wire \text_in_r[61] ;
 wire \text_in_r[62] ;
 wire \text_in_r[63] ;
 wire \text_in_r[64] ;
 wire \text_in_r[65] ;
 wire \text_in_r[66] ;
 wire \text_in_r[67] ;
 wire \text_in_r[68] ;
 wire \text_in_r[69] ;
 wire \text_in_r[6] ;
 wire \text_in_r[70] ;
 wire \text_in_r[71] ;
 wire \text_in_r[72] ;
 wire \text_in_r[73] ;
 wire \text_in_r[74] ;
 wire \text_in_r[75] ;
 wire \text_in_r[76] ;
 wire \text_in_r[77] ;
 wire \text_in_r[78] ;
 wire \text_in_r[79] ;
 wire \text_in_r[7] ;
 wire \text_in_r[80] ;
 wire \text_in_r[81] ;
 wire \text_in_r[82] ;
 wire \text_in_r[83] ;
 wire \text_in_r[84] ;
 wire \text_in_r[85] ;
 wire \text_in_r[86] ;
 wire \text_in_r[87] ;
 wire \text_in_r[88] ;
 wire \text_in_r[89] ;
 wire \text_in_r[8] ;
 wire \text_in_r[90] ;
 wire \text_in_r[91] ;
 wire \text_in_r[92] ;
 wire \text_in_r[93] ;
 wire \text_in_r[94] ;
 wire \text_in_r[95] ;
 wire \text_in_r[96] ;
 wire \text_in_r[97] ;
 wire \text_in_r[98] ;
 wire \text_in_r[99] ;
 wire \text_in_r[9] ;
 wire \u0.r0.out[24] ;
 wire \u0.r0.out[25] ;
 wire \u0.r0.out[26] ;
 wire \u0.r0.out[27] ;
 wire \u0.r0.out[28] ;
 wire \u0.r0.out[29] ;
 wire \u0.r0.out[30] ;
 wire \u0.r0.out[31] ;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt[2] ;
 wire \u0.r0.rcnt[3] ;
 wire \u0.r0.rcnt_next[0] ;
 wire \u0.r0.rcnt_next[1] ;
 wire \u0.subword[0] ;
 wire \u0.subword[10] ;
 wire \u0.subword[11] ;
 wire \u0.subword[12] ;
 wire \u0.subword[13] ;
 wire \u0.subword[14] ;
 wire \u0.subword[15] ;
 wire \u0.subword[16] ;
 wire \u0.subword[17] ;
 wire \u0.subword[18] ;
 wire \u0.subword[19] ;
 wire \u0.subword[1] ;
 wire \u0.subword[20] ;
 wire \u0.subword[21] ;
 wire \u0.subword[22] ;
 wire \u0.subword[23] ;
 wire \u0.subword[24] ;
 wire \u0.subword[25] ;
 wire \u0.subword[26] ;
 wire \u0.subword[27] ;
 wire \u0.subword[28] ;
 wire \u0.subword[29] ;
 wire \u0.subword[2] ;
 wire \u0.subword[30] ;
 wire \u0.subword[31] ;
 wire \u0.subword[3] ;
 wire \u0.subword[4] ;
 wire \u0.subword[5] ;
 wire \u0.subword[6] ;
 wire \u0.subword[7] ;
 wire \u0.subword[8] ;
 wire \u0.subword[9] ;
 wire \u0.tmp_w[0] ;
 wire \u0.tmp_w[10] ;
 wire \u0.tmp_w[11] ;
 wire \u0.tmp_w[12] ;
 wire \u0.tmp_w[13] ;
 wire \u0.tmp_w[14] ;
 wire \u0.tmp_w[15] ;
 wire \u0.tmp_w[16] ;
 wire \u0.tmp_w[17] ;
 wire \u0.tmp_w[18] ;
 wire \u0.tmp_w[19] ;
 wire \u0.tmp_w[1] ;
 wire \u0.tmp_w[20] ;
 wire \u0.tmp_w[21] ;
 wire \u0.tmp_w[22] ;
 wire \u0.tmp_w[23] ;
 wire \u0.tmp_w[24] ;
 wire \u0.tmp_w[25] ;
 wire \u0.tmp_w[26] ;
 wire \u0.tmp_w[27] ;
 wire \u0.tmp_w[28] ;
 wire \u0.tmp_w[29] ;
 wire \u0.tmp_w[2] ;
 wire \u0.tmp_w[30] ;
 wire \u0.tmp_w[31] ;
 wire \u0.tmp_w[3] ;
 wire \u0.tmp_w[4] ;
 wire \u0.tmp_w[5] ;
 wire \u0.tmp_w[6] ;
 wire \u0.tmp_w[7] ;
 wire \u0.tmp_w[8] ;
 wire \u0.tmp_w[9] ;
 wire \u0.w[0][0] ;
 wire \u0.w[0][10] ;
 wire \u0.w[0][11] ;
 wire \u0.w[0][12] ;
 wire \u0.w[0][13] ;
 wire \u0.w[0][14] ;
 wire \u0.w[0][15] ;
 wire \u0.w[0][16] ;
 wire \u0.w[0][17] ;
 wire \u0.w[0][18] ;
 wire \u0.w[0][19] ;
 wire \u0.w[0][1] ;
 wire \u0.w[0][20] ;
 wire \u0.w[0][21] ;
 wire \u0.w[0][22] ;
 wire \u0.w[0][23] ;
 wire \u0.w[0][24] ;
 wire \u0.w[0][25] ;
 wire \u0.w[0][26] ;
 wire \u0.w[0][27] ;
 wire \u0.w[0][28] ;
 wire \u0.w[0][29] ;
 wire \u0.w[0][2] ;
 wire \u0.w[0][30] ;
 wire \u0.w[0][31] ;
 wire \u0.w[0][3] ;
 wire \u0.w[0][4] ;
 wire \u0.w[0][5] ;
 wire \u0.w[0][6] ;
 wire \u0.w[0][7] ;
 wire \u0.w[0][8] ;
 wire \u0.w[0][9] ;
 wire \u0.w[1][0] ;
 wire \u0.w[1][10] ;
 wire \u0.w[1][11] ;
 wire \u0.w[1][12] ;
 wire \u0.w[1][13] ;
 wire \u0.w[1][14] ;
 wire \u0.w[1][15] ;
 wire \u0.w[1][16] ;
 wire \u0.w[1][17] ;
 wire \u0.w[1][18] ;
 wire \u0.w[1][19] ;
 wire \u0.w[1][1] ;
 wire \u0.w[1][20] ;
 wire \u0.w[1][21] ;
 wire \u0.w[1][22] ;
 wire \u0.w[1][23] ;
 wire \u0.w[1][24] ;
 wire \u0.w[1][25] ;
 wire \u0.w[1][26] ;
 wire \u0.w[1][27] ;
 wire \u0.w[1][28] ;
 wire \u0.w[1][29] ;
 wire \u0.w[1][2] ;
 wire \u0.w[1][30] ;
 wire \u0.w[1][31] ;
 wire \u0.w[1][3] ;
 wire \u0.w[1][4] ;
 wire \u0.w[1][5] ;
 wire \u0.w[1][6] ;
 wire \u0.w[1][7] ;
 wire \u0.w[1][8] ;
 wire \u0.w[1][9] ;
 wire \u0.w[2][0] ;
 wire \u0.w[2][10] ;
 wire \u0.w[2][11] ;
 wire \u0.w[2][12] ;
 wire \u0.w[2][13] ;
 wire \u0.w[2][14] ;
 wire \u0.w[2][15] ;
 wire \u0.w[2][16] ;
 wire \u0.w[2][17] ;
 wire \u0.w[2][18] ;
 wire \u0.w[2][19] ;
 wire \u0.w[2][1] ;
 wire \u0.w[2][20] ;
 wire \u0.w[2][21] ;
 wire \u0.w[2][22] ;
 wire \u0.w[2][23] ;
 wire \u0.w[2][24] ;
 wire \u0.w[2][25] ;
 wire \u0.w[2][26] ;
 wire \u0.w[2][27] ;
 wire \u0.w[2][28] ;
 wire \u0.w[2][29] ;
 wire \u0.w[2][2] ;
 wire \u0.w[2][30] ;
 wire \u0.w[2][31] ;
 wire \u0.w[2][3] ;
 wire \u0.w[2][4] ;
 wire \u0.w[2][5] ;
 wire \u0.w[2][6] ;
 wire \u0.w[2][7] ;
 wire \u0.w[2][8] ;
 wire \u0.w[2][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net928;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net647;
 wire net64;
 wire net66;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net45;
 wire net55;
 wire net56;
 wire net65;
 wire net67;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net787;
 wire net788;
 wire net789;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net943;
 wire net944;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net63;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net556;
 wire net557;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net832;
 wire net833;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net885;
 wire net886;
 wire net892;
 wire net895;
 wire net896;
 wire net918;
 wire net919;
 wire net920;
 wire net926;
 wire net927;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net940;
 wire net941;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net979;
 wire net980;
 wire net993;
 wire net1011;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1146;
 wire net1147;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1273;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16211_ (.A1(\u0.w[0][19] ),
    .A2(\u0.w[2][19] ),
    .ZN(_07232_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16212_ (.A1(\u0.w[1][19] ),
    .A2(\u0.subword[19] ),
    .Z(_07243_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16213_ (.A1(\u0.tmp_w[19] ),
    .A2(_07243_),
    .Z(_07254_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16214_ (.A1(_07232_),
    .A2(_07254_),
    .Z(_07265_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16215_ (.I(net216),
    .ZN(_07276_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16216_ (.I(_07276_),
    .Z(_07286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16217_ (.A1(_07265_),
    .A2(_07286_),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16218_ (.A1(_07276_),
    .A2(net126),
    .Z(_07308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16219_ (.A1(_07297_),
    .A2(_07308_),
    .ZN(_07319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16220_ (.I(_07319_),
    .ZN(_07330_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16221_ (.I(_07330_),
    .Z(_07341_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16222_ (.I(_07341_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16223_ (.A1(\u0.w[0][16] ),
    .A2(\u0.w[2][16] ),
    .ZN(_07361_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16224_ (.A1(\u0.subword[16] ),
    .A2(\u0.w[1][16] ),
    .Z(_07372_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16225_ (.A1(\u0.tmp_w[16] ),
    .A2(_07372_),
    .Z(_07383_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16226_ (.A1(_07361_),
    .A2(_07383_),
    .Z(_07394_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16227_ (.I(_07286_),
    .Z(_07404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16228_ (.A1(_07394_),
    .A2(_07404_),
    .ZN(_07415_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16229_ (.I(net123),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16230_ (.I(net216),
    .Z(_07437_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16231_ (.A1(_07426_),
    .A2(_07437_),
    .Z(_07448_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16232_ (.I(_07448_),
    .ZN(_07458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16233_ (.A1(_07458_),
    .A2(_07415_),
    .ZN(_15543_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16234_ (.A1(\u0.w[0][17] ),
    .A2(\u0.w[2][17] ),
    .ZN(_07463_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16235_ (.A1(\u0.w[1][17] ),
    .A2(\u0.subword[17] ),
    .Z(_07464_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16236_ (.A1(\u0.tmp_w[17] ),
    .A2(_07464_),
    .Z(_07465_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16237_ (.A1(_07465_),
    .A2(_07463_),
    .Z(_07466_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _16238_ (.I(_07276_),
    .Z(_07467_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _16239_ (.I(_07467_),
    .Z(_07468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16240_ (.A1(_07468_),
    .A2(_07466_),
    .ZN(_07469_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16241_ (.I(net124),
    .ZN(_07470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16242_ (.A1(_07470_),
    .A2(_07437_),
    .Z(_07471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16243_ (.I(_07471_),
    .ZN(_07472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16244_ (.A1(_07472_),
    .A2(_07469_),
    .ZN(_15548_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16245_ (.A1(\u0.w[0][21] ),
    .A2(\u0.w[2][21] ),
    .ZN(_07473_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16246_ (.A1(\u0.w[1][21] ),
    .A2(\u0.subword[21] ),
    .Z(_07475_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16247_ (.A1(\u0.tmp_w[21] ),
    .A2(_07475_),
    .Z(_07477_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16248_ (.A1(_07473_),
    .A2(_07477_),
    .Z(_07479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16249_ (.A1(_07479_),
    .A2(_07404_),
    .Z(_07481_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16250_ (.A1(_07468_),
    .A2(net129),
    .ZN(_07482_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16251_ (.A1(_07481_),
    .A2(_07482_),
    .ZN(_07484_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16252_ (.I(_07484_),
    .Z(_07486_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16253_ (.I(_07486_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16254_ (.A1(\u0.w[0][20] ),
    .A2(\u0.w[2][20] ),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16255_ (.A1(\u0.w[1][20] ),
    .A2(\u0.subword[20] ),
    .Z(_07491_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16256_ (.A1(\u0.tmp_w[20] ),
    .A2(_07491_),
    .Z(_07493_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16257_ (.A1(_07489_),
    .A2(_07493_),
    .Z(_07495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16258_ (.A1(_07495_),
    .A2(_07286_),
    .Z(_07497_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16259_ (.I(net128),
    .ZN(_07498_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16260_ (.A1(_07498_),
    .A2(_07437_),
    .Z(_07504_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16261_ (.A1(_07497_),
    .A2(_07504_),
    .ZN(_07513_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16262_ (.I(_07513_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16263_ (.A1(\u0.w[0][18] ),
    .A2(\u0.w[2][18] ),
    .Z(_07526_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16264_ (.A1(\u0.subword[18] ),
    .A2(\u0.w[1][18] ),
    .Z(_07531_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16265_ (.A1(\u0.tmp_w[18] ),
    .A2(_07531_),
    .Z(_07532_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16266_ (.A1(_07526_),
    .A2(_07532_),
    .Z(_07533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16267_ (.A1(_07533_),
    .A2(_07276_),
    .ZN(_07534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16268_ (.A1(net216),
    .A2(net125),
    .ZN(_07535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16269_ (.A1(_07534_),
    .A2(_07535_),
    .ZN(_07536_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16270_ (.I(_07536_),
    .Z(_07537_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16271_ (.I(_07537_),
    .Z(_15562_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16272_ (.A1(\u0.w[0][0] ),
    .A2(\u0.w[2][0] ),
    .ZN(_07538_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16273_ (.A1(\u0.subword[0] ),
    .A2(\u0.w[1][0] ),
    .Z(_07539_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16274_ (.A1(\u0.tmp_w[0] ),
    .A2(_07539_),
    .Z(_07540_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _16275_ (.A1(_07540_),
    .A2(_07538_),
    .Z(_07541_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _16276_ (.I(_07467_),
    .Z(_07542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16277_ (.A1(_07541_),
    .A2(_07542_),
    .ZN(_07543_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16278_ (.I(net45),
    .ZN(_07544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16279_ (.A1(_07544_),
    .A2(_07437_),
    .Z(_07545_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16280_ (.I(_07545_),
    .ZN(_07546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16281_ (.A1(_07546_),
    .A2(_07543_),
    .ZN(_15611_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16282_ (.A1(\u0.w[0][1] ),
    .A2(\u0.w[2][1] ),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16283_ (.A1(\u0.subword[1] ),
    .A2(\u0.w[1][1] ),
    .Z(_07548_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16284_ (.A1(\u0.tmp_w[1] ),
    .A2(_07548_),
    .Z(_07549_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16285_ (.A1(_07549_),
    .A2(_07547_),
    .Z(_07550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16286_ (.A1(_07550_),
    .A2(_07404_),
    .ZN(_07551_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16287_ (.I(net127),
    .ZN(_07552_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16288_ (.A1(_07552_),
    .A2(_07437_),
    .Z(_07553_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16289_ (.I(_07553_),
    .ZN(_07554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16290_ (.A1(_07554_),
    .A2(_07551_),
    .ZN(_15616_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16291_ (.A1(\u0.w[0][2] ),
    .A2(\u0.w[2][2] ),
    .ZN(_07555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16292_ (.I(\u0.tmp_w[2] ),
    .ZN(_07556_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16293_ (.A1(\u0.subword[2] ),
    .A2(\u0.w[1][2] ),
    .Z(_07557_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16294_ (.A1(_07556_),
    .A2(_07557_),
    .Z(_07558_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _16295_ (.A1(_07555_),
    .A2(_07558_),
    .Z(_07559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16296_ (.A1(_07559_),
    .A2(_07467_),
    .ZN(_07560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16297_ (.A1(net216),
    .A2(net138),
    .Z(_07561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16298_ (.I(_07561_),
    .ZN(_07562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16299_ (.A1(_07560_),
    .A2(_07562_),
    .ZN(_07563_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16300_ (.I(_07563_),
    .Z(_15630_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16301_ (.A1(\u0.w[0][3] ),
    .A2(\u0.w[2][3] ),
    .ZN(_07564_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16302_ (.A1(\u0.w[1][3] ),
    .A2(\u0.subword[3] ),
    .Z(_07565_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16303_ (.A1(\u0.tmp_w[3] ),
    .A2(_07565_),
    .Z(_07566_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16304_ (.A1(_07564_),
    .A2(_07566_),
    .Z(_07567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16305_ (.A1(_07567_),
    .A2(_07467_),
    .ZN(_07568_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16306_ (.A1(_07286_),
    .A2(net149),
    .Z(_07569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16307_ (.A1(_07568_),
    .A2(_07569_),
    .ZN(_07570_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16308_ (.I(_07570_),
    .ZN(_07571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16309_ (.I(_07571_),
    .Z(_07572_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16310_ (.I(_07572_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16311_ (.A1(\u0.w[0][4] ),
    .A2(\u0.w[2][4] ),
    .ZN(_07573_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16312_ (.A1(\u0.w[1][4] ),
    .A2(\u0.subword[4] ),
    .Z(_07574_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16313_ (.A1(\u0.tmp_w[4] ),
    .A2(_07574_),
    .Z(_07575_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16314_ (.A1(_07573_),
    .A2(_07575_),
    .Z(_07576_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16315_ (.A1(_07286_),
    .A2(net160),
    .ZN(_07577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16316_ (.A1(_07576_),
    .A2(_07467_),
    .B(_07577_),
    .ZN(_07578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16317_ (.I(_07578_),
    .Z(_07579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16318_ (.I(_07579_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16319_ (.A1(\u0.w[0][5] ),
    .A2(\u0.w[2][5] ),
    .ZN(_07580_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16320_ (.A1(\u0.w[1][5] ),
    .A2(\u0.subword[5] ),
    .Z(_07581_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16321_ (.A1(\u0.tmp_w[5] ),
    .A2(_07581_),
    .Z(_07582_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16322_ (.A1(_07580_),
    .A2(_07582_),
    .Z(_07583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16323_ (.A1(_07583_),
    .A2(_07404_),
    .Z(_07584_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16324_ (.A1(_07468_),
    .A2(net171),
    .ZN(_07585_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16325_ (.A1(_07584_),
    .A2(_07585_),
    .ZN(_07586_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16326_ (.I(_07586_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16327_ (.A1(\u0.w[1][6] ),
    .A2(\u0.subword[6] ),
    .Z(_07587_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16328_ (.A1(\u0.w[0][6] ),
    .A2(\u0.w[2][6] ),
    .ZN(_07588_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16329_ (.A1(\u0.tmp_w[6] ),
    .A2(_07587_),
    .A3(_07588_),
    .Z(_07589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16330_ (.A1(_07589_),
    .A2(_07542_),
    .Z(_07590_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16331_ (.A1(_07542_),
    .A2(net182),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16332_ (.A1(_07590_),
    .A2(_07591_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16333_ (.A1(\u0.w[1][7] ),
    .A2(\u0.subword[7] ),
    .Z(_07592_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16334_ (.A1(\u0.w[0][7] ),
    .A2(\u0.w[2][7] ),
    .ZN(_07593_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16335_ (.A1(\u0.tmp_w[7] ),
    .A2(_07592_),
    .A3(_07593_),
    .Z(_07594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16336_ (.A1(_07594_),
    .A2(_07542_),
    .Z(_07595_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16337_ (.I(_07468_),
    .Z(_07596_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16338_ (.A1(_07596_),
    .A2(net193),
    .ZN(_07597_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16339_ (.A1(_07595_),
    .A2(_07597_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16340_ (.A1(\u0.w[0][8] ),
    .A2(\u0.w[2][8] ),
    .ZN(_07598_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16341_ (.A1(\u0.subword[8] ),
    .A2(\u0.w[1][8] ),
    .Z(_07599_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16342_ (.A1(\u0.tmp_w[8] ),
    .A2(_07599_),
    .Z(_07600_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _16343_ (.A1(_07600_),
    .A2(_07598_),
    .Z(_07601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16344_ (.A1(_07601_),
    .A2(_07468_),
    .ZN(_07602_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16345_ (.I(net204),
    .ZN(_07603_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16346_ (.A1(_07603_),
    .A2(net216),
    .Z(_07604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16347_ (.I(_07604_),
    .ZN(_07605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16348_ (.A1(_07605_),
    .A2(_07602_),
    .ZN(_15577_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16349_ (.A1(\u0.w[0][9] ),
    .A2(\u0.w[2][9] ),
    .ZN(_07606_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16350_ (.A1(\u0.subword[9] ),
    .A2(\u0.w[1][9] ),
    .Z(_07607_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16351_ (.A1(\u0.tmp_w[9] ),
    .A2(_07607_),
    .Z(_07608_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _16352_ (.A1(_07608_),
    .A2(_07606_),
    .Z(_07609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16353_ (.A1(_07404_),
    .A2(_07609_),
    .ZN(_07610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16354_ (.I(net215),
    .ZN(_07611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16355_ (.A1(_07611_),
    .A2(_07437_),
    .Z(_07612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16356_ (.I(_07612_),
    .ZN(_07613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16357_ (.A1(_07613_),
    .A2(_07610_),
    .ZN(_15582_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16358_ (.A1(\u0.w[0][10] ),
    .A2(\u0.w[2][10] ),
    .ZN(_07614_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _16359_ (.I(\u0.tmp_w[10] ),
    .ZN(_07615_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16360_ (.A1(\u0.w[1][10] ),
    .A2(\u0.subword[10] ),
    .Z(_07616_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16361_ (.A1(_07615_),
    .A2(_07616_),
    .Z(_07617_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _16362_ (.A1(_07617_),
    .A2(_07614_),
    .Z(_07618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16363_ (.A1(_07618_),
    .A2(_07286_),
    .ZN(_07619_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16364_ (.A1(net216),
    .A2(net99),
    .Z(_07620_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16365_ (.I(_07620_),
    .ZN(_07621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16366_ (.A1(_07621_),
    .A2(_07619_),
    .ZN(_07622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16367_ (.I(_07622_),
    .Z(_15596_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16368_ (.A1(\u0.w[0][11] ),
    .A2(\u0.w[2][11] ),
    .ZN(_07623_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16369_ (.A1(\u0.w[1][11] ),
    .A2(\u0.subword[11] ),
    .Z(_07624_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16370_ (.A1(\u0.tmp_w[11] ),
    .A2(_07624_),
    .Z(_07625_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16371_ (.A1(_07623_),
    .A2(_07625_),
    .Z(_07626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16372_ (.A1(_07626_),
    .A2(_07286_),
    .ZN(_07627_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16373_ (.A1(_07276_),
    .A2(net110),
    .Z(_07628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16374_ (.A1(_07627_),
    .A2(_07628_),
    .ZN(_07629_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16375_ (.I(_07629_),
    .ZN(_07630_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16376_ (.I(_07630_),
    .Z(_07631_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16377_ (.I(_07631_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16378_ (.A1(\u0.w[0][12] ),
    .A2(\u0.w[2][12] ),
    .ZN(_07632_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16379_ (.A1(\u0.w[1][12] ),
    .A2(\u0.subword[12] ),
    .Z(_07633_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16380_ (.A1(\u0.tmp_w[12] ),
    .A2(_07633_),
    .Z(_07634_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16381_ (.A1(_07632_),
    .A2(_07634_),
    .Z(_07635_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16382_ (.I(net119),
    .ZN(_07636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16383_ (.I0(_07635_),
    .I1(_07636_),
    .S(net216),
    .Z(_07637_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16384_ (.I(_07637_),
    .Z(_07638_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16385_ (.I(_07638_),
    .ZN(_07639_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16386_ (.I(_07639_),
    .Z(_07640_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16387_ (.I(_07640_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16388_ (.A1(\u0.w[0][13] ),
    .A2(\u0.w[2][13] ),
    .ZN(_07641_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16389_ (.A1(\u0.w[1][13] ),
    .A2(\u0.subword[13] ),
    .Z(_07642_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16390_ (.A1(\u0.tmp_w[13] ),
    .A2(_07642_),
    .Z(_07643_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16391_ (.A1(_07641_),
    .A2(_07643_),
    .Z(_07644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16392_ (.A1(_07644_),
    .A2(_07404_),
    .Z(_07645_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16393_ (.A1(_07468_),
    .A2(net120),
    .ZN(_07646_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16394_ (.A1(_07645_),
    .A2(_07646_),
    .ZN(_07647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16395_ (.I(_07647_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16396_ (.A1(\u0.w[0][14] ),
    .A2(\u0.w[2][14] ),
    .ZN(_07648_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16397_ (.A1(\u0.w[1][14] ),
    .A2(\u0.subword[14] ),
    .Z(_07649_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16398_ (.A1(\u0.tmp_w[14] ),
    .A2(_07649_),
    .Z(_07650_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16399_ (.A1(_07648_),
    .A2(_07650_),
    .Z(_07651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16400_ (.A1(_07651_),
    .A2(_07542_),
    .Z(_07652_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16401_ (.A1(_07596_),
    .A2(net121),
    .ZN(_07653_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16402_ (.A1(_07652_),
    .A2(_07653_),
    .ZN(_07654_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16403_ (.I(_07654_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16404_ (.A1(\u0.w[1][15] ),
    .A2(\u0.subword[15] ),
    .Z(_07655_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16405_ (.A1(\u0.w[0][15] ),
    .A2(\u0.w[2][15] ),
    .ZN(_07656_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16406_ (.A1(\u0.tmp_w[15] ),
    .A2(_07655_),
    .A3(_07656_),
    .Z(_07657_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16407_ (.A1(_07657_),
    .A2(_07596_),
    .Z(_07658_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16408_ (.A1(_07596_),
    .A2(net122),
    .ZN(_07659_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16409_ (.A1(_07658_),
    .A2(_07659_),
    .ZN(_07660_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16410_ (.I(_07660_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16411_ (.A1(\u0.w[1][22] ),
    .A2(\u0.subword[22] ),
    .Z(_07661_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16412_ (.A1(\u0.w[0][22] ),
    .A2(\u0.w[2][22] ),
    .ZN(_07662_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16413_ (.A1(\u0.tmp_w[22] ),
    .A2(_07661_),
    .A3(_07662_),
    .Z(_07663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16414_ (.A1(_07663_),
    .A2(_07542_),
    .Z(_07664_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16415_ (.A1(_07542_),
    .A2(net130),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16416_ (.A1(_07664_),
    .A2(_07665_),
    .ZN(_07666_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16417_ (.I(_07666_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16418_ (.A1(\u0.w[1][23] ),
    .A2(\u0.subword[23] ),
    .Z(_07667_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16419_ (.A1(\u0.w[0][23] ),
    .A2(\u0.w[2][23] ),
    .ZN(_07668_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16420_ (.A1(\u0.tmp_w[23] ),
    .A2(_07667_),
    .A3(_07668_),
    .Z(_07669_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16421_ (.A1(_07669_),
    .A2(_07596_),
    .Z(_07670_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16422_ (.A1(_07596_),
    .A2(net131),
    .ZN(_07671_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16423_ (.A1(_07670_),
    .A2(_07671_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _16424_ (.I(\u0.w[0][24] ),
    .ZN(_07672_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16425_ (.A1(\u0.r0.out[24] ),
    .A2(\u0.w[2][24] ),
    .Z(_07673_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16426_ (.A1(_07672_),
    .A2(_07673_),
    .Z(_07674_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16427_ (.A1(\u0.w[1][24] ),
    .A2(\u0.subword[24] ),
    .Z(_07675_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16428_ (.A1(_07675_),
    .A2(\u0.tmp_w[24] ),
    .Z(_07676_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16429_ (.A1(_07676_),
    .A2(_07674_),
    .Z(_07677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16430_ (.A1(_07674_),
    .A2(_07676_),
    .ZN(_07678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16431_ (.A1(_07677_),
    .A2(_07678_),
    .ZN(_07679_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16432_ (.A1(_07437_),
    .A2(net132),
    .Z(_07680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16433_ (.A1(net764),
    .A2(_07542_),
    .B(_07680_),
    .ZN(_15645_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16434_ (.A1(\u0.w[2][25] ),
    .A2(\u0.w[0][25] ),
    .Z(_07681_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16435_ (.A1(\u0.r0.out[25] ),
    .A2(_07681_),
    .Z(_07682_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16436_ (.A1(\u0.tmp_w[25] ),
    .A2(\u0.w[1][25] ),
    .Z(_07683_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16437_ (.A1(\u0.subword[25] ),
    .A2(_07683_),
    .Z(_07684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16438_ (.A1(_07682_),
    .A2(_07684_),
    .Z(_07685_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16439_ (.A1(_07682_),
    .A2(_07684_),
    .ZN(_07686_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _16440_ (.A1(_07685_),
    .A2(_07686_),
    .B(_07467_),
    .ZN(_07687_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16441_ (.A1(_07467_),
    .A2(net133),
    .Z(_07688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16442_ (.A1(_07687_),
    .A2(_07688_),
    .ZN(_15650_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16443_ (.I(\u0.w[0][26] ),
    .ZN(_07689_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16444_ (.A1(\u0.w[2][26] ),
    .A2(\u0.r0.out[26] ),
    .Z(_07690_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16445_ (.A1(_07689_),
    .A2(_07690_),
    .Z(_07691_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16446_ (.A1(\u0.w[1][26] ),
    .A2(\u0.subword[26] ),
    .Z(_07692_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16447_ (.A1(\u0.tmp_w[26] ),
    .A2(_07692_),
    .Z(_07693_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16448_ (.A1(_07693_),
    .A2(_07691_),
    .Z(_07694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16449_ (.A1(_07694_),
    .A2(_07286_),
    .ZN(_07695_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16450_ (.A1(_07286_),
    .A2(net134),
    .Z(_07696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16451_ (.A1(_07696_),
    .A2(_07695_),
    .ZN(_07697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16452_ (.I(_07697_),
    .Z(_15664_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16453_ (.A1(\u0.w[0][27] ),
    .A2(\u0.w[2][27] ),
    .Z(_07698_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16454_ (.A1(\u0.r0.out[27] ),
    .A2(_07698_),
    .Z(_07699_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16455_ (.A1(\u0.tmp_w[27] ),
    .A2(\u0.w[1][27] ),
    .Z(_07700_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16456_ (.A1(\u0.subword[27] ),
    .A2(_07700_),
    .Z(_07701_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16457_ (.A1(_07699_),
    .A2(_07701_),
    .Z(_07702_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16458_ (.A1(_07699_),
    .A2(_07701_),
    .ZN(_07703_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16459_ (.A1(_07702_),
    .A2(net216),
    .A3(_07703_),
    .Z(_07704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16460_ (.A1(net216),
    .A2(net135),
    .ZN(_07705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16461_ (.A1(_07705_),
    .A2(_07704_),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16462_ (.I(net825),
    .Z(_07707_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16463_ (.I(_07707_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16464_ (.A1(\u0.w[0][28] ),
    .A2(\u0.w[2][28] ),
    .Z(_07708_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16465_ (.A1(\u0.r0.out[28] ),
    .A2(_07708_),
    .Z(_07709_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16466_ (.A1(\u0.tmp_w[28] ),
    .A2(\u0.w[1][28] ),
    .Z(_07710_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16467_ (.A1(\u0.subword[28] ),
    .A2(_07710_),
    .Z(_07711_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16468_ (.A1(_07709_),
    .A2(_07711_),
    .Z(_07712_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16469_ (.A1(_07709_),
    .A2(_07711_),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16470_ (.A1(_07712_),
    .A2(_07713_),
    .B(_07404_),
    .ZN(_07714_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16471_ (.A1(_07467_),
    .A2(net136),
    .Z(_07715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16472_ (.A1(_07714_),
    .A2(_07715_),
    .ZN(_07716_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16473_ (.I(_07716_),
    .ZN(_07717_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16474_ (.I(_07717_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16475_ (.A1(\u0.w[0][29] ),
    .A2(\u0.w[2][29] ),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16476_ (.A1(\u0.r0.out[29] ),
    .A2(_07718_),
    .Z(_07719_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16477_ (.A1(\u0.tmp_w[29] ),
    .A2(\u0.w[1][29] ),
    .Z(_07720_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16478_ (.A1(\u0.subword[29] ),
    .A2(_07720_),
    .Z(_07721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16479_ (.A1(_07719_),
    .A2(_07721_),
    .Z(_07722_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16480_ (.A1(_07719_),
    .A2(_07721_),
    .ZN(_07723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16481_ (.A1(_07722_),
    .A2(_07723_),
    .B(_07468_),
    .ZN(_07724_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16482_ (.A1(_07404_),
    .A2(net137),
    .Z(_07725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16483_ (.A1(_07724_),
    .A2(_07725_),
    .ZN(_07726_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16484_ (.I(_07726_),
    .ZN(_07727_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16485_ (.I(_07727_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16486_ (.A1(\u0.w[0][30] ),
    .A2(\u0.w[2][30] ),
    .A3(\u0.r0.out[30] ),
    .Z(_07728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16487_ (.I(\u0.w[1][30] ),
    .ZN(_07729_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16488_ (.A1(\u0.tmp_w[30] ),
    .A2(\u0.subword[30] ),
    .A3(_07729_),
    .Z(_07730_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16489_ (.A1(_07728_),
    .A2(_07730_),
    .Z(_07731_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16490_ (.I(net139),
    .ZN(_07732_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16491_ (.I(_07437_),
    .Z(_07733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16492_ (.A1(_07732_),
    .A2(_07733_),
    .Z(_07734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16493_ (.A1(_07731_),
    .A2(_07542_),
    .B(_07734_),
    .ZN(_07735_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16494_ (.I(_07735_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16495_ (.A1(\u0.w[0][31] ),
    .A2(\u0.w[2][31] ),
    .Z(_07736_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16496_ (.A1(\u0.r0.out[31] ),
    .A2(_07736_),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16497_ (.A1(\u0.w[1][31] ),
    .A2(\u0.subword[31] ),
    .A3(_07737_),
    .Z(_07738_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _16498_ (.I(\u0.tmp_w[31] ),
    .ZN(_07739_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16499_ (.A1(_07738_),
    .A2(_07739_),
    .Z(_07740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16500_ (.A1(_07738_),
    .A2(_07739_),
    .ZN(_07741_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16501_ (.A1(_07740_),
    .A2(_07596_),
    .A3(_07741_),
    .Z(_07742_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16502_ (.A1(_07596_),
    .A2(net140),
    .ZN(_07743_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16503_ (.A1(_07742_),
    .A2(_07743_),
    .Z(_07744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16504_ (.I(_07744_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16505_ (.A1(_07539_),
    .A2(_07538_),
    .ZN(_07745_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16506_ (.I(_07733_),
    .Z(_07746_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16507_ (.I(_07746_),
    .Z(_07747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16508_ (.I0(_07745_),
    .I1(net141),
    .S(_07747_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16509_ (.A1(_07548_),
    .A2(_07547_),
    .ZN(_07748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16510_ (.I0(_07748_),
    .I1(net142),
    .S(_07747_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16511_ (.A1(_07557_),
    .A2(_07555_),
    .ZN(_07749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16512_ (.I0(_07749_),
    .I1(net143),
    .S(_07747_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16513_ (.A1(_07565_),
    .A2(_07564_),
    .ZN(_07750_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16514_ (.I(_07746_),
    .Z(_07751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16515_ (.I0(_07750_),
    .I1(net144),
    .S(_07751_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16516_ (.A1(_07574_),
    .A2(_07573_),
    .ZN(_07752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16517_ (.I0(_07752_),
    .I1(net145),
    .S(_07751_),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16518_ (.A1(_07581_),
    .A2(_07580_),
    .ZN(_07753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16519_ (.I0(_07753_),
    .I1(net146),
    .S(_07751_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16520_ (.A1(_07587_),
    .A2(_07588_),
    .ZN(_07754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16521_ (.I0(_07754_),
    .I1(net147),
    .S(_07751_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16522_ (.A1(_07592_),
    .A2(_07593_),
    .ZN(_07755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16523_ (.I0(_07755_),
    .I1(net148),
    .S(_07751_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16524_ (.A1(_07599_),
    .A2(_07598_),
    .ZN(_07756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16525_ (.I0(_07756_),
    .I1(net150),
    .S(_07751_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16526_ (.A1(_07607_),
    .A2(_07606_),
    .ZN(_07757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16527_ (.I0(_07757_),
    .I1(net151),
    .S(_07751_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16528_ (.A1(_07616_),
    .A2(_07614_),
    .ZN(_07758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16529_ (.I0(_07758_),
    .I1(net152),
    .S(_07751_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16530_ (.A1(_07624_),
    .A2(_07623_),
    .ZN(_07759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16531_ (.I0(_07759_),
    .I1(net153),
    .S(_07751_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16532_ (.A1(_07633_),
    .A2(_07632_),
    .ZN(_07760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16533_ (.I0(_07760_),
    .I1(net154),
    .S(_07751_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16534_ (.A1(_07642_),
    .A2(_07641_),
    .ZN(_07761_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16535_ (.I(_07746_),
    .Z(_07762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16536_ (.I0(_07761_),
    .I1(net155),
    .S(_07762_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16537_ (.A1(_07649_),
    .A2(_07648_),
    .ZN(_07763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16538_ (.I0(_07763_),
    .I1(net156),
    .S(_07762_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16539_ (.A1(_07655_),
    .A2(_07656_),
    .ZN(_07764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16540_ (.I0(_07764_),
    .I1(net157),
    .S(_07762_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16541_ (.A1(_07372_),
    .A2(_07361_),
    .ZN(_07765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16542_ (.I0(_07765_),
    .I1(net158),
    .S(_07762_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16543_ (.A1(_07464_),
    .A2(_07463_),
    .ZN(_07766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16544_ (.I0(_07766_),
    .I1(net159),
    .S(_07762_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16545_ (.A1(_07526_),
    .A2(_07531_),
    .Z(_07767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16546_ (.I0(_07767_),
    .I1(net161),
    .S(_07762_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16547_ (.A1(_07243_),
    .A2(_07232_),
    .ZN(_07768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16548_ (.I0(_07768_),
    .I1(net162),
    .S(_07762_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16549_ (.A1(_07491_),
    .A2(_07489_),
    .ZN(_07769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16550_ (.I0(_07769_),
    .I1(net163),
    .S(_07762_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16551_ (.A1(_07475_),
    .A2(_07473_),
    .ZN(_07770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16552_ (.I0(_07770_),
    .I1(net164),
    .S(_07762_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16553_ (.A1(_07661_),
    .A2(_07662_),
    .ZN(_07771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16554_ (.I0(_07771_),
    .I1(net165),
    .S(_07762_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16555_ (.A1(_07667_),
    .A2(_07668_),
    .ZN(_07772_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _16556_ (.I(_07733_),
    .Z(_07773_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16557_ (.I(_07773_),
    .Z(_07774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16558_ (.I0(_07772_),
    .I1(net166),
    .S(_07774_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16559_ (.A1(_07675_),
    .A2(net708),
    .ZN(_07775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16560_ (.I0(_07775_),
    .I1(net167),
    .S(_07774_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16561_ (.A1(\u0.w[1][25] ),
    .A2(\u0.subword[25] ),
    .A3(net710),
    .Z(_07776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16562_ (.I0(_07776_),
    .I1(net168),
    .S(_07774_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16563_ (.A1(_07692_),
    .A2(_07691_),
    .ZN(_07777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16564_ (.I0(_07777_),
    .I1(net169),
    .S(_07774_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16565_ (.A1(\u0.w[1][27] ),
    .A2(\u0.subword[27] ),
    .A3(_07699_),
    .Z(_07778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16566_ (.I0(_07778_),
    .I1(net170),
    .S(_07774_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16567_ (.A1(\u0.w[1][28] ),
    .A2(\u0.subword[28] ),
    .A3(_07709_),
    .Z(_07779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16568_ (.I0(_07779_),
    .I1(net172),
    .S(_07774_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16569_ (.A1(\u0.w[1][29] ),
    .A2(\u0.subword[29] ),
    .A3(_07719_),
    .Z(_07780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16570_ (.I0(_07780_),
    .I1(net173),
    .S(_07774_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16571_ (.A1(\u0.w[1][30] ),
    .A2(\u0.subword[30] ),
    .A3(_07728_),
    .Z(_07781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16572_ (.I0(_07781_),
    .I1(net174),
    .S(_07774_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16573_ (.I0(_07738_),
    .I1(net175),
    .S(_07774_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16574_ (.I(\u0.w[1][0] ),
    .ZN(_07782_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _16575_ (.I(_07733_),
    .Z(_07783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16576_ (.I0(\u0.w[1][0] ),
    .I1(net176),
    .S(_07783_),
    .Z(_07784_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16577_ (.A1(\u0.w[0][0] ),
    .A2(\u0.subword[0] ),
    .Z(_07785_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16578_ (.I(_07733_),
    .Z(_07786_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16579_ (.A1(\u0.w[0][0] ),
    .A2(\u0.subword[0] ),
    .ZN(_07787_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16580_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_07787_),
    .Z(_07788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16581_ (.I0(_07782_),
    .I1(_07784_),
    .S(_07788_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _16582_ (.I(_07733_),
    .Z(_07789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16583_ (.I0(\u0.w[1][1] ),
    .I1(net177),
    .S(_07789_),
    .Z(_07790_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16584_ (.I(\u0.w[1][1] ),
    .ZN(_07791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16585_ (.A1(\u0.w[0][1] ),
    .A2(\u0.subword[1] ),
    .Z(_07792_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16586_ (.I(_07596_),
    .Z(_07793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16587_ (.A1(\u0.w[0][1] ),
    .A2(\u0.subword[1] ),
    .ZN(_07794_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16588_ (.A1(_07792_),
    .A2(_07793_),
    .A3(_07794_),
    .Z(_07795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16589_ (.I0(_07790_),
    .I1(_07791_),
    .S(_07795_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16590_ (.I(\u0.w[1][2] ),
    .ZN(_07796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16591_ (.I0(\u0.w[1][2] ),
    .I1(net178),
    .S(_07783_),
    .Z(_07797_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16592_ (.A1(\u0.subword[2] ),
    .A2(\u0.w[0][2] ),
    .Z(_07798_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16593_ (.A1(\u0.subword[2] ),
    .A2(\u0.w[0][2] ),
    .ZN(_07799_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16594_ (.A1(_07798_),
    .A2(_07786_),
    .A3(_07799_),
    .Z(_07800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16595_ (.I0(_07796_),
    .I1(_07797_),
    .S(_07800_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16596_ (.I(\u0.w[1][3] ),
    .ZN(_07801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16597_ (.I0(\u0.w[1][3] ),
    .I1(net179),
    .S(_07783_),
    .Z(_07802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16598_ (.A1(\u0.w[0][3] ),
    .A2(\u0.subword[3] ),
    .Z(_07803_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16599_ (.A1(\u0.w[0][3] ),
    .A2(\u0.subword[3] ),
    .ZN(_07804_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16600_ (.A1(_07803_),
    .A2(_07786_),
    .A3(_07804_),
    .Z(_07805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16601_ (.I0(_07801_),
    .I1(_07802_),
    .S(_07805_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16602_ (.I(_07733_),
    .Z(_07806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16603_ (.I0(\u0.w[1][4] ),
    .I1(net180),
    .S(_07806_),
    .Z(_07807_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16604_ (.I(\u0.w[1][4] ),
    .ZN(_07808_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16605_ (.A1(\u0.w[0][4] ),
    .A2(\u0.subword[4] ),
    .Z(_07809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16606_ (.A1(\u0.w[0][4] ),
    .A2(\u0.subword[4] ),
    .ZN(_07810_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16607_ (.A1(_07809_),
    .A2(_07793_),
    .A3(_07810_),
    .Z(_07811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16608_ (.I0(_07807_),
    .I1(_07808_),
    .S(_07811_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16609_ (.A1(\u0.w[0][5] ),
    .A2(\u0.subword[5] ),
    .Z(_07812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16610_ (.A1(\u0.w[0][5] ),
    .A2(\u0.subword[5] ),
    .ZN(_07813_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16611_ (.A1(_07812_),
    .A2(_07793_),
    .A3(_07813_),
    .Z(_07814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16612_ (.I0(\u0.w[1][5] ),
    .I1(net181),
    .S(_07789_),
    .Z(_07815_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16613_ (.A1(_07814_),
    .A2(_07815_),
    .ZN(_07816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16614_ (.A1(\u0.w[1][5] ),
    .A2(_07814_),
    .B(_07816_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16615_ (.A1(\u0.w[0][6] ),
    .A2(\u0.subword[6] ),
    .Z(_07817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16616_ (.A1(\u0.w[0][6] ),
    .A2(\u0.subword[6] ),
    .ZN(_07818_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16617_ (.A1(_07817_),
    .A2(_07793_),
    .A3(_07818_),
    .Z(_07819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16618_ (.I0(\u0.w[1][6] ),
    .I1(net183),
    .S(_07789_),
    .Z(_07820_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16619_ (.A1(_07819_),
    .A2(_07820_),
    .ZN(_07821_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16620_ (.A1(\u0.w[1][6] ),
    .A2(_07819_),
    .B(_07821_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16621_ (.A1(\u0.w[0][7] ),
    .A2(\u0.subword[7] ),
    .Z(_07822_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16622_ (.A1(\u0.w[0][7] ),
    .A2(\u0.subword[7] ),
    .ZN(_07823_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16623_ (.A1(_07822_),
    .A2(_07746_),
    .A3(_07823_),
    .Z(_07824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16624_ (.I0(\u0.w[1][7] ),
    .I1(net184),
    .S(_07789_),
    .Z(_07825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16625_ (.A1(_07824_),
    .A2(_07825_),
    .ZN(_07826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16626_ (.A1(\u0.w[1][7] ),
    .A2(_07824_),
    .B(_07826_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16627_ (.I0(\u0.w[1][8] ),
    .I1(net185),
    .S(_07806_),
    .Z(_07827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16628_ (.I(\u0.w[1][8] ),
    .ZN(_07828_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16629_ (.A1(\u0.w[0][8] ),
    .A2(\u0.subword[8] ),
    .Z(_07829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16630_ (.A1(\u0.w[0][8] ),
    .A2(\u0.subword[8] ),
    .ZN(_07830_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16631_ (.A1(_07829_),
    .A2(_07793_),
    .A3(_07830_),
    .Z(_07831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16632_ (.I0(_07827_),
    .I1(_07828_),
    .S(_07831_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16633_ (.I0(\u0.w[1][9] ),
    .I1(net186),
    .S(_07806_),
    .Z(_07832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16634_ (.I(\u0.w[1][9] ),
    .ZN(_07833_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16635_ (.A1(\u0.w[0][9] ),
    .A2(\u0.subword[9] ),
    .Z(_07834_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16636_ (.I(_07596_),
    .Z(_07835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16637_ (.A1(\u0.w[0][9] ),
    .A2(\u0.subword[9] ),
    .ZN(_07836_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16638_ (.A1(_07834_),
    .A2(_07835_),
    .A3(_07836_),
    .Z(_07837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16639_ (.I0(_07832_),
    .I1(_07833_),
    .S(_07837_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16640_ (.I0(\u0.w[1][10] ),
    .I1(net187),
    .S(_07806_),
    .Z(_07838_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16641_ (.I(\u0.w[1][10] ),
    .ZN(_07839_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16642_ (.A1(\u0.subword[10] ),
    .A2(\u0.w[0][10] ),
    .Z(_07840_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16643_ (.A1(\u0.subword[10] ),
    .A2(\u0.w[0][10] ),
    .ZN(_07841_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16644_ (.A1(_07840_),
    .A2(_07835_),
    .A3(_07841_),
    .Z(_07842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16645_ (.I0(_07838_),
    .I1(_07839_),
    .S(_07842_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16646_ (.I(\u0.w[1][11] ),
    .ZN(_07843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16647_ (.I0(\u0.w[1][11] ),
    .I1(net188),
    .S(_07783_),
    .Z(_07844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16648_ (.A1(\u0.w[0][11] ),
    .A2(\u0.subword[11] ),
    .Z(_07845_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16649_ (.A1(\u0.w[0][11] ),
    .A2(\u0.subword[11] ),
    .ZN(_07846_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16650_ (.A1(_07845_),
    .A2(_07786_),
    .A3(_07846_),
    .Z(_07847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16651_ (.I0(_07843_),
    .I1(_07844_),
    .S(_07847_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16652_ (.I0(\u0.w[1][12] ),
    .I1(net189),
    .S(_07806_),
    .Z(_07848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16653_ (.I(\u0.w[1][12] ),
    .ZN(_07849_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16654_ (.A1(\u0.w[0][12] ),
    .A2(\u0.subword[12] ),
    .Z(_07850_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16655_ (.A1(\u0.w[0][12] ),
    .A2(\u0.subword[12] ),
    .ZN(_07851_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16656_ (.A1(_07850_),
    .A2(_07835_),
    .A3(_07851_),
    .Z(_07852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16657_ (.I0(_07848_),
    .I1(_07849_),
    .S(_07852_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16658_ (.A1(\u0.w[0][13] ),
    .A2(\u0.subword[13] ),
    .Z(_07853_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16659_ (.A1(\u0.w[0][13] ),
    .A2(\u0.subword[13] ),
    .ZN(_07854_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16660_ (.A1(_07853_),
    .A2(_07746_),
    .A3(_07854_),
    .Z(_07855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16661_ (.I0(\u0.w[1][13] ),
    .I1(net190),
    .S(_07789_),
    .Z(_07856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16662_ (.A1(_07855_),
    .A2(_07856_),
    .ZN(_07857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16663_ (.A1(\u0.w[1][13] ),
    .A2(_07855_),
    .B(_07857_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16664_ (.A1(\u0.w[0][14] ),
    .A2(\u0.subword[14] ),
    .Z(_07858_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16665_ (.A1(\u0.w[0][14] ),
    .A2(\u0.subword[14] ),
    .ZN(_07859_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16666_ (.A1(_07858_),
    .A2(_07746_),
    .A3(_07859_),
    .Z(_07860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16667_ (.I0(\u0.w[1][14] ),
    .I1(net191),
    .S(_07789_),
    .Z(_07861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16668_ (.A1(_07860_),
    .A2(_07861_),
    .ZN(_07862_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16669_ (.A1(\u0.w[1][14] ),
    .A2(_07860_),
    .B(_07862_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16670_ (.A1(\u0.w[0][15] ),
    .A2(\u0.subword[15] ),
    .Z(_07863_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16671_ (.A1(\u0.w[0][15] ),
    .A2(\u0.subword[15] ),
    .ZN(_07864_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16672_ (.A1(_07863_),
    .A2(_07746_),
    .A3(_07864_),
    .Z(_07865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16673_ (.I0(\u0.w[1][15] ),
    .I1(net192),
    .S(_07789_),
    .Z(_07866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16674_ (.A1(_07865_),
    .A2(_07866_),
    .ZN(_07867_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16675_ (.A1(\u0.w[1][15] ),
    .A2(_07865_),
    .B(_07867_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16676_ (.I0(\u0.w[1][16] ),
    .I1(net194),
    .S(_07806_),
    .Z(_07868_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16677_ (.I(\u0.w[1][16] ),
    .ZN(_07869_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16678_ (.A1(\u0.w[0][16] ),
    .A2(\u0.subword[16] ),
    .Z(_07870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16679_ (.A1(\u0.w[0][16] ),
    .A2(\u0.subword[16] ),
    .ZN(_07871_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16680_ (.A1(_07870_),
    .A2(_07835_),
    .A3(_07871_),
    .Z(_07872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16681_ (.I0(_07868_),
    .I1(_07869_),
    .S(_07872_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16682_ (.I0(net1033),
    .I1(net195),
    .S(_07806_),
    .Z(_07873_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16683_ (.I(net1030),
    .ZN(_07874_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16684_ (.A1(\u0.w[0][17] ),
    .A2(net1035),
    .Z(_07875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16685_ (.A1(\u0.w[0][17] ),
    .A2(net1035),
    .ZN(_07876_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16686_ (.A1(_07875_),
    .A2(_07835_),
    .A3(_07876_),
    .Z(_07877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16687_ (.I0(_07873_),
    .I1(_07874_),
    .S(_07877_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16688_ (.I0(\u0.w[1][18] ),
    .I1(net196),
    .S(_07806_),
    .Z(_07878_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16689_ (.I(\u0.w[1][18] ),
    .ZN(_07879_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16690_ (.A1(\u0.subword[18] ),
    .A2(\u0.w[0][18] ),
    .Z(_07880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16691_ (.A1(\u0.subword[18] ),
    .A2(\u0.w[0][18] ),
    .ZN(_07881_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16692_ (.A1(_07880_),
    .A2(_07835_),
    .A3(_07881_),
    .Z(_07882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16693_ (.I0(_07878_),
    .I1(_07879_),
    .S(_07882_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16694_ (.I0(\u0.w[1][19] ),
    .I1(net197),
    .S(_07806_),
    .Z(_07883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16695_ (.I(\u0.w[1][19] ),
    .ZN(_07884_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16696_ (.A1(\u0.w[0][19] ),
    .A2(\u0.subword[19] ),
    .Z(_07885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16697_ (.A1(\u0.w[0][19] ),
    .A2(\u0.subword[19] ),
    .ZN(_07886_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16698_ (.A1(_07885_),
    .A2(_07835_),
    .A3(_07886_),
    .Z(_07887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16699_ (.I0(_07883_),
    .I1(_07884_),
    .S(_07887_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16700_ (.I(\u0.w[1][20] ),
    .ZN(_07888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16701_ (.I0(\u0.w[1][20] ),
    .I1(net198),
    .S(_07783_),
    .Z(_07889_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16702_ (.A1(\u0.w[0][20] ),
    .A2(\u0.subword[20] ),
    .Z(_07890_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16703_ (.A1(\u0.w[0][20] ),
    .A2(\u0.subword[20] ),
    .ZN(_07891_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16704_ (.A1(_07890_),
    .A2(_07786_),
    .A3(_07891_),
    .Z(_07892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16705_ (.I0(_07888_),
    .I1(_07889_),
    .S(_07892_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16706_ (.I(\u0.w[1][21] ),
    .ZN(_07893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16707_ (.I0(\u0.w[1][21] ),
    .I1(net199),
    .S(_07783_),
    .Z(_07894_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16708_ (.A1(\u0.w[0][21] ),
    .A2(\u0.subword[21] ),
    .Z(_07895_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16709_ (.A1(\u0.w[0][21] ),
    .A2(\u0.subword[21] ),
    .ZN(_07896_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16710_ (.A1(_07895_),
    .A2(_07733_),
    .A3(_07896_),
    .Z(_07897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16711_ (.I0(_07893_),
    .I1(_07894_),
    .S(_07897_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16712_ (.I0(\u0.w[1][22] ),
    .I1(net200),
    .S(_07806_),
    .Z(_07898_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16713_ (.I(\u0.w[1][22] ),
    .ZN(_07899_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16714_ (.A1(\u0.w[0][22] ),
    .A2(\u0.subword[22] ),
    .Z(_07900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16715_ (.A1(\u0.w[0][22] ),
    .A2(\u0.subword[22] ),
    .ZN(_07901_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16716_ (.A1(_07900_),
    .A2(_07835_),
    .A3(_07901_),
    .Z(_07902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16717_ (.I0(_07898_),
    .I1(_07899_),
    .S(_07902_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16718_ (.I0(\u0.w[1][23] ),
    .I1(net201),
    .S(_07783_),
    .Z(_07903_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16719_ (.I(\u0.w[1][23] ),
    .ZN(_07904_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16720_ (.A1(\u0.w[0][23] ),
    .A2(\u0.subword[23] ),
    .Z(_07905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16721_ (.A1(\u0.w[0][23] ),
    .A2(\u0.subword[23] ),
    .ZN(_07906_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16722_ (.A1(_07905_),
    .A2(_07835_),
    .A3(_07906_),
    .Z(_07907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16723_ (.I0(_07903_),
    .I1(_07904_),
    .S(_07907_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16724_ (.I(net697),
    .ZN(_07908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16725_ (.I0(net696),
    .I1(net202),
    .S(_07783_),
    .Z(_07909_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16726_ (.A1(\u0.w[0][24] ),
    .A2(\u0.subword[24] ),
    .A3(\u0.r0.out[24] ),
    .Z(_07910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16727_ (.I(_07835_),
    .Z(_07911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16728_ (.A1(_07910_),
    .A2(_07911_),
    .ZN(_07912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16729_ (.I0(_07908_),
    .I1(_07909_),
    .S(_07912_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16730_ (.I(net652),
    .ZN(_07913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16731_ (.I0(net653),
    .I1(net203),
    .S(_07783_),
    .Z(_07914_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16732_ (.A1(net629),
    .A2(\u0.subword[25] ),
    .A3(\u0.r0.out[25] ),
    .Z(_07915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16733_ (.A1(_07915_),
    .A2(_07911_),
    .ZN(_07916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16734_ (.I0(_07913_),
    .I1(_07914_),
    .S(_07916_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16735_ (.I(net766),
    .ZN(_07917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16736_ (.I0(net766),
    .I1(net205),
    .S(_07783_),
    .Z(_07918_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16737_ (.A1(\u0.w[0][26] ),
    .A2(\u0.subword[26] ),
    .A3(\u0.r0.out[26] ),
    .Z(_07919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16738_ (.A1(_07919_),
    .A2(_07911_),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16739_ (.I0(_07917_),
    .I1(_07918_),
    .S(_07920_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16740_ (.I(\u0.w[1][27] ),
    .ZN(_07921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16741_ (.I0(\u0.w[1][27] ),
    .I1(net206),
    .S(_07786_),
    .Z(_07922_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16742_ (.A1(\u0.w[0][27] ),
    .A2(\u0.subword[27] ),
    .A3(\u0.r0.out[27] ),
    .Z(_07923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16743_ (.A1(_07923_),
    .A2(_07793_),
    .ZN(_07924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16744_ (.I0(_07921_),
    .I1(_07922_),
    .S(_07924_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16745_ (.I(\u0.w[1][28] ),
    .ZN(_07925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16746_ (.I0(\u0.w[1][28] ),
    .I1(net207),
    .S(_07786_),
    .Z(_07926_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16747_ (.A1(\u0.w[0][28] ),
    .A2(\u0.subword[28] ),
    .A3(\u0.r0.out[28] ),
    .Z(_07927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16748_ (.A1(_07927_),
    .A2(_07793_),
    .ZN(_07928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16749_ (.I0(_07925_),
    .I1(_07926_),
    .S(_07928_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16750_ (.I(\u0.w[1][29] ),
    .ZN(_07929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16751_ (.I0(\u0.w[1][29] ),
    .I1(net208),
    .S(_07786_),
    .Z(_07930_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16752_ (.A1(\u0.w[0][29] ),
    .A2(\u0.subword[29] ),
    .A3(\u0.r0.out[29] ),
    .Z(_07931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16753_ (.A1(_07931_),
    .A2(_07793_),
    .ZN(_07932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16754_ (.I0(_07929_),
    .I1(_07930_),
    .S(_07932_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16755_ (.I0(\u0.w[1][30] ),
    .I1(net209),
    .S(_07786_),
    .Z(_07933_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16756_ (.A1(\u0.w[0][30] ),
    .A2(\u0.subword[30] ),
    .A3(\u0.r0.out[30] ),
    .Z(_07934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16757_ (.A1(_07934_),
    .A2(_07793_),
    .ZN(_07935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16758_ (.I0(_07729_),
    .I1(_07933_),
    .S(_07935_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16759_ (.I(\u0.w[1][31] ),
    .ZN(_07936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16760_ (.I0(\u0.w[1][31] ),
    .I1(net210),
    .S(_07786_),
    .Z(_07937_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16761_ (.A1(\u0.w[0][31] ),
    .A2(\u0.subword[31] ),
    .A3(\u0.r0.out[31] ),
    .Z(_07938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16762_ (.A1(_07938_),
    .A2(_07793_),
    .ZN(_07939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16763_ (.I0(_07936_),
    .I1(_07937_),
    .S(_07939_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16764_ (.I(_07746_),
    .Z(_07940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16765_ (.A1(_07940_),
    .A2(net211),
    .ZN(_07941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16766_ (.A1(_07788_),
    .A2(_07941_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16767_ (.I(_07733_),
    .Z(_07942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16768_ (.A1(_07942_),
    .A2(net212),
    .Z(_07943_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16769_ (.A1(_07795_),
    .A2(_07943_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16770_ (.A1(_07940_),
    .A2(net213),
    .ZN(_07944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16771_ (.A1(_07800_),
    .A2(_07944_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16772_ (.A1(_07940_),
    .A2(net214),
    .ZN(_07945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16773_ (.A1(_07805_),
    .A2(_07945_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16774_ (.A1(_07942_),
    .A2(net55),
    .Z(_07946_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16775_ (.A1(_07811_),
    .A2(_07946_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16776_ (.A1(_07942_),
    .A2(net56),
    .Z(_07947_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16777_ (.A1(_07814_),
    .A2(_07947_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16778_ (.I(_07733_),
    .Z(_07948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16779_ (.A1(_07948_),
    .A2(net65),
    .Z(_07949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16780_ (.A1(_07819_),
    .A2(_07949_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16781_ (.A1(_07940_),
    .A2(net67),
    .ZN(_07950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16782_ (.A1(_07824_),
    .A2(_07950_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16783_ (.A1(_07948_),
    .A2(net93),
    .Z(_07951_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16784_ (.A1(_07831_),
    .A2(_07951_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16785_ (.A1(_07948_),
    .A2(net94),
    .Z(_07952_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16786_ (.A1(_07837_),
    .A2(_07952_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16787_ (.A1(_07948_),
    .A2(net95),
    .Z(_07953_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16788_ (.A1(_07842_),
    .A2(_07953_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16789_ (.I(_07746_),
    .Z(_07954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16790_ (.A1(_07954_),
    .A2(net96),
    .ZN(_07955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16791_ (.A1(_07847_),
    .A2(_07955_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16792_ (.A1(_07948_),
    .A2(net97),
    .Z(_07956_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16793_ (.A1(_07852_),
    .A2(_07956_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16794_ (.A1(_07954_),
    .A2(net98),
    .ZN(_07957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16795_ (.A1(_07855_),
    .A2(_07957_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16796_ (.A1(_07954_),
    .A2(net100),
    .ZN(_07958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16797_ (.A1(_07860_),
    .A2(_07958_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16798_ (.A1(_07954_),
    .A2(net101),
    .ZN(_07959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16799_ (.A1(_07865_),
    .A2(_07959_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16800_ (.A1(_07948_),
    .A2(net102),
    .Z(_07960_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16801_ (.A1(_07872_),
    .A2(_07960_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16802_ (.A1(_07948_),
    .A2(net103),
    .Z(_07961_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16803_ (.A1(_07877_),
    .A2(_07961_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16804_ (.A1(_07948_),
    .A2(net104),
    .Z(_07962_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16805_ (.A1(_07882_),
    .A2(_07962_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16806_ (.A1(_07948_),
    .A2(net105),
    .Z(_07963_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16807_ (.A1(_07887_),
    .A2(_07963_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16808_ (.A1(_07954_),
    .A2(net106),
    .ZN(_07964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16809_ (.A1(_07892_),
    .A2(_07964_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16810_ (.A1(_07954_),
    .A2(net107),
    .ZN(_07965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16811_ (.A1(_07897_),
    .A2(_07965_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16812_ (.A1(_07948_),
    .A2(net108),
    .Z(_07966_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16813_ (.A1(_07902_),
    .A2(_07966_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16814_ (.A1(_07746_),
    .A2(net109),
    .Z(_07967_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16815_ (.A1(_07907_),
    .A2(_07967_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16816_ (.A1(_07954_),
    .A2(net111),
    .ZN(_07968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16817_ (.A1(_07912_),
    .A2(_07968_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16818_ (.A1(_07954_),
    .A2(net112),
    .ZN(_07969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16819_ (.A1(_07916_),
    .A2(_07969_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16820_ (.A1(_07954_),
    .A2(net113),
    .ZN(_07970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16821_ (.A1(_07920_),
    .A2(_07970_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16822_ (.A1(_07954_),
    .A2(net114),
    .ZN(_07971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16823_ (.A1(_07924_),
    .A2(_07971_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16824_ (.A1(_07747_),
    .A2(net115),
    .ZN(_07972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16825_ (.A1(_07928_),
    .A2(_07972_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16826_ (.A1(_07747_),
    .A2(net116),
    .ZN(_07973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16827_ (.A1(_07932_),
    .A2(_07973_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16828_ (.A1(_07747_),
    .A2(net117),
    .ZN(_07974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16829_ (.A1(_07935_),
    .A2(_07974_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16830_ (.A1(_07747_),
    .A2(net118),
    .ZN(_07975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16831_ (.A1(_07939_),
    .A2(_07975_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16832_ (.A1(_07466_),
    .A2(_07468_),
    .B(_07471_),
    .ZN(_15537_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16833_ (.I(_07536_),
    .ZN(_07976_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16834_ (.I(_07976_),
    .Z(_15557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16835_ (.A1(_07394_),
    .A2(_07468_),
    .B(_07448_),
    .ZN(_15538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16836_ (.I(_15553_),
    .ZN(_07977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16837_ (.A1(_15557_),
    .A2(_07977_),
    .ZN(_07978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16838_ (.I(_07978_),
    .ZN(_07979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16839_ (.I(_15549_),
    .ZN(_07980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16840_ (.A1(_15562_),
    .A2(_07980_),
    .ZN(_07981_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16841_ (.I(_07981_),
    .ZN(_07982_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16842_ (.A1(_07979_),
    .A2(_07982_),
    .B(_00390_),
    .ZN(_07983_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16843_ (.I(_07513_),
    .ZN(_07984_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16844_ (.I(_07984_),
    .Z(_07985_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16845_ (.I(_07985_),
    .Z(_07986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16846_ (.I(_15540_),
    .ZN(_07987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16847_ (.A1(_07536_),
    .A2(_07987_),
    .ZN(_07988_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16848_ (.I(_07319_),
    .Z(_07989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16849_ (.A1(_07988_),
    .A2(_07989_),
    .Z(_07990_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16850_ (.I(_07534_),
    .Z(_07991_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _16851_ (.I(_07535_),
    .Z(_07992_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16852_ (.A1(_07991_),
    .A2(_15539_),
    .A3(_07992_),
    .ZN(_07993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16853_ (.A1(_07990_),
    .A2(_07993_),
    .ZN(_07994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16854_ (.A1(_07983_),
    .A2(_07986_),
    .A3(_07994_),
    .ZN(_07995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16855_ (.A1(_07537_),
    .A2(_15538_),
    .ZN(_07996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16856_ (.A1(_07996_),
    .A2(_07989_),
    .Z(_07997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16857_ (.A1(net1038),
    .A2(net82),
    .ZN(_07998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16858_ (.A1(_07997_),
    .A2(_07998_),
    .ZN(_07999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16859_ (.A1(_07998_),
    .A2(_07996_),
    .ZN(_08000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16860_ (.I(_07330_),
    .Z(_08001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16861_ (.A1(_08000_),
    .A2(_08001_),
    .ZN(_08002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16862_ (.A1(_07999_),
    .A2(_08002_),
    .A3(_00391_),
    .ZN(_08003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16863_ (.A1(_07995_),
    .A2(_08003_),
    .A3(_00392_),
    .ZN(_08004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16864_ (.A1(_15557_),
    .A2(net6),
    .ZN(_08005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16865_ (.A1(_15562_),
    .A2(_15540_),
    .ZN(_08006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16866_ (.A1(_08005_),
    .A2(_08006_),
    .ZN(_08007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16867_ (.I(_07319_),
    .Z(_08008_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16868_ (.I(_08008_),
    .Z(_08009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16869_ (.A1(_08007_),
    .A2(_08009_),
    .ZN(_08010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16870_ (.A1(_07987_),
    .A2(_07992_),
    .A3(_07991_),
    .ZN(_08011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16871_ (.I(_08011_),
    .ZN(_08012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16872_ (.A1(_07341_),
    .A2(_08012_),
    .ZN(_08013_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16873_ (.A1(_08010_),
    .A2(_00391_),
    .A3(_08013_),
    .ZN(_08014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16874_ (.A1(_07537_),
    .A2(_07977_),
    .ZN(_08015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16875_ (.I(_08015_),
    .ZN(_08016_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16876_ (.I(_07989_),
    .Z(_08017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16877_ (.I(_07513_),
    .Z(_08018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16878_ (.A1(_08016_),
    .A2(_08017_),
    .B(_08018_),
    .ZN(_08019_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16879_ (.A1(_07991_),
    .A2(_15553_),
    .A3(_07992_),
    .ZN(_08020_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16880_ (.I(_07341_),
    .Z(_08021_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16881_ (.A1(net61),
    .A2(_08020_),
    .A3(_08021_),
    .ZN(_08022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16882_ (.A1(_15557_),
    .A2(_07980_),
    .ZN(_08023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16883_ (.I(_08023_),
    .ZN(_08024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16884_ (.A1(_08024_),
    .A2(_08017_),
    .ZN(_08025_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16885_ (.A1(_08019_),
    .A2(_08022_),
    .A3(_08025_),
    .ZN(_08026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16886_ (.I(_07484_),
    .ZN(_08027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16887_ (.I(_08027_),
    .Z(_08028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16888_ (.A1(_08014_),
    .A2(_08026_),
    .A3(_08028_),
    .ZN(_08029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16889_ (.I(_07666_),
    .ZN(_08030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16890_ (.I(_08030_),
    .Z(_08031_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16891_ (.A1(_08004_),
    .A2(_08029_),
    .A3(_08031_),
    .ZN(_08032_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16892_ (.A1(_07537_),
    .A2(_15537_),
    .ZN(_08033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16893_ (.A1(_08033_),
    .A2(_08008_),
    .ZN(_08034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16894_ (.I(_07984_),
    .Z(_08035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16895_ (.A1(_08034_),
    .A2(_08035_),
    .Z(_08036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16896_ (.A1(_07976_),
    .A2(net1037),
    .ZN(_08037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16897_ (.A1(_07537_),
    .A2(_15539_),
    .ZN(_08038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16898_ (.A1(_08037_),
    .A2(_07341_),
    .A3(_08038_),
    .ZN(_08039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16899_ (.A1(_07537_),
    .A2(_15555_),
    .Z(_08040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16900_ (.A1(_08040_),
    .A2(_08008_),
    .ZN(_08041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16901_ (.A1(_08036_),
    .A2(_08039_),
    .A3(_08041_),
    .ZN(_08042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16902_ (.I(_15541_),
    .ZN(_08043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16903_ (.A1(_15562_),
    .A2(_08043_),
    .ZN(_08044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16904_ (.A1(_08044_),
    .A2(_07341_),
    .Z(_08045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16905_ (.A1(_08045_),
    .A2(_08037_),
    .ZN(_08046_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16906_ (.I(_08018_),
    .Z(_08047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16907_ (.A1(_15548_),
    .A2(_07537_),
    .ZN(_08048_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16908_ (.I(_08008_),
    .Z(_08049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16909_ (.A1(_07991_),
    .A2(_15544_),
    .A3(_07992_),
    .ZN(_08050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16910_ (.A1(_08048_),
    .A2(_08049_),
    .A3(_08050_),
    .ZN(_08051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16911_ (.A1(_08046_),
    .A2(_08047_),
    .A3(_08051_),
    .ZN(_08052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16912_ (.A1(_08042_),
    .A2(_08052_),
    .A3(_08028_),
    .ZN(_08053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16913_ (.A1(_08050_),
    .A2(_07319_),
    .ZN(_08054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16914_ (.I(_08054_),
    .ZN(_08055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16915_ (.A1(net1036),
    .A2(_07537_),
    .ZN(_08056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16916_ (.A1(_08055_),
    .A2(_08056_),
    .ZN(_08057_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16917_ (.A1(_08043_),
    .A2(_07534_),
    .A3(_07535_),
    .ZN(_08058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16918_ (.A1(_08058_),
    .A2(_07330_),
    .ZN(_08059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16919_ (.I(_08059_),
    .ZN(_08060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16920_ (.A1(_08060_),
    .A2(net61),
    .ZN(_08061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16921_ (.A1(_08057_),
    .A2(_08061_),
    .A3(_08047_),
    .ZN(_08062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16922_ (.I(_07330_),
    .Z(_08063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16923_ (.A1(_08050_),
    .A2(_08063_),
    .ZN(_08064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16924_ (.I(_08064_),
    .ZN(_08065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16925_ (.I(_15546_),
    .ZN(_08066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16926_ (.A1(_15562_),
    .A2(_08066_),
    .ZN(_08067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16927_ (.A1(_08065_),
    .A2(_08067_),
    .ZN(_08068_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16928_ (.I(_08035_),
    .Z(_08069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16929_ (.A1(_08037_),
    .A2(_07989_),
    .ZN(_08070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16930_ (.A1(_08068_),
    .A2(_08069_),
    .A3(_08070_),
    .ZN(_08071_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16931_ (.I(_07484_),
    .Z(_08072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16932_ (.A1(_08062_),
    .A2(_08071_),
    .A3(_08072_),
    .ZN(_08073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16933_ (.A1(_08053_),
    .A2(_08073_),
    .A3(_00393_),
    .ZN(_08074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16934_ (.I(_00394_),
    .ZN(_08075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16935_ (.I(_08075_),
    .Z(_08076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16936_ (.A1(_08032_),
    .A2(_08074_),
    .A3(_08076_),
    .ZN(_08077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16937_ (.A1(_07979_),
    .A2(_08040_),
    .B(_08017_),
    .ZN(_08078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16938_ (.A1(_08067_),
    .A2(_08063_),
    .Z(_08079_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16939_ (.I(_08035_),
    .Z(_08080_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16940_ (.A1(_08079_),
    .A2(_08080_),
    .ZN(_08081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16941_ (.I(_08027_),
    .Z(_08082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16942_ (.A1(_08078_),
    .A2(_08081_),
    .B(_08082_),
    .ZN(_08083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16943_ (.A1(_07537_),
    .A2(_15537_),
    .ZN(_08084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16944_ (.A1(_08084_),
    .A2(_07989_),
    .Z(_08085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16945_ (.A1(_07991_),
    .A2(_07992_),
    .A3(_15540_),
    .ZN(_08086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16946_ (.A1(_08085_),
    .A2(_08086_),
    .ZN(_08087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16947_ (.A1(_07991_),
    .A2(_15549_),
    .A3(_07992_),
    .ZN(_08088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16948_ (.A1(_08056_),
    .A2(_08021_),
    .A3(_08088_),
    .ZN(_08089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16949_ (.A1(_08087_),
    .A2(_08069_),
    .A3(_08089_),
    .ZN(_08090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16950_ (.I(_08030_),
    .Z(_08091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16951_ (.A1(_08083_),
    .A2(_08090_),
    .B(_08091_),
    .ZN(_08092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16952_ (.A1(_07330_),
    .A2(_07988_),
    .ZN(_08093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16953_ (.I(_08093_),
    .ZN(_08094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _16954_ (.I(_15551_),
    .ZN(_08095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16955_ (.A1(_07991_),
    .A2(_07992_),
    .B(_08095_),
    .ZN(_08096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16956_ (.A1(_08008_),
    .A2(_08096_),
    .Z(_08097_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16957_ (.A1(_08094_),
    .A2(_08097_),
    .A3(_08080_),
    .ZN(_08098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16958_ (.A1(_08039_),
    .A2(_08035_),
    .Z(_08099_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16959_ (.A1(_07991_),
    .A2(_15546_),
    .A3(_07992_),
    .ZN(_08100_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16960_ (.A1(_08063_),
    .A2(_08100_),
    .Z(_08101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16961_ (.A1(_08099_),
    .A2(_08098_),
    .B(_08101_),
    .ZN(_08102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16962_ (.A1(_08102_),
    .A2(_08028_),
    .ZN(_08103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16963_ (.A1(_08103_),
    .A2(_08092_),
    .ZN(_08104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16964_ (.I(_15544_),
    .ZN(_08105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16965_ (.A1(_15562_),
    .A2(_08105_),
    .Z(_08106_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16966_ (.I(_07319_),
    .Z(_08107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16967_ (.A1(_08106_),
    .A2(_08107_),
    .B(_08035_),
    .ZN(_08108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16968_ (.A1(_08040_),
    .A2(_08063_),
    .ZN(_08109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16969_ (.A1(_08108_),
    .A2(_08025_),
    .A3(_08109_),
    .ZN(_08110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16970_ (.A1(_07991_),
    .A2(_07992_),
    .A3(_08095_),
    .ZN(_08111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16971_ (.A1(_07330_),
    .A2(_08111_),
    .ZN(_08112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16972_ (.I(_08112_),
    .ZN(_08113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16973_ (.A1(_07537_),
    .A2(_15544_),
    .ZN(_08114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16974_ (.A1(_08114_),
    .A2(_08113_),
    .ZN(_08115_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16975_ (.I(_08035_),
    .Z(_08116_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16976_ (.A1(_08041_),
    .A2(_08116_),
    .A3(_08115_),
    .ZN(_08117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16977_ (.A1(_08110_),
    .A2(_08117_),
    .A3(_08072_),
    .ZN(_08118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16978_ (.A1(_15562_),
    .A2(_15553_),
    .ZN(_08119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16979_ (.A1(_08037_),
    .A2(_08001_),
    .A3(_08119_),
    .ZN(_08120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16980_ (.A1(_15557_),
    .A2(net5),
    .ZN(_08121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16981_ (.A1(_08121_),
    .A2(_08049_),
    .A3(_08114_),
    .ZN(_08122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16982_ (.A1(_08120_),
    .A2(_08122_),
    .A3(_08116_),
    .ZN(_08123_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16983_ (.I(_08027_),
    .Z(_08124_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _16984_ (.I(_08063_),
    .Z(_08125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16985_ (.A1(_08125_),
    .A2(_15565_),
    .ZN(_08126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _16986_ (.I(_07513_),
    .Z(_08127_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16987_ (.A1(_00390_),
    .A2(_08086_),
    .B(_08126_),
    .C(_08127_),
    .ZN(_08128_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16988_ (.A1(_08123_),
    .A2(_08124_),
    .A3(_08128_),
    .ZN(_08129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16989_ (.A1(_08031_),
    .A2(_08129_),
    .A3(_08118_),
    .ZN(_08130_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16990_ (.A1(_08104_),
    .A2(_08130_),
    .A3(_00394_),
    .ZN(_08131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16991_ (.A1(_08077_),
    .A2(_08131_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16992_ (.A1(_08056_),
    .A2(_08008_),
    .Z(_08132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16993_ (.A1(_08132_),
    .A2(_08020_),
    .ZN(_08133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16994_ (.A1(_08065_),
    .A2(_08038_),
    .ZN(_08134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16995_ (.A1(_08133_),
    .A2(_08072_),
    .A3(_08134_),
    .ZN(_08135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16996_ (.A1(_08135_),
    .A2(_00391_),
    .ZN(_08136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16997_ (.A1(_07997_),
    .A2(_08005_),
    .ZN(_08137_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16998_ (.I(_08033_),
    .ZN(_08138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16999_ (.A1(_08079_),
    .A2(_08138_),
    .ZN(_08139_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17000_ (.A1(_08137_),
    .A2(_08139_),
    .A3(_08124_),
    .Z(_08140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17001_ (.A1(_08088_),
    .A2(_07319_),
    .ZN(_08141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17002_ (.I(_08141_),
    .ZN(_08142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17003_ (.A1(_08142_),
    .A2(_08038_),
    .ZN(_08143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17004_ (.I(_08143_),
    .ZN(_08144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17005_ (.I(_15567_),
    .ZN(_08145_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17006_ (.A1(_08027_),
    .A2(_08145_),
    .A3(_08125_),
    .Z(_08146_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17007_ (.A1(_08144_),
    .A2(_08146_),
    .B(_07986_),
    .ZN(_08147_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17008_ (.A1(_08136_),
    .A2(_08140_),
    .B(_08031_),
    .C(_08147_),
    .ZN(_08148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17009_ (.I(_08121_),
    .ZN(_08149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17010_ (.A1(_08149_),
    .A2(_08107_),
    .ZN(_08150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17011_ (.A1(_08150_),
    .A2(_08041_),
    .Z(_08151_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17012_ (.I(_08086_),
    .ZN(_08152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17013_ (.A1(_08152_),
    .A2(_07341_),
    .ZN(_08153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17014_ (.A1(_08153_),
    .A2(_07513_),
    .Z(_08154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17015_ (.A1(_08016_),
    .A2(_08001_),
    .ZN(_08155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17016_ (.A1(_08151_),
    .A2(_08154_),
    .A3(_08155_),
    .ZN(_08156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17017_ (.A1(_07997_),
    .A2(_08020_),
    .ZN(_08157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17018_ (.A1(_08157_),
    .A2(_08139_),
    .A3(_08069_),
    .ZN(_08158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17019_ (.A1(_08156_),
    .A2(_00392_),
    .A3(_08158_),
    .ZN(_08159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17020_ (.A1(_08121_),
    .A2(_07985_),
    .ZN(_08160_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17021_ (.A1(_08094_),
    .A2(_08160_),
    .ZN(_08161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17022_ (.I(_15539_),
    .ZN(_08162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17023_ (.A1(_15562_),
    .A2(_08162_),
    .ZN(_08163_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17024_ (.A1(_08163_),
    .A2(_08001_),
    .Z(_08164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17025_ (.A1(_08161_),
    .A2(_08164_),
    .B(_07486_),
    .ZN(_08165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17026_ (.A1(_08044_),
    .A2(_08008_),
    .ZN(_08166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17027_ (.I(_08166_),
    .ZN(_08167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17028_ (.A1(_15562_),
    .A2(_15555_),
    .Z(_08168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17029_ (.A1(_08167_),
    .A2(_08168_),
    .ZN(_08169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17030_ (.A1(_07993_),
    .A2(_08063_),
    .ZN(_08170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17031_ (.I(_08170_),
    .ZN(_08171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17032_ (.A1(_08171_),
    .A2(_08006_),
    .ZN(_08172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17033_ (.A1(_08169_),
    .A2(_08172_),
    .A3(_08047_),
    .ZN(_08173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17034_ (.A1(_08165_),
    .A2(_08173_),
    .B(_08091_),
    .ZN(_08174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17035_ (.A1(_08159_),
    .A2(_08174_),
    .ZN(_08175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17036_ (.A1(_08148_),
    .A2(_08175_),
    .A3(_08076_),
    .ZN(_08176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17037_ (.A1(_15562_),
    .A2(_15546_),
    .Z(_08177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17038_ (.A1(_08177_),
    .A2(_08049_),
    .B(_08018_),
    .ZN(_08178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17039_ (.A1(_08178_),
    .A2(_08172_),
    .B(_08082_),
    .ZN(_08179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17040_ (.A1(_08060_),
    .A2(_08048_),
    .ZN(_08180_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17041_ (.A1(_08180_),
    .A2(_08047_),
    .A3(_08164_),
    .ZN(_08181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17042_ (.A1(_08179_),
    .A2(_08181_),
    .B(_08091_),
    .ZN(_08182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17043_ (.A1(_07997_),
    .A2(net896),
    .ZN(_08183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17044_ (.A1(net5),
    .A2(net6),
    .ZN(_08184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17045_ (.A1(_08056_),
    .A2(_08184_),
    .A3(_08125_),
    .ZN(_08185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17046_ (.A1(_08183_),
    .A2(_08080_),
    .A3(_08185_),
    .ZN(_08186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17047_ (.A1(_08094_),
    .A2(_08100_),
    .ZN(_08187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17048_ (.A1(_08121_),
    .A2(_08107_),
    .A3(_08015_),
    .ZN(_08188_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17049_ (.A1(_08187_),
    .A2(_08188_),
    .A3(_08127_),
    .ZN(_08189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17050_ (.A1(_08189_),
    .A2(_08186_),
    .ZN(_08190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17051_ (.A1(_08190_),
    .A2(_08028_),
    .ZN(_08191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17052_ (.A1(_08191_),
    .A2(_08182_),
    .B(_08076_),
    .ZN(_08192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17053_ (.I(_08037_),
    .ZN(_08193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17054_ (.A1(_08067_),
    .A2(_08008_),
    .ZN(_08194_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17055_ (.A1(_08193_),
    .A2(_08093_),
    .B1(_08194_),
    .B2(_08149_),
    .ZN(_08195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17056_ (.A1(_08085_),
    .A2(_07998_),
    .ZN(_08196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17057_ (.A1(_08063_),
    .A2(_15557_),
    .Z(_08197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17058_ (.A1(_08197_),
    .A2(_08105_),
    .ZN(_08198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17059_ (.A1(_08196_),
    .A2(_08116_),
    .A3(_08198_),
    .ZN(_08199_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17060_ (.A1(_08195_),
    .A2(_07986_),
    .B(_08199_),
    .C(_08072_),
    .ZN(_08200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17061_ (.A1(_07989_),
    .A2(net82),
    .ZN(_08201_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17062_ (.A1(_08201_),
    .A2(_15557_),
    .Z(_08202_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17063_ (.A1(_07989_),
    .A2(_15558_),
    .Z(_08203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17064_ (.A1(_08202_),
    .A2(_08203_),
    .Z(_08204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17065_ (.A1(_08101_),
    .A2(_07513_),
    .Z(_08205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17066_ (.A1(_08204_),
    .A2(_08205_),
    .B(_07486_),
    .ZN(_08206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17067_ (.A1(_08106_),
    .A2(_08107_),
    .ZN(_08207_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17068_ (.A1(_08207_),
    .A2(_08035_),
    .A3(_08101_),
    .Z(_08208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17069_ (.A1(_08045_),
    .A2(_08011_),
    .ZN(_08209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17070_ (.A1(_08208_),
    .A2(_08209_),
    .ZN(_08210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17071_ (.A1(_08206_),
    .A2(_08210_),
    .B(_00393_),
    .ZN(_08211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17072_ (.A1(_08200_),
    .A2(_08211_),
    .ZN(_08212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17073_ (.A1(_08212_),
    .A2(_08192_),
    .ZN(_08213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17074_ (.A1(_08176_),
    .A2(_08213_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17075_ (.A1(_08056_),
    .A2(_07989_),
    .A3(_08111_),
    .Z(_08214_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17076_ (.A1(_07988_),
    .A2(_08001_),
    .A3(_08086_),
    .Z(_08215_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17077_ (.A1(_08214_),
    .A2(_08215_),
    .B(_08080_),
    .ZN(_08216_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17078_ (.I(_08096_),
    .ZN(_08217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17079_ (.A1(_08138_),
    .A2(_08217_),
    .A3(_08125_),
    .ZN(_08218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17080_ (.A1(_07991_),
    .A2(_15541_),
    .A3(_07992_),
    .ZN(_08219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17081_ (.A1(_07996_),
    .A2(_08107_),
    .A3(_08219_),
    .ZN(_08220_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17082_ (.A1(_08218_),
    .A2(_08127_),
    .A3(_08220_),
    .ZN(_08221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17083_ (.A1(_08216_),
    .A2(_08221_),
    .ZN(_08222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17084_ (.A1(_08222_),
    .A2(_00392_),
    .ZN(_08223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17085_ (.A1(_08217_),
    .A2(_08100_),
    .ZN(_08224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17086_ (.A1(_08224_),
    .A2(_08009_),
    .ZN(_08225_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17087_ (.A1(_15557_),
    .A2(_08066_),
    .ZN(_08226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17088_ (.A1(_08226_),
    .A2(_08021_),
    .A3(_08048_),
    .ZN(_08227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17089_ (.A1(_08225_),
    .A2(_08227_),
    .A3(_08069_),
    .ZN(_08228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17090_ (.A1(_08096_),
    .A2(_08049_),
    .B(_07985_),
    .ZN(_08229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17091_ (.A1(_08226_),
    .A2(_08021_),
    .A3(_08056_),
    .ZN(_08230_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17092_ (.A1(_08219_),
    .A2(_08001_),
    .Z(_08231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17093_ (.A1(_08229_),
    .A2(_08230_),
    .A3(_08231_),
    .ZN(_08232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17094_ (.A1(_08228_),
    .A2(_08232_),
    .A3(_08124_),
    .ZN(_08233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17095_ (.A1(_08223_),
    .A2(_00393_),
    .A3(_08233_),
    .ZN(_08234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17096_ (.I(_08087_),
    .ZN(_08235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17097_ (.A1(_08100_),
    .A2(_08063_),
    .ZN(_08236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17098_ (.A1(_08236_),
    .A2(_08106_),
    .B(_08035_),
    .ZN(_08237_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17099_ (.A1(_08235_),
    .A2(_08237_),
    .ZN(_08238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17100_ (.A1(_08065_),
    .A2(_08084_),
    .ZN(_08239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17101_ (.A1(_08067_),
    .A2(_08058_),
    .A3(_08017_),
    .ZN(_08240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17102_ (.A1(_08239_),
    .A2(_08240_),
    .B(_08116_),
    .ZN(_08241_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17103_ (.A1(_08238_),
    .A2(_08241_),
    .B(_08124_),
    .ZN(_08242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17104_ (.A1(_15557_),
    .A2(_15555_),
    .ZN(_08243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17105_ (.I(_08243_),
    .ZN(_08244_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17106_ (.I(_07996_),
    .ZN(_08245_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17107_ (.A1(_08244_),
    .A2(_08245_),
    .B(_08021_),
    .ZN(_08246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17108_ (.A1(_08005_),
    .A2(_08049_),
    .A3(net61),
    .ZN(_08247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17109_ (.A1(_08246_),
    .A2(_00391_),
    .A3(_08247_),
    .ZN(_08248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17110_ (.A1(_08054_),
    .A2(_08035_),
    .Z(_08249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17111_ (.A1(_08171_),
    .A2(_08044_),
    .ZN(_08250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17112_ (.A1(_08249_),
    .A2(_08250_),
    .B(_08082_),
    .ZN(_08251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17113_ (.A1(_08248_),
    .A2(_08251_),
    .ZN(_08252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17114_ (.A1(_08242_),
    .A2(_08031_),
    .A3(_08252_),
    .ZN(_08253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17115_ (.A1(_08234_),
    .A2(_08253_),
    .A3(_08076_),
    .ZN(_08254_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17116_ (.A1(_08245_),
    .A2(_15560_),
    .B(_08125_),
    .ZN(_08255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17117_ (.A1(_08087_),
    .A2(_08255_),
    .B(_08116_),
    .ZN(_08256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17118_ (.A1(_08114_),
    .A2(_07341_),
    .ZN(_08257_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17119_ (.A1(_08012_),
    .A2(_08257_),
    .Z(_08258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17120_ (.A1(_08017_),
    .A2(_15565_),
    .ZN(_08259_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17121_ (.I(_07513_),
    .Z(_08260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17122_ (.A1(_08259_),
    .A2(_08258_),
    .B(_08260_),
    .ZN(_08261_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17123_ (.A1(_08261_),
    .A2(_08256_),
    .B(_00393_),
    .ZN(_08262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17124_ (.A1(_08094_),
    .A2(_08226_),
    .ZN(_08263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17125_ (.A1(_08263_),
    .A2(_08019_),
    .B(_07666_),
    .ZN(_08264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17126_ (.A1(_08171_),
    .A2(_07996_),
    .ZN(_08265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17127_ (.A1(_08143_),
    .A2(_08265_),
    .A3(_08260_),
    .ZN(_08266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17128_ (.A1(_08264_),
    .A2(_08266_),
    .B(_08124_),
    .ZN(_08267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17129_ (.A1(_08267_),
    .A2(_08262_),
    .ZN(_08268_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17130_ (.A1(_08107_),
    .A2(_15563_),
    .Z(_08269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17131_ (.A1(_08269_),
    .A2(_08249_),
    .B(_07666_),
    .ZN(_08270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17132_ (.A1(_08049_),
    .A2(_15560_),
    .ZN(_08271_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17133_ (.A1(_08239_),
    .A2(_08260_),
    .A3(_08271_),
    .ZN(_08272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17134_ (.A1(_08270_),
    .A2(_08272_),
    .B(_08072_),
    .ZN(_08273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17135_ (.A1(_07978_),
    .A2(_08084_),
    .ZN(_08274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17136_ (.A1(_08274_),
    .A2(_08009_),
    .ZN(_08275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17137_ (.A1(_07982_),
    .A2(_00390_),
    .ZN(_08276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17138_ (.A1(_08154_),
    .A2(_08275_),
    .A3(_08276_),
    .ZN(_08277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17139_ (.A1(_07998_),
    .A2(_08084_),
    .A3(_08125_),
    .ZN(_08278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17140_ (.A1(_08049_),
    .A2(_08145_),
    .ZN(_08279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17141_ (.A1(_08278_),
    .A2(_08116_),
    .A3(_08279_),
    .ZN(_08280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17142_ (.A1(_08277_),
    .A2(_00393_),
    .A3(_08280_),
    .ZN(_08281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17143_ (.A1(_08273_),
    .A2(_08281_),
    .ZN(_08282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17144_ (.A1(_08268_),
    .A2(_00394_),
    .A3(_08282_),
    .ZN(_08283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17145_ (.A1(_08283_),
    .A2(_08254_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17146_ (.I(_08214_),
    .ZN(_08284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17147_ (.A1(_08096_),
    .A2(_08001_),
    .ZN(_08285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17148_ (.A1(_08284_),
    .A2(_07486_),
    .A3(_08285_),
    .ZN(_08286_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17149_ (.I(_08070_),
    .ZN(_08287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17150_ (.A1(_08287_),
    .A2(_07988_),
    .ZN(_08288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17151_ (.A1(_08060_),
    .A2(_07996_),
    .ZN(_08289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17152_ (.A1(_08288_),
    .A2(_08027_),
    .A3(_08289_),
    .ZN(_08290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17153_ (.A1(_08286_),
    .A2(_08290_),
    .ZN(_08291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17154_ (.A1(_08291_),
    .A2(_07986_),
    .ZN(_08292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17155_ (.A1(_08142_),
    .A2(_08084_),
    .Z(_08293_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17156_ (.I(_08013_),
    .ZN(_08294_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17157_ (.A1(_08293_),
    .A2(_08294_),
    .B(_08027_),
    .ZN(_08295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17158_ (.A1(_08109_),
    .A2(_07513_),
    .Z(_08296_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17159_ (.A1(_08027_),
    .A2(_07988_),
    .A3(_08063_),
    .Z(_08297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17160_ (.A1(_08296_),
    .A2(_08297_),
    .Z(_08298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17161_ (.A1(_08295_),
    .A2(_08298_),
    .B(_07666_),
    .ZN(_08299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17162_ (.A1(_08292_),
    .A2(_08299_),
    .ZN(_08300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17163_ (.A1(_08193_),
    .A2(_08096_),
    .B(_07341_),
    .ZN(_08301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17164_ (.A1(_07990_),
    .A2(_08058_),
    .ZN(_08302_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17165_ (.A1(_08301_),
    .A2(_08127_),
    .A3(_08302_),
    .ZN(_08303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17166_ (.A1(_08196_),
    .A2(_08120_),
    .A3(_07985_),
    .ZN(_08304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17167_ (.A1(_08303_),
    .A2(_08304_),
    .ZN(_08305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17168_ (.A1(_08305_),
    .A2(_08072_),
    .ZN(_08306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17169_ (.A1(_08113_),
    .A2(_07996_),
    .ZN(_08307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17170_ (.A1(_08143_),
    .A2(_08307_),
    .ZN(_08308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17171_ (.A1(_08308_),
    .A2(_08080_),
    .ZN(_08309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17172_ (.A1(_08220_),
    .A2(_08127_),
    .B(_07486_),
    .ZN(_08310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17173_ (.A1(_08309_),
    .A2(_08310_),
    .B(_08091_),
    .ZN(_08311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17174_ (.A1(_08306_),
    .A2(_08311_),
    .ZN(_08312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17175_ (.A1(_08300_),
    .A2(_08312_),
    .ZN(_08313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17176_ (.A1(_08313_),
    .A2(_08076_),
    .ZN(_08314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17177_ (.A1(_08038_),
    .A2(_07989_),
    .Z(_08315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17178_ (.A1(_08315_),
    .A2(_08011_),
    .ZN(_08316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17179_ (.A1(_15557_),
    .A2(_08105_),
    .ZN(_08317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17180_ (.A1(_08317_),
    .A2(_07981_),
    .ZN(_08318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17181_ (.A1(_08318_),
    .A2(_08001_),
    .ZN(_08319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17182_ (.A1(_08316_),
    .A2(_08319_),
    .ZN(_08320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17183_ (.A1(_08320_),
    .A2(_08080_),
    .ZN(_08321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17184_ (.A1(_07990_),
    .A2(_08023_),
    .ZN(_08322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17185_ (.A1(_08322_),
    .A2(_08002_),
    .A3(_08127_),
    .ZN(_08323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17186_ (.A1(_08321_),
    .A2(_08323_),
    .ZN(_08324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17187_ (.A1(_08324_),
    .A2(_00392_),
    .ZN(_08325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17188_ (.A1(_08121_),
    .A2(_07998_),
    .ZN(_08326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17189_ (.A1(_08326_),
    .A2(_08017_),
    .ZN(_08327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17190_ (.A1(_08064_),
    .A2(_07985_),
    .Z(_08328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17191_ (.A1(_08327_),
    .A2(_08328_),
    .B(_07486_),
    .ZN(_08329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17192_ (.A1(_08111_),
    .A2(_07319_),
    .ZN(_08330_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17193_ (.I(_08330_),
    .ZN(_08331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17194_ (.A1(_08331_),
    .A2(_08006_),
    .ZN(_08332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17195_ (.A1(_08180_),
    .A2(_08332_),
    .A3(_08260_),
    .ZN(_08333_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17196_ (.A1(_08329_),
    .A2(_08333_),
    .B(_08091_),
    .ZN(_08334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17197_ (.A1(_08325_),
    .A2(_08334_),
    .B(_08075_),
    .ZN(_08335_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17198_ (.A1(_08155_),
    .A2(_08018_),
    .Z(_08336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17199_ (.A1(_08149_),
    .A2(_07982_),
    .B(_08049_),
    .ZN(_08337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17200_ (.A1(_08336_),
    .A2(_08337_),
    .A3(_08013_),
    .ZN(_08338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17201_ (.I(_08006_),
    .ZN(_08339_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17202_ (.A1(_08339_),
    .A2(_08001_),
    .A3(_08033_),
    .Z(_08340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17203_ (.A1(_08045_),
    .A2(_08226_),
    .ZN(_08341_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17204_ (.A1(_08340_),
    .A2(_08069_),
    .A3(_08341_),
    .ZN(_08342_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17205_ (.A1(_08338_),
    .A2(_08342_),
    .A3(_00392_),
    .ZN(_08343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17206_ (.A1(_08094_),
    .A2(_08138_),
    .ZN(_08344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17207_ (.A1(_08327_),
    .A2(_08344_),
    .B(_08260_),
    .ZN(_08345_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17208_ (.A1(_08245_),
    .A2(_15560_),
    .ZN(_08346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17209_ (.A1(_08127_),
    .A2(_08013_),
    .ZN(_08347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17210_ (.A1(_08009_),
    .A2(_08346_),
    .B(_08347_),
    .ZN(_08348_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17211_ (.A1(_08348_),
    .A2(_08345_),
    .B(_08124_),
    .ZN(_08349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17212_ (.A1(_08343_),
    .A2(_08031_),
    .A3(_08349_),
    .ZN(_08350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17213_ (.A1(_08335_),
    .A2(_08350_),
    .ZN(_08351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17214_ (.A1(_08351_),
    .A2(_08314_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17215_ (.A1(_08078_),
    .A2(_07986_),
    .A3(_08002_),
    .ZN(_08352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17216_ (.A1(_08048_),
    .A2(_08184_),
    .ZN(_08353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17217_ (.A1(_08353_),
    .A2(_08009_),
    .ZN(_08354_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17218_ (.A1(_08354_),
    .A2(_08307_),
    .A3(_08047_),
    .ZN(_08355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17219_ (.A1(_08352_),
    .A2(_08028_),
    .A3(_08355_),
    .ZN(_08356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17220_ (.A1(_08113_),
    .A2(_08048_),
    .ZN(_08357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17221_ (.A1(_08108_),
    .A2(_08357_),
    .ZN(_08358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17222_ (.A1(_08017_),
    .A2(_08162_),
    .ZN(_08359_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17223_ (.A1(_08152_),
    .A2(_08009_),
    .B(_08080_),
    .C(_08359_),
    .ZN(_08360_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17224_ (.A1(_08358_),
    .A2(_08360_),
    .A3(_00392_),
    .ZN(_08361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17225_ (.A1(_08356_),
    .A2(_08031_),
    .A3(_08361_),
    .ZN(_08362_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17226_ (.A1(_08194_),
    .A2(_08152_),
    .Z(_08363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17227_ (.A1(_08099_),
    .A2(_08363_),
    .ZN(_08364_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17228_ (.A1(_08170_),
    .A2(_08018_),
    .Z(_08365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17229_ (.A1(_08168_),
    .A2(_08008_),
    .ZN(_08366_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17230_ (.A1(_08365_),
    .A2(_08366_),
    .B(_08082_),
    .ZN(_08367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17231_ (.A1(_08364_),
    .A2(_08367_),
    .ZN(_08368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17232_ (.A1(_07997_),
    .A2(_08058_),
    .ZN(_08369_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17233_ (.A1(_08197_),
    .A2(_08127_),
    .ZN(_08370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17234_ (.A1(_08369_),
    .A2(_08370_),
    .B(_07486_),
    .ZN(_08371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17235_ (.A1(_08016_),
    .A2(_08017_),
    .B(_07985_),
    .ZN(_08372_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17236_ (.A1(_08139_),
    .A2(_08372_),
    .A3(_08034_),
    .ZN(_08373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17237_ (.A1(_08371_),
    .A2(_08373_),
    .ZN(_08374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17238_ (.A1(_08368_),
    .A2(_08374_),
    .A3(_00393_),
    .ZN(_08375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17239_ (.A1(_08362_),
    .A2(_08076_),
    .A3(_08375_),
    .ZN(_08376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17240_ (.A1(_08005_),
    .A2(_08015_),
    .ZN(_08377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17241_ (.A1(_08377_),
    .A2(_00390_),
    .ZN(_08378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17242_ (.A1(_08208_),
    .A2(_08378_),
    .ZN(_08379_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17243_ (.A1(_08033_),
    .A2(_08257_),
    .B(_08240_),
    .C(_08260_),
    .ZN(_08380_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17244_ (.A1(_08379_),
    .A2(_08380_),
    .A3(_08028_),
    .ZN(_08381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17245_ (.A1(_08153_),
    .A2(_08217_),
    .Z(_08382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17246_ (.A1(_08205_),
    .A2(_08382_),
    .B(_08082_),
    .ZN(_08383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17247_ (.A1(_08167_),
    .A2(_08011_),
    .ZN(_08384_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17248_ (.A1(_08384_),
    .A2(_08115_),
    .A3(_08069_),
    .ZN(_08385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17249_ (.A1(_08383_),
    .A2(_08385_),
    .B(_00393_),
    .ZN(_08386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17250_ (.A1(_08381_),
    .A2(_08386_),
    .ZN(_08387_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17251_ (.A1(_08245_),
    .A2(_15569_),
    .B(_08125_),
    .ZN(_08388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17252_ (.A1(_08133_),
    .A2(_08388_),
    .A3(_08069_),
    .ZN(_08389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17253_ (.A1(_08040_),
    .A2(_07985_),
    .ZN(_08390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17254_ (.A1(_08390_),
    .A2(_08112_),
    .B(_08027_),
    .ZN(_08391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17255_ (.A1(_08389_),
    .A2(_08391_),
    .B(_08091_),
    .ZN(_08392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17256_ (.A1(_08353_),
    .A2(_08125_),
    .Z(_08393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17257_ (.A1(_08274_),
    .A2(_00390_),
    .ZN(_08394_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17258_ (.A1(_08393_),
    .A2(_08394_),
    .A3(_08260_),
    .ZN(_08395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17259_ (.A1(_08137_),
    .A2(_08116_),
    .A3(_08278_),
    .ZN(_08396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17260_ (.A1(_08395_),
    .A2(_08396_),
    .A3(_08124_),
    .ZN(_08397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17261_ (.A1(_08392_),
    .A2(_08397_),
    .ZN(_08398_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17262_ (.A1(_08387_),
    .A2(_00394_),
    .A3(_08398_),
    .ZN(_08399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17263_ (.A1(_08376_),
    .A2(_08399_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17264_ (.A1(_00390_),
    .A2(net5),
    .ZN(_08400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17265_ (.A1(_07999_),
    .A2(_07986_),
    .A3(_08400_),
    .ZN(_08401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17266_ (.A1(_08331_),
    .A2(_08048_),
    .ZN(_08402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17267_ (.A1(_08065_),
    .A2(net61),
    .ZN(_08403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17268_ (.A1(_08402_),
    .A2(_08403_),
    .A3(_00391_),
    .ZN(_08404_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17269_ (.A1(_08401_),
    .A2(_08404_),
    .A3(_00392_),
    .ZN(_08405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17270_ (.A1(_08024_),
    .A2(_00390_),
    .B(_08080_),
    .ZN(_08406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17271_ (.A1(_08315_),
    .A2(_08058_),
    .ZN(_08407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17272_ (.A1(_08406_),
    .A2(_08407_),
    .B(_07486_),
    .ZN(_08408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17273_ (.A1(_08132_),
    .A2(_08226_),
    .ZN(_08409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17274_ (.A1(_08099_),
    .A2(_08409_),
    .ZN(_08410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17275_ (.A1(_08408_),
    .A2(_08410_),
    .ZN(_08411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17276_ (.A1(_08405_),
    .A2(_08411_),
    .A3(_08076_),
    .ZN(_08412_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17277_ (.I(_07990_),
    .ZN(_08413_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17278_ (.A1(_08301_),
    .A2(_08413_),
    .A3(_07986_),
    .ZN(_08414_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17279_ (.A1(_08194_),
    .A2(_08018_),
    .A3(_08317_),
    .Z(_08415_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17280_ (.A1(_08415_),
    .A2(_08072_),
    .ZN(_08416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17281_ (.A1(_08414_),
    .A2(_08416_),
    .B(_08075_),
    .ZN(_08417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17282_ (.A1(_08079_),
    .A2(_08058_),
    .ZN(_08418_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17283_ (.A1(_08036_),
    .A2(_08418_),
    .A3(_08041_),
    .ZN(_08419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17284_ (.A1(_07996_),
    .A2(_07341_),
    .Z(_08420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17285_ (.A1(_08420_),
    .A2(_08226_),
    .ZN(_08421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17286_ (.A1(_08331_),
    .A2(_08114_),
    .ZN(_08422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17287_ (.A1(_08421_),
    .A2(_00391_),
    .A3(_08422_),
    .ZN(_08423_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17288_ (.A1(_08419_),
    .A2(_08423_),
    .A3(_00392_),
    .ZN(_08424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17289_ (.A1(_08424_),
    .A2(_08417_),
    .ZN(_08425_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17290_ (.A1(_08412_),
    .A2(_08425_),
    .A3(_00393_),
    .ZN(_08426_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17291_ (.I(_08366_),
    .ZN(_08427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17292_ (.A1(_08427_),
    .A2(_08084_),
    .ZN(_08428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17293_ (.A1(_08428_),
    .A2(_08154_),
    .B(_07486_),
    .ZN(_08429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17294_ (.A1(_07978_),
    .A2(net61),
    .Z(_08430_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17295_ (.A1(_08430_),
    .A2(_08009_),
    .B(_08116_),
    .C(_08231_),
    .ZN(_08431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17296_ (.A1(_08429_),
    .A2(_08431_),
    .ZN(_08432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17297_ (.A1(_08107_),
    .A2(net5),
    .ZN(_08433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17298_ (.A1(_08433_),
    .A2(net6),
    .ZN(_08434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17299_ (.A1(_08036_),
    .A2(_08434_),
    .B(_08082_),
    .ZN(_08435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17300_ (.A1(_08023_),
    .A2(_08163_),
    .ZN(_08436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17301_ (.A1(_08436_),
    .A2(_00390_),
    .ZN(_08437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17302_ (.A1(_08037_),
    .A2(_08184_),
    .ZN(_08438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17303_ (.A1(_08438_),
    .A2(_08009_),
    .ZN(_08439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17304_ (.A1(_08437_),
    .A2(_08439_),
    .A3(_08047_),
    .ZN(_08440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17305_ (.A1(_08435_),
    .A2(_08440_),
    .ZN(_08441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17306_ (.A1(_08432_),
    .A2(_08441_),
    .A3(_00394_),
    .ZN(_08442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17307_ (.A1(_08094_),
    .A2(_08088_),
    .ZN(_08443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17308_ (.A1(_08006_),
    .A2(_08058_),
    .A3(_08017_),
    .ZN(_08444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17309_ (.A1(_08443_),
    .A2(_08047_),
    .A3(_08444_),
    .ZN(_08445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17310_ (.A1(_07341_),
    .A2(_07980_),
    .Z(_08446_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17311_ (.A1(_08315_),
    .A2(_08127_),
    .A3(_08446_),
    .Z(_08447_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17312_ (.A1(_08445_),
    .A2(_08447_),
    .A3(_08124_),
    .ZN(_08448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17313_ (.A1(_08055_),
    .A2(_08038_),
    .ZN(_08449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17314_ (.I(_08420_),
    .ZN(_08450_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17315_ (.A1(_08449_),
    .A2(_08450_),
    .A3(_08116_),
    .ZN(_08451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17316_ (.A1(_08205_),
    .A2(_08059_),
    .ZN(_08452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17317_ (.A1(_08451_),
    .A2(_08452_),
    .A3(_08072_),
    .ZN(_08453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17318_ (.A1(_08448_),
    .A2(_08076_),
    .A3(_08453_),
    .ZN(_08454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17319_ (.A1(_08442_),
    .A2(_08454_),
    .A3(_08031_),
    .ZN(_08455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17320_ (.A1(_08426_),
    .A2(_08455_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17321_ (.A1(_08060_),
    .A2(_08006_),
    .ZN(_08456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17322_ (.A1(_08456_),
    .A2(_08150_),
    .A3(_08018_),
    .ZN(_08457_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17323_ (.A1(_08008_),
    .A2(_15559_),
    .Z(_08458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17324_ (.A1(_08402_),
    .A2(_07985_),
    .A3(_08458_),
    .ZN(_08459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17325_ (.A1(_08457_),
    .A2(_08459_),
    .ZN(_08460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17326_ (.A1(_08460_),
    .A2(_08072_),
    .ZN(_08461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17327_ (.A1(_08357_),
    .A2(_08141_),
    .ZN(_08462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17328_ (.A1(_08462_),
    .A2(_08260_),
    .ZN(_08463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17329_ (.A1(_08237_),
    .A2(_08027_),
    .Z(_08464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17330_ (.A1(_08463_),
    .A2(_08464_),
    .ZN(_08465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17331_ (.A1(_08461_),
    .A2(_08091_),
    .A3(_08465_),
    .ZN(_08466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17332_ (.A1(_08339_),
    .A2(_08107_),
    .ZN(_08467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17333_ (.A1(_08301_),
    .A2(_08467_),
    .ZN(_08468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17334_ (.A1(_08468_),
    .A2(_08116_),
    .ZN(_08469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17335_ (.A1(_08057_),
    .A2(_08203_),
    .ZN(_08470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17336_ (.A1(_08470_),
    .A2(_08127_),
    .ZN(_08471_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17337_ (.A1(_08469_),
    .A2(_08124_),
    .A3(_08471_),
    .ZN(_08472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17338_ (.A1(_07998_),
    .A2(_08063_),
    .ZN(_08473_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17339_ (.A1(_08473_),
    .A2(_08149_),
    .Z(_08474_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17340_ (.A1(_08048_),
    .A2(_07989_),
    .Z(_08475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17341_ (.A1(_08475_),
    .A2(_08317_),
    .ZN(_08476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17342_ (.A1(_08474_),
    .A2(_08476_),
    .A3(_08080_),
    .ZN(_08477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17343_ (.A1(_08473_),
    .A2(_08166_),
    .ZN(_08478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17344_ (.A1(_08121_),
    .A2(_07513_),
    .Z(_08479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17345_ (.A1(_08478_),
    .A2(_08479_),
    .B(_08027_),
    .ZN(_08480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17346_ (.A1(_08477_),
    .A2(_08480_),
    .B(_08091_),
    .ZN(_08481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17347_ (.A1(_08472_),
    .A2(_08481_),
    .ZN(_08482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17348_ (.A1(_08466_),
    .A2(_08482_),
    .ZN(_08483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17349_ (.A1(_08483_),
    .A2(_08076_),
    .ZN(_08484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17350_ (.A1(_08217_),
    .A2(_08243_),
    .ZN(_08485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17351_ (.A1(_00390_),
    .A2(_08485_),
    .ZN(_08486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17352_ (.A1(_08372_),
    .A2(_08486_),
    .B(_08082_),
    .ZN(_08487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17353_ (.A1(_08353_),
    .A2(_08021_),
    .ZN(_08488_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17354_ (.A1(_08488_),
    .A2(_08069_),
    .A3(_08201_),
    .ZN(_08489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17355_ (.A1(_08489_),
    .A2(_08487_),
    .B(_08091_),
    .ZN(_08490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17356_ (.A1(_07997_),
    .A2(_08086_),
    .ZN(_08491_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17357_ (.A1(_08301_),
    .A2(_08491_),
    .A3(_08047_),
    .ZN(_08492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17358_ (.A1(_08040_),
    .A2(_08021_),
    .B(_08018_),
    .ZN(_08493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17359_ (.A1(_08331_),
    .A2(_08044_),
    .ZN(_08494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17360_ (.A1(_08197_),
    .A2(_08162_),
    .ZN(_08495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17361_ (.A1(_08493_),
    .A2(_08494_),
    .A3(_08495_),
    .ZN(_08496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17362_ (.A1(_08492_),
    .A2(_08028_),
    .A3(_08496_),
    .ZN(_08497_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17363_ (.A1(_08497_),
    .A2(_08490_),
    .B(_08075_),
    .ZN(_08498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17364_ (.A1(_08005_),
    .A2(_08114_),
    .ZN(_08499_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17365_ (.A1(_08009_),
    .A2(_08499_),
    .B(_08025_),
    .C(_08260_),
    .ZN(_08500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17366_ (.A1(_08121_),
    .A2(_08021_),
    .A3(_08114_),
    .ZN(_08501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17367_ (.A1(_08491_),
    .A2(_08069_),
    .A3(_08501_),
    .ZN(_08502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17368_ (.A1(_08500_),
    .A2(_08028_),
    .A3(_08502_),
    .ZN(_08503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17369_ (.A1(_08427_),
    .A2(_08006_),
    .ZN(_08504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17370_ (.A1(_08065_),
    .A2(_08048_),
    .ZN(_08505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17371_ (.A1(_08504_),
    .A2(_07986_),
    .A3(_08505_),
    .ZN(_08506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17372_ (.A1(_07990_),
    .A2(_08050_),
    .ZN(_08507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17373_ (.A1(_08507_),
    .A2(_08047_),
    .A3(_08269_),
    .ZN(_08508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17374_ (.A1(_08506_),
    .A2(_08508_),
    .A3(_08072_),
    .ZN(_08509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17375_ (.A1(_08503_),
    .A2(_08509_),
    .A3(_08031_),
    .ZN(_08510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17376_ (.A1(_08510_),
    .A2(_08498_),
    .ZN(_08511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17377_ (.A1(_08511_),
    .A2(_08484_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17378_ (.A1(_08287_),
    .A2(_08114_),
    .ZN(_08512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17379_ (.A1(_08336_),
    .A2(_08512_),
    .A3(_08495_),
    .ZN(_08513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17380_ (.A1(_08166_),
    .A2(_07985_),
    .Z(_08514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17381_ (.A1(_08514_),
    .A2(_08357_),
    .B(_08082_),
    .ZN(_08515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17382_ (.A1(_08513_),
    .A2(_08515_),
    .B(_08091_),
    .ZN(_08516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17383_ (.A1(_08288_),
    .A2(_00391_),
    .A3(_08209_),
    .ZN(_08517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17384_ (.A1(_08255_),
    .A2(_08494_),
    .A3(_07986_),
    .ZN(_08518_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17385_ (.A1(_08517_),
    .A2(_08518_),
    .A3(_08028_),
    .ZN(_08519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17386_ (.A1(_08516_),
    .A2(_08519_),
    .ZN(_08520_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17387_ (.A1(_08006_),
    .A2(_07993_),
    .A3(_08107_),
    .ZN(_08521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17388_ (.A1(_08521_),
    .A2(_08257_),
    .ZN(_08522_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17389_ (.A1(_08522_),
    .A2(_08260_),
    .ZN(_08523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17390_ (.A1(_08163_),
    .A2(_08125_),
    .ZN(_08524_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17391_ (.A1(_08413_),
    .A2(_08524_),
    .A3(_08080_),
    .ZN(_08525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17392_ (.A1(_08523_),
    .A2(_08525_),
    .ZN(_08526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17393_ (.A1(_08526_),
    .A2(_08028_),
    .ZN(_08527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17394_ (.A1(_08420_),
    .A2(_08138_),
    .ZN(_08528_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17395_ (.A1(_08433_),
    .A2(_08018_),
    .Z(_08529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17396_ (.A1(_08528_),
    .A2(_08529_),
    .B(_08082_),
    .ZN(_08530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17397_ (.A1(_08475_),
    .A2(_07993_),
    .ZN(_08531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17398_ (.A1(_08531_),
    .A2(_07986_),
    .A3(_08278_),
    .ZN(_08532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17399_ (.A1(_08530_),
    .A2(_08532_),
    .ZN(_08533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17400_ (.A1(_08527_),
    .A2(_08533_),
    .A3(_08031_),
    .ZN(_08534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17401_ (.A1(_08520_),
    .A2(_08534_),
    .A3(_08076_),
    .ZN(_08535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17402_ (.A1(_08085_),
    .A2(_07993_),
    .ZN(_08536_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17403_ (.A1(_08536_),
    .A2(_00391_),
    .A3(_08307_),
    .ZN(_08537_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17404_ (.A1(_08006_),
    .A2(_08088_),
    .A3(_08021_),
    .ZN(_08538_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17405_ (.A1(_08119_),
    .A2(_07993_),
    .A3(_08049_),
    .ZN(_08539_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17406_ (.A1(_08538_),
    .A2(_08539_),
    .A3(_08069_),
    .ZN(_08540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17407_ (.A1(_08537_),
    .A2(_08540_),
    .A3(_00392_),
    .ZN(_08541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17408_ (.A1(_08009_),
    .A2(_15546_),
    .ZN(_08542_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17409_ (.A1(_08488_),
    .A2(_08047_),
    .A3(_08542_),
    .ZN(_08543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17410_ (.A1(_08033_),
    .A2(_08021_),
    .B(_08018_),
    .ZN(_08544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17411_ (.A1(_08244_),
    .A2(_08017_),
    .ZN(_08545_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17412_ (.A1(_08544_),
    .A2(_08545_),
    .A3(_08015_),
    .ZN(_08546_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17413_ (.A1(_08543_),
    .A2(_08546_),
    .A3(_08124_),
    .ZN(_08547_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17414_ (.A1(_08541_),
    .A2(_08547_),
    .A3(_00393_),
    .ZN(_08548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17415_ (.A1(_08006_),
    .A2(_08011_),
    .A3(_08125_),
    .ZN(_08549_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17416_ (.A1(_00391_),
    .A2(_08150_),
    .A3(_08549_),
    .A4(_08259_),
    .ZN(_08550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17417_ (.A1(_08001_),
    .A2(_15569_),
    .ZN(_08551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17418_ (.A1(_08551_),
    .A2(_07985_),
    .ZN(_08552_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17419_ (.A1(_08552_),
    .A2(_08097_),
    .ZN(_08553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17420_ (.A1(_08012_),
    .A2(_08049_),
    .ZN(_08554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17421_ (.A1(_08553_),
    .A2(_08554_),
    .B(_07486_),
    .ZN(_08555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17422_ (.A1(_08550_),
    .A2(_08555_),
    .ZN(_08556_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17423_ (.A1(_15539_),
    .A2(_08107_),
    .B(_08035_),
    .ZN(_08557_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17424_ (.I(_08557_),
    .ZN(_08558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17425_ (.A1(_08558_),
    .A2(_08545_),
    .B(_08082_),
    .ZN(_08559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17426_ (.A1(_08139_),
    .A2(_08108_),
    .A3(_08034_),
    .ZN(_08560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17427_ (.A1(_08559_),
    .A2(_08560_),
    .ZN(_08561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17428_ (.A1(_08556_),
    .A2(_08561_),
    .A3(_08031_),
    .ZN(_08562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17429_ (.A1(_08548_),
    .A2(_08562_),
    .A3(_00394_),
    .ZN(_08563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17430_ (.A1(_08535_),
    .A2(_08563_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17431_ (.A1(_07404_),
    .A2(_07609_),
    .B(_07612_),
    .ZN(_15571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17432_ (.A1(_07286_),
    .A2(_07618_),
    .B(_07620_),
    .ZN(_08564_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17433_ (.I(_08564_),
    .Z(_15591_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17434_ (.A1(_07467_),
    .A2(_07601_),
    .B(_07604_),
    .ZN(_15572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17435_ (.A1(_15582_),
    .A2(_08564_),
    .ZN(_08565_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17436_ (.I(_08565_),
    .ZN(_08566_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17437_ (.I(_07629_),
    .Z(_08567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17438_ (.A1(_08566_),
    .A2(_08567_),
    .ZN(_08568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17439_ (.A1(_07622_),
    .A2(_15589_),
    .Z(_08569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17440_ (.A1(_08569_),
    .A2(_08567_),
    .ZN(_08570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17441_ (.A1(_08568_),
    .A2(_08570_),
    .ZN(_08571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17442_ (.I(_08571_),
    .ZN(_08572_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17443_ (.I(_07638_),
    .Z(_08573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17444_ (.I(_08573_),
    .Z(_08574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17445_ (.A1(_08564_),
    .A2(_15572_),
    .ZN(_08575_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17446_ (.I(_08575_),
    .ZN(_08576_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17447_ (.I(_15573_),
    .ZN(_08577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17448_ (.A1(_07622_),
    .A2(_08577_),
    .ZN(_08578_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _17449_ (.I(_08578_),
    .ZN(_08579_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17450_ (.I(_07630_),
    .Z(_08580_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17451_ (.A1(_08576_),
    .A2(_08579_),
    .B(_08580_),
    .ZN(_08581_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17452_ (.A1(_08572_),
    .A2(_08574_),
    .A3(_08581_),
    .ZN(_08582_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17453_ (.I(_08564_),
    .Z(_08583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17454_ (.A1(_08583_),
    .A2(_15578_),
    .ZN(_08584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17455_ (.A1(_08584_),
    .A2(_07629_),
    .ZN(_08585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17456_ (.I(_08585_),
    .ZN(_08586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17457_ (.A1(net78),
    .A2(_07622_),
    .ZN(_08587_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17458_ (.I(_08587_),
    .Z(_08588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17459_ (.A1(_08586_),
    .A2(_08588_),
    .ZN(_08589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17460_ (.A1(_15577_),
    .A2(_08583_),
    .ZN(_08590_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17461_ (.I(_15575_),
    .ZN(_08591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17462_ (.A1(_08591_),
    .A2(_15596_),
    .ZN(_08592_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17463_ (.A1(_08590_),
    .A2(_08592_),
    .A3(_00385_),
    .ZN(_08593_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17464_ (.A1(_08589_),
    .A2(_08593_),
    .A3(_00386_),
    .ZN(_08594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17465_ (.I(_07647_),
    .ZN(_08595_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17466_ (.I(_08595_),
    .Z(_08596_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17467_ (.I(_08596_),
    .Z(_08597_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17468_ (.A1(_08582_),
    .A2(_08594_),
    .A3(_08597_),
    .ZN(_08598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17469_ (.A1(_08564_),
    .A2(_08591_),
    .ZN(_08599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17470_ (.A1(_08599_),
    .A2(_07630_),
    .ZN(_08600_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17471_ (.I(_08600_),
    .ZN(_08601_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17472_ (.I(_15574_),
    .ZN(_08602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17473_ (.A1(_08602_),
    .A2(_15596_),
    .ZN(_08603_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17474_ (.I(_08603_),
    .Z(_08604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17475_ (.A1(_08601_),
    .A2(net79),
    .ZN(_08605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17476_ (.A1(_15577_),
    .A2(_15596_),
    .ZN(_08606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17477_ (.A1(_08586_),
    .A2(_08606_),
    .ZN(_08607_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17478_ (.A1(_08605_),
    .A2(_08607_),
    .A3(_00386_),
    .ZN(_08608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17479_ (.A1(_08584_),
    .A2(_07631_),
    .ZN(_08609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17480_ (.I(_08609_),
    .ZN(_08610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17481_ (.I(_15580_),
    .ZN(_08611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17482_ (.A1(_07622_),
    .A2(_08611_),
    .ZN(_08612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17483_ (.A1(_08610_),
    .A2(_08612_),
    .ZN(_08613_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17484_ (.I(_08573_),
    .Z(_08614_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17485_ (.I(_07629_),
    .Z(_08615_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17486_ (.A1(_08590_),
    .A2(_08615_),
    .Z(_08616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17487_ (.I(_08616_),
    .ZN(_08617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17488_ (.A1(_08613_),
    .A2(_08614_),
    .A3(_08617_),
    .ZN(_08618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17489_ (.A1(_08608_),
    .A2(_08618_),
    .A3(_00387_),
    .ZN(_08619_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17490_ (.A1(_08598_),
    .A2(_08619_),
    .A3(_00388_),
    .ZN(_08620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17491_ (.A1(_07622_),
    .A2(_15572_),
    .ZN(_08621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17492_ (.A1(_08621_),
    .A2(_08615_),
    .Z(_08622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17493_ (.A1(_15577_),
    .A2(net78),
    .ZN(_08623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17494_ (.A1(_08622_),
    .A2(_08623_),
    .ZN(_08624_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17495_ (.I(_08621_),
    .ZN(_08625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17496_ (.A1(net77),
    .A2(net30),
    .ZN(_08626_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17497_ (.I(_07630_),
    .Z(_08627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17498_ (.A1(_08625_),
    .A2(_08626_),
    .B(_08627_),
    .ZN(_08628_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17499_ (.A1(_08624_),
    .A2(_08628_),
    .A3(_00386_),
    .ZN(_08629_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17500_ (.I(_15583_),
    .ZN(_08630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17501_ (.A1(_15596_),
    .A2(_08630_),
    .ZN(_08631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17502_ (.I(_08631_),
    .ZN(_08632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17503_ (.I(_15587_),
    .ZN(_08633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17504_ (.A1(_15591_),
    .A2(_08633_),
    .ZN(_08634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17505_ (.I(_08634_),
    .ZN(_08635_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17506_ (.A1(_08632_),
    .A2(_08635_),
    .B(_00385_),
    .ZN(_08636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17507_ (.A1(_08583_),
    .A2(_15573_),
    .ZN(_08637_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17508_ (.I(_08567_),
    .Z(_08638_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17509_ (.A1(net79),
    .A2(_08637_),
    .A3(_08638_),
    .ZN(_08639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17510_ (.A1(_08639_),
    .A2(_08614_),
    .A3(_08636_),
    .ZN(_08640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17511_ (.A1(_08629_),
    .A2(_08640_),
    .A3(_00387_),
    .ZN(_08641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17512_ (.I(_07654_),
    .ZN(_08642_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17513_ (.I(_08642_),
    .Z(_08643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17514_ (.A1(_08583_),
    .A2(_08630_),
    .ZN(_08644_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17515_ (.I(_08644_),
    .ZN(_08645_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17516_ (.A1(_08583_),
    .A2(_15587_),
    .ZN(_08646_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17517_ (.A1(_08645_),
    .A2(_08646_),
    .B(_08638_),
    .ZN(_08647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17518_ (.A1(net84),
    .A2(_15587_),
    .ZN(_08648_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17519_ (.I(_07631_),
    .Z(_08649_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17520_ (.A1(_08604_),
    .A2(_08648_),
    .A3(_08649_),
    .ZN(_08650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17521_ (.I(_08573_),
    .Z(_08651_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17522_ (.A1(_08647_),
    .A2(_08650_),
    .A3(_08651_),
    .ZN(_08652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17523_ (.A1(_15591_),
    .A2(net30),
    .ZN(_08653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17524_ (.A1(_07622_),
    .A2(_15574_),
    .ZN(_08654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17525_ (.A1(_08653_),
    .A2(_08654_),
    .ZN(_08655_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17526_ (.I(_07629_),
    .Z(_08656_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17527_ (.I(_08656_),
    .Z(_08657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17528_ (.A1(_08655_),
    .A2(_08657_),
    .ZN(_08658_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17529_ (.I(_07640_),
    .Z(_08659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17530_ (.A1(_08602_),
    .A2(_08583_),
    .ZN(_08660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17531_ (.I(_08660_),
    .ZN(_08661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17532_ (.A1(_07631_),
    .A2(_08661_),
    .ZN(_08662_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17533_ (.A1(_08658_),
    .A2(_08659_),
    .A3(_08662_),
    .ZN(_08663_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17534_ (.I(_08595_),
    .Z(_08664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17535_ (.A1(_08652_),
    .A2(_08663_),
    .A3(_08664_),
    .ZN(_08665_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17536_ (.A1(_08665_),
    .A2(_08643_),
    .A3(_08641_),
    .ZN(_08666_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17537_ (.I(_07660_),
    .ZN(_08667_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17538_ (.I(_08667_),
    .Z(_08668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17539_ (.A1(_08620_),
    .A2(_08666_),
    .A3(_08668_),
    .ZN(_08669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17540_ (.A1(_08569_),
    .A2(_07630_),
    .ZN(_08670_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17541_ (.I(_07629_),
    .Z(_08671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17542_ (.A1(_08645_),
    .A2(_08671_),
    .ZN(_08672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17543_ (.A1(_08670_),
    .A2(_08672_),
    .Z(_08673_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17544_ (.I(_15578_),
    .ZN(_08674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17545_ (.A1(_15596_),
    .A2(_08674_),
    .Z(_08675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17546_ (.A1(_08675_),
    .A2(_08656_),
    .B(_07638_),
    .ZN(_08676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17547_ (.A1(_08673_),
    .A2(_08676_),
    .B(_07654_),
    .ZN(_08677_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17548_ (.I(_15585_),
    .ZN(_08678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17549_ (.A1(_08678_),
    .A2(_08564_),
    .ZN(_08679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17550_ (.A1(_08679_),
    .A2(_07630_),
    .ZN(_08680_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17551_ (.I(_08680_),
    .ZN(_08681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17552_ (.A1(_15596_),
    .A2(_15578_),
    .ZN(_08682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17553_ (.A1(_08681_),
    .A2(_08682_),
    .ZN(_08683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17554_ (.A1(_08683_),
    .A2(_08614_),
    .A3(_08570_),
    .ZN(_08684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17555_ (.A1(_08677_),
    .A2(_08684_),
    .B(_08664_),
    .ZN(_08685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17556_ (.A1(_07622_),
    .A2(_15571_),
    .ZN(_08686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17557_ (.A1(_08686_),
    .A2(_08615_),
    .Z(_08687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17558_ (.A1(_15574_),
    .A2(_08564_),
    .ZN(_08688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17559_ (.A1(_08687_),
    .A2(_08688_),
    .ZN(_08689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17560_ (.A1(net84),
    .A2(_15583_),
    .ZN(_08690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17561_ (.A1(_08606_),
    .A2(_08690_),
    .A3(_08649_),
    .ZN(_08691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17562_ (.A1(_08689_),
    .A2(_08691_),
    .B(_08659_),
    .ZN(_08692_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17563_ (.I(_08615_),
    .Z(_08693_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17564_ (.A1(_08569_),
    .A2(_08635_),
    .B(_08693_),
    .ZN(_08694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17565_ (.A1(_08612_),
    .A2(_07631_),
    .ZN(_08695_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17566_ (.I(_08573_),
    .Z(_08696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17567_ (.A1(_08694_),
    .A2(_08695_),
    .B(_08696_),
    .ZN(_08697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17568_ (.I(_07654_),
    .Z(_08698_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17569_ (.A1(_08692_),
    .A2(_08697_),
    .B(_08698_),
    .ZN(_08699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17570_ (.A1(_08685_),
    .A2(_08699_),
    .ZN(_08700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17571_ (.A1(_08583_),
    .A2(_15580_),
    .ZN(_08701_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17572_ (.I(_08701_),
    .ZN(_08702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17573_ (.A1(_08702_),
    .A2(_08657_),
    .ZN(_08703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17574_ (.A1(_08581_),
    .A2(_08614_),
    .A3(_08703_),
    .ZN(_08704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17575_ (.A1(_15596_),
    .A2(_15585_),
    .ZN(_08705_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17576_ (.I(_08705_),
    .ZN(_08706_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17577_ (.A1(_08706_),
    .A2(_08702_),
    .B(_08693_),
    .ZN(_08707_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17578_ (.I(_07640_),
    .Z(_08708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17579_ (.A1(_07630_),
    .A2(_08603_),
    .ZN(_08709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17580_ (.A1(_08707_),
    .A2(_08708_),
    .A3(_08709_),
    .ZN(_08710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17581_ (.A1(_08704_),
    .A2(_08710_),
    .A3(_08698_),
    .ZN(_08711_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17582_ (.A1(_08576_),
    .A2(_08646_),
    .B(_08580_),
    .ZN(_08712_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17583_ (.A1(_08575_),
    .A2(_08682_),
    .A3(_08638_),
    .ZN(_08713_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17584_ (.A1(_08712_),
    .A2(_08713_),
    .A3(_08651_),
    .ZN(_08714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17585_ (.A1(_08627_),
    .A2(_15599_),
    .ZN(_08715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17586_ (.A1(_08715_),
    .A2(_07640_),
    .ZN(_08716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17587_ (.I(_08716_),
    .ZN(_08717_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17588_ (.I(_08688_),
    .ZN(_08718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17589_ (.A1(_08718_),
    .A2(_08638_),
    .ZN(_08719_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17590_ (.A1(_08717_),
    .A2(_08719_),
    .B(_07654_),
    .ZN(_08720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17591_ (.A1(_08714_),
    .A2(_08720_),
    .ZN(_08721_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17592_ (.A1(_08711_),
    .A2(_08597_),
    .A3(_08721_),
    .ZN(_08722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17593_ (.A1(_08700_),
    .A2(_08722_),
    .A3(_00389_),
    .ZN(_08723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17594_ (.A1(_08669_),
    .A2(_08723_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17595_ (.A1(_08567_),
    .A2(_15592_),
    .B(_07639_),
    .ZN(_08724_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17596_ (.I(_08724_),
    .ZN(_08725_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17597_ (.A1(_08611_),
    .A2(_07619_),
    .A3(_07621_),
    .ZN(_08726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17598_ (.A1(_08687_),
    .A2(_08726_),
    .ZN(_08727_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _17599_ (.I(_07647_),
    .Z(_08728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17600_ (.A1(_08725_),
    .A2(_08727_),
    .B(_08728_),
    .ZN(_08729_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17601_ (.A1(_08592_),
    .A2(_08660_),
    .A3(_08580_),
    .ZN(_08730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17602_ (.A1(_08682_),
    .A2(_08726_),
    .A3(_08638_),
    .ZN(_08731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17603_ (.A1(_08730_),
    .A2(_08731_),
    .A3(_08574_),
    .ZN(_08732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17604_ (.A1(_08729_),
    .A2(_08732_),
    .B(_00388_),
    .ZN(_08733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17605_ (.A1(_08612_),
    .A2(_08615_),
    .Z(_08734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17606_ (.A1(_08734_),
    .A2(_08575_),
    .ZN(_08735_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17607_ (.I(_08709_),
    .ZN(_08736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17608_ (.A1(_08736_),
    .A2(_08590_),
    .ZN(_08737_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17609_ (.A1(_08735_),
    .A2(_08737_),
    .A3(_00386_),
    .ZN(_08738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17610_ (.A1(_08687_),
    .A2(_08623_),
    .ZN(_08739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17611_ (.A1(_07631_),
    .A2(net84),
    .Z(_08740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17612_ (.A1(_08740_),
    .A2(_08674_),
    .ZN(_08741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17613_ (.A1(_08739_),
    .A2(_08574_),
    .A3(_08741_),
    .ZN(_08742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17614_ (.A1(_08738_),
    .A2(_08742_),
    .A3(_00387_),
    .ZN(_08743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17615_ (.A1(_08743_),
    .A2(_08733_),
    .ZN(_08744_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17616_ (.A1(_15577_),
    .A2(net30),
    .B(_08590_),
    .C(_08649_),
    .ZN(_08745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17617_ (.A1(_08606_),
    .A2(_08567_),
    .Z(_08746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17618_ (.A1(_08746_),
    .A2(_08688_),
    .ZN(_08747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17619_ (.A1(_08745_),
    .A2(_08574_),
    .A3(_08747_),
    .ZN(_08748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17620_ (.A1(_08576_),
    .A2(_08567_),
    .B(_07638_),
    .ZN(_08749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17621_ (.A1(_08726_),
    .A2(_07630_),
    .ZN(_08750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17622_ (.I(_08750_),
    .ZN(_08751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17623_ (.A1(_08751_),
    .A2(_08654_),
    .ZN(_08752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17624_ (.A1(_08646_),
    .A2(_08567_),
    .ZN(_08753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17625_ (.A1(_08749_),
    .A2(_08752_),
    .A3(_08753_),
    .ZN(_08754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17626_ (.A1(_08748_),
    .A2(_08754_),
    .A3(_08597_),
    .ZN(_08755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17627_ (.A1(_15596_),
    .A2(_15580_),
    .Z(_08756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17628_ (.I(_07639_),
    .Z(_08757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17629_ (.A1(_08756_),
    .A2(_08657_),
    .B(_08757_),
    .ZN(_08758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17630_ (.A1(_08637_),
    .A2(_07630_),
    .ZN(_08759_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17631_ (.I(_08759_),
    .ZN(_08760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17632_ (.A1(_08760_),
    .A2(_08654_),
    .ZN(_08761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17633_ (.A1(_08758_),
    .A2(_08761_),
    .B(_08596_),
    .ZN(_08762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17634_ (.A1(_08601_),
    .A2(_08588_),
    .ZN(_08763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17635_ (.A1(_08567_),
    .A2(_08579_),
    .ZN(_08764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17636_ (.A1(_08763_),
    .A2(_08708_),
    .A3(_08764_),
    .ZN(_08765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17637_ (.A1(_08762_),
    .A2(_08765_),
    .B(_08642_),
    .ZN(_08766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17638_ (.A1(_08755_),
    .A2(_08766_),
    .ZN(_08767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17639_ (.A1(_08744_),
    .A2(_08767_),
    .A3(_00389_),
    .ZN(_08768_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17640_ (.A1(_08695_),
    .A2(_08566_),
    .Z(_08769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17641_ (.A1(_08622_),
    .A2(_08653_),
    .ZN(_08770_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17642_ (.A1(_08769_),
    .A2(_08770_),
    .A3(_08664_),
    .ZN(_08771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17643_ (.A1(_08746_),
    .A2(_08648_),
    .ZN(_08772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17644_ (.A1(_08579_),
    .A2(_08649_),
    .B(_08595_),
    .ZN(_08773_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17645_ (.A1(_08772_),
    .A2(_08773_),
    .A3(_08741_),
    .ZN(_08774_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17646_ (.A1(_08771_),
    .A2(_08774_),
    .A3(_00386_),
    .ZN(_08775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17647_ (.A1(_08578_),
    .A2(_08644_),
    .B(_08627_),
    .ZN(_08776_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17648_ (.I(_08776_),
    .ZN(_08777_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17649_ (.A1(_07647_),
    .A2(_15601_),
    .A3(_08671_),
    .Z(_08778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17650_ (.A1(_08777_),
    .A2(_08778_),
    .ZN(_08779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17651_ (.A1(_08779_),
    .A2(_08574_),
    .B(_08698_),
    .ZN(_08780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17652_ (.A1(_08775_),
    .A2(_08780_),
    .B(_00389_),
    .ZN(_08781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17653_ (.A1(_08646_),
    .A2(_08627_),
    .ZN(_08782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17654_ (.A1(_08615_),
    .A2(_08688_),
    .ZN(_08783_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _17655_ (.I(_08783_),
    .ZN(_08784_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17656_ (.A1(_08570_),
    .A2(_08749_),
    .A3(_08782_),
    .A4(_08784_),
    .ZN(_08785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17657_ (.A1(_08622_),
    .A2(_08648_),
    .ZN(_08786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17658_ (.A1(_08769_),
    .A2(_08786_),
    .A3(_08574_),
    .ZN(_08787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17659_ (.A1(_08785_),
    .A2(_00387_),
    .A3(_08787_),
    .ZN(_08788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17660_ (.A1(_08764_),
    .A2(_08573_),
    .ZN(_08789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17661_ (.I(_08789_),
    .ZN(_08790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17662_ (.A1(_08709_),
    .A2(_08575_),
    .Z(_08791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17663_ (.A1(_08790_),
    .A2(_08791_),
    .B(_08728_),
    .ZN(_08792_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17664_ (.I(_15589_),
    .ZN(_08793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17665_ (.A1(_08583_),
    .A2(_08793_),
    .ZN(_08794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17666_ (.A1(_08794_),
    .A2(_08615_),
    .ZN(_08795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17667_ (.I(_08795_),
    .ZN(_08796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17668_ (.A1(_08796_),
    .A2(_08592_),
    .ZN(_08797_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17669_ (.A1(_08761_),
    .A2(_08797_),
    .A3(_08708_),
    .ZN(_08798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17670_ (.A1(_08792_),
    .A2(_08798_),
    .B(_08643_),
    .ZN(_08799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17671_ (.A1(_08799_),
    .A2(_08788_),
    .ZN(_08800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17672_ (.A1(_08781_),
    .A2(_08800_),
    .ZN(_08801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17673_ (.A1(_08768_),
    .A2(_08801_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17674_ (.A1(net84),
    .A2(_15575_),
    .ZN(_08802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17675_ (.A1(_08622_),
    .A2(_08802_),
    .ZN(_08803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17676_ (.A1(_08565_),
    .A2(_08705_),
    .A3(_08580_),
    .ZN(_08804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17677_ (.A1(_08803_),
    .A2(_08804_),
    .A3(_08659_),
    .ZN(_08805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17678_ (.A1(_08606_),
    .A2(_08679_),
    .A3(_08656_),
    .ZN(_08806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17679_ (.A1(_08603_),
    .A2(_08688_),
    .A3(_08627_),
    .ZN(_08807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17680_ (.A1(_08806_),
    .A2(_08807_),
    .ZN(_08808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17681_ (.A1(_08808_),
    .A2(_08696_),
    .ZN(_08809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17682_ (.A1(_08805_),
    .A2(_08809_),
    .ZN(_08810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17683_ (.A1(_08810_),
    .A2(_00387_),
    .ZN(_08811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17684_ (.A1(_08751_),
    .A2(_08588_),
    .ZN(_08812_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17685_ (.A1(_08707_),
    .A2(_08812_),
    .A3(_08574_),
    .ZN(_08813_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17686_ (.I(_08802_),
    .ZN(_08814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17687_ (.A1(_08814_),
    .A2(_08693_),
    .B(_08573_),
    .ZN(_08815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17688_ (.A1(_08751_),
    .A2(_08606_),
    .ZN(_08816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17689_ (.A1(_08706_),
    .A2(_08656_),
    .ZN(_08817_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17690_ (.A1(_08815_),
    .A2(_08816_),
    .A3(_08817_),
    .ZN(_08818_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17691_ (.A1(_08813_),
    .A2(_08818_),
    .A3(_08664_),
    .ZN(_08819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17692_ (.A1(_08811_),
    .A2(_08819_),
    .A3(_00388_),
    .ZN(_08820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17693_ (.I(_08689_),
    .ZN(_08821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17694_ (.A1(_08701_),
    .A2(_07631_),
    .ZN(_08822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17695_ (.A1(_08822_),
    .A2(_08675_),
    .B(_07638_),
    .ZN(_08823_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17696_ (.A1(_08821_),
    .A2(_08823_),
    .ZN(_08824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17697_ (.A1(_08686_),
    .A2(_08584_),
    .A3(_08580_),
    .ZN(_08825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17698_ (.A1(_08612_),
    .A2(_08599_),
    .A3(_08693_),
    .ZN(_08826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17699_ (.A1(_08825_),
    .A2(_08826_),
    .B(_08696_),
    .ZN(_08827_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17700_ (.A1(_08824_),
    .A2(_08827_),
    .B(_08664_),
    .ZN(_08828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17701_ (.A1(_08585_),
    .A2(_08573_),
    .Z(_08829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17702_ (.A1(_08760_),
    .A2(_08592_),
    .ZN(_08830_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17703_ (.A1(_08829_),
    .A2(_08830_),
    .B(_08596_),
    .ZN(_08831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17704_ (.A1(_15591_),
    .A2(_15589_),
    .ZN(_08832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17705_ (.I(_08832_),
    .ZN(_08833_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17706_ (.A1(_08625_),
    .A2(_08833_),
    .B(_00385_),
    .ZN(_08834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17707_ (.A1(_08653_),
    .A2(net79),
    .A3(_08638_),
    .ZN(_08835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17708_ (.A1(_08834_),
    .A2(_08708_),
    .A3(_08835_),
    .ZN(_08836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17709_ (.A1(_08831_),
    .A2(_08836_),
    .ZN(_08837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17710_ (.A1(_08828_),
    .A2(_08643_),
    .A3(_08837_),
    .ZN(_08838_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17711_ (.A1(_08820_),
    .A2(_08838_),
    .A3(_08668_),
    .ZN(_08839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17712_ (.A1(_08623_),
    .A2(_08686_),
    .A3(_08580_),
    .ZN(_08840_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17713_ (.A1(_15601_),
    .A2(_00385_),
    .B(_08840_),
    .C(_08651_),
    .ZN(_08841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17714_ (.A1(_08784_),
    .A2(_07640_),
    .Z(_08842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17715_ (.A1(_08632_),
    .A2(_00385_),
    .ZN(_08843_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17716_ (.A1(_08588_),
    .A2(_08648_),
    .A3(_08638_),
    .ZN(_08844_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17717_ (.A1(_08842_),
    .A2(_08843_),
    .A3(_08844_),
    .ZN(_08845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17718_ (.A1(_08841_),
    .A2(_08597_),
    .A3(_08845_),
    .ZN(_08846_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17719_ (.A1(_08625_),
    .A2(_15594_),
    .B(_08649_),
    .ZN(_08847_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17720_ (.A1(_08689_),
    .A2(_08847_),
    .A3(_00386_),
    .ZN(_08848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17721_ (.A1(_08682_),
    .A2(_07630_),
    .ZN(_08849_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17722_ (.A1(_08567_),
    .A2(_15599_),
    .Z(_08850_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17723_ (.I(_08850_),
    .ZN(_08851_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17724_ (.A1(_08849_),
    .A2(_08661_),
    .B(_08851_),
    .C(_08696_),
    .ZN(_08852_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17725_ (.A1(_08848_),
    .A2(_00387_),
    .A3(_08852_),
    .ZN(_08853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17726_ (.A1(_08846_),
    .A2(_08853_),
    .A3(_00388_),
    .ZN(_08854_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17727_ (.A1(_08615_),
    .A2(_15597_),
    .Z(_08855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17728_ (.A1(_08829_),
    .A2(_08855_),
    .B(_07647_),
    .ZN(_08856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17729_ (.A1(_08657_),
    .A2(_15594_),
    .ZN(_08857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17730_ (.A1(_08825_),
    .A2(_08708_),
    .A3(_08857_),
    .ZN(_08858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17731_ (.A1(_08856_),
    .A2(_08858_),
    .B(_08698_),
    .ZN(_08859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17732_ (.A1(_08760_),
    .A2(_08621_),
    .ZN(_08860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17733_ (.A1(_08777_),
    .A2(_08860_),
    .A3(_08708_),
    .ZN(_08861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17734_ (.A1(_08736_),
    .A2(_08726_),
    .ZN(_08862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17735_ (.A1(_08862_),
    .A2(_08651_),
    .A3(_08753_),
    .ZN(_08863_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17736_ (.A1(_08861_),
    .A2(_08863_),
    .A3(_08728_),
    .ZN(_08864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17737_ (.A1(_08859_),
    .A2(_08864_),
    .B(_08668_),
    .ZN(_08865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17738_ (.A1(_08854_),
    .A2(_08865_),
    .ZN(_08866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17739_ (.A1(_08839_),
    .A2(_08866_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17740_ (.A1(_08576_),
    .A2(_08626_),
    .B(_08638_),
    .ZN(_08867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17741_ (.A1(_08655_),
    .A2(_00385_),
    .ZN(_08868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17742_ (.A1(_08867_),
    .A2(_08868_),
    .A3(_08614_),
    .ZN(_08869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17743_ (.I(_15594_),
    .ZN(_08870_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17744_ (.A1(_08621_),
    .A2(_08870_),
    .A3(_08693_),
    .ZN(_08871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17745_ (.A1(_08871_),
    .A2(_08662_),
    .ZN(_08872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17746_ (.A1(_08872_),
    .A2(_00386_),
    .ZN(_08873_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17747_ (.A1(_08869_),
    .A2(_08873_),
    .A3(_08664_),
    .ZN(_08874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17748_ (.A1(_08575_),
    .A2(_08631_),
    .ZN(_08875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17749_ (.A1(_08875_),
    .A2(_08657_),
    .ZN(_08876_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _17750_ (.I(_07638_),
    .Z(_08877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17751_ (.A1(_08646_),
    .A2(_08649_),
    .B(_08877_),
    .ZN(_08878_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17752_ (.A1(_08876_),
    .A2(_08878_),
    .A3(_08662_),
    .ZN(_08879_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17753_ (.A1(_08565_),
    .A2(_08654_),
    .A3(_08638_),
    .ZN(_08880_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17754_ (.A1(_08592_),
    .A2(_08726_),
    .A3(_08649_),
    .ZN(_08881_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17755_ (.A1(_08880_),
    .A2(_08881_),
    .A3(_08651_),
    .ZN(_08882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17756_ (.A1(_08879_),
    .A2(_08882_),
    .A3(_08728_),
    .ZN(_08883_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17757_ (.A1(_08874_),
    .A2(_08883_),
    .A3(_08643_),
    .ZN(_08884_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17758_ (.A1(_08609_),
    .A2(_08573_),
    .Z(_08885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17759_ (.A1(_08867_),
    .A2(_08885_),
    .B(_07647_),
    .ZN(_08886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17760_ (.A1(_08679_),
    .A2(_07629_),
    .ZN(_08887_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17761_ (.I(_08887_),
    .ZN(_08888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17762_ (.A1(_08888_),
    .A2(_08654_),
    .ZN(_08889_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17763_ (.A1(_08763_),
    .A2(_08889_),
    .A3(_08708_),
    .ZN(_08890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17764_ (.A1(_08886_),
    .A2(_08890_),
    .B(_08642_),
    .ZN(_08891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17765_ (.A1(_08604_),
    .A2(_08644_),
    .A3(_08671_),
    .ZN(_08892_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17766_ (.A1(_08628_),
    .A2(_08757_),
    .A3(_08892_),
    .ZN(_08893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17767_ (.A1(_08583_),
    .A2(_08674_),
    .ZN(_08894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17768_ (.A1(_08631_),
    .A2(_08894_),
    .B(_08671_),
    .ZN(_08895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17769_ (.A1(_08578_),
    .A2(_08688_),
    .B(_08580_),
    .ZN(_08896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17770_ (.A1(_08895_),
    .A2(_08896_),
    .B(_08877_),
    .ZN(_08897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17771_ (.A1(_08893_),
    .A2(_08897_),
    .ZN(_08898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17772_ (.A1(_08898_),
    .A2(_00387_),
    .ZN(_08899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17773_ (.A1(_08891_),
    .A2(_08899_),
    .ZN(_08900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17774_ (.A1(_08884_),
    .A2(_08900_),
    .B(_08668_),
    .ZN(_08901_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17775_ (.A1(_08670_),
    .A2(_07640_),
    .Z(_08902_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17776_ (.A1(_08583_),
    .A2(_15574_),
    .ZN(_08903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17777_ (.A1(_08903_),
    .A2(_08615_),
    .Z(_08904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17778_ (.A1(_08904_),
    .A2(_07647_),
    .ZN(_08905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17779_ (.A1(_08902_),
    .A2(_08905_),
    .Z(_08906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17780_ (.A1(_08588_),
    .A2(_08644_),
    .B(_08580_),
    .ZN(_08907_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17781_ (.I(_08662_),
    .ZN(_08908_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17782_ (.A1(_08907_),
    .A2(_08908_),
    .B(_08595_),
    .ZN(_08909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17783_ (.A1(_08906_),
    .A2(_08909_),
    .ZN(_08910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17784_ (.A1(_08910_),
    .A2(_08643_),
    .ZN(_08911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17785_ (.A1(_08601_),
    .A2(_08621_),
    .ZN(_08912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17786_ (.A1(_08590_),
    .A2(_08604_),
    .A3(_08693_),
    .ZN(_08913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17787_ (.A1(_08912_),
    .A2(_08596_),
    .A3(_08913_),
    .ZN(_08914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17788_ (.A1(_08706_),
    .A2(_08649_),
    .ZN(_08915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17789_ (.A1(_08806_),
    .A2(_07647_),
    .A3(_08915_),
    .ZN(_08916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17790_ (.A1(_08914_),
    .A2(_08916_),
    .B(_00386_),
    .ZN(_08917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17791_ (.A1(_08911_),
    .A2(_08917_),
    .B(_08668_),
    .ZN(_08918_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17792_ (.A1(_08680_),
    .A2(_08625_),
    .ZN(_08919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17793_ (.A1(_08919_),
    .A2(_08776_),
    .B(_08877_),
    .ZN(_08920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17794_ (.A1(_08803_),
    .A2(_08757_),
    .ZN(_08921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17795_ (.A1(_08920_),
    .A2(_08921_),
    .ZN(_08922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17796_ (.A1(_08922_),
    .A2(_08597_),
    .ZN(_08923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17797_ (.A1(_08739_),
    .A2(_08712_),
    .A3(_08651_),
    .ZN(_08924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17798_ (.A1(_08590_),
    .A2(_08705_),
    .ZN(_08925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17799_ (.A1(_08925_),
    .A2(_08627_),
    .ZN(_08926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17800_ (.A1(_08604_),
    .A2(_08599_),
    .A3(_08693_),
    .ZN(_08927_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17801_ (.A1(_08926_),
    .A2(_08927_),
    .A3(_08659_),
    .ZN(_08928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17802_ (.A1(_08924_),
    .A2(_08728_),
    .A3(_08928_),
    .ZN(_08929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17803_ (.A1(_08923_),
    .A2(_08929_),
    .B(_08643_),
    .ZN(_08930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17804_ (.A1(_08930_),
    .A2(_08918_),
    .ZN(_08931_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17805_ (.A1(_08901_),
    .A2(_08931_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17806_ (.A1(_08628_),
    .A2(_08694_),
    .A3(_08574_),
    .ZN(_08932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17807_ (.I(_08919_),
    .ZN(_08933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17808_ (.A1(net77),
    .A2(net30),
    .ZN(_08934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17809_ (.A1(_08587_),
    .A2(_08934_),
    .ZN(_08935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17810_ (.A1(_08935_),
    .A2(_08671_),
    .ZN(_08936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17811_ (.A1(_08933_),
    .A2(_08936_),
    .A3(_00386_),
    .ZN(_08937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17812_ (.A1(_08932_),
    .A2(_08937_),
    .A3(_08597_),
    .ZN(_08938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17813_ (.A1(_08656_),
    .A2(_15573_),
    .Z(_08939_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17814_ (.A1(_08939_),
    .A2(_08783_),
    .B(_08877_),
    .ZN(_08940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17815_ (.A1(_08940_),
    .A2(_07647_),
    .ZN(_08941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17816_ (.A1(_08681_),
    .A2(_08588_),
    .ZN(_08942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17817_ (.A1(_08676_),
    .A2(_08942_),
    .Z(_08943_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17818_ (.A1(_08943_),
    .A2(_08941_),
    .Z(_08944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17819_ (.A1(_08944_),
    .A2(_08643_),
    .A3(_08938_),
    .ZN(_08945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17820_ (.A1(_08622_),
    .A2(_08599_),
    .ZN(_08946_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17821_ (.A1(_08740_),
    .A2(_08757_),
    .ZN(_08947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17822_ (.A1(_08946_),
    .A2(_08947_),
    .B(_08728_),
    .ZN(_08948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17823_ (.A1(_08753_),
    .A2(_07640_),
    .Z(_08949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17824_ (.A1(_08949_),
    .A2(_08769_),
    .A3(_08568_),
    .ZN(_08950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17825_ (.A1(_08948_),
    .A2(_08950_),
    .ZN(_08951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17826_ (.A1(_08734_),
    .A2(_08688_),
    .ZN(_08952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17827_ (.A1(_08581_),
    .A2(_08952_),
    .A3(_08574_),
    .ZN(_08953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17828_ (.A1(_08759_),
    .A2(_08757_),
    .Z(_08954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17829_ (.A1(_08954_),
    .A2(_08795_),
    .B(_08596_),
    .ZN(_08955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17830_ (.A1(_08953_),
    .A2(_08955_),
    .ZN(_08956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17831_ (.A1(_08951_),
    .A2(_08956_),
    .A3(_00388_),
    .ZN(_08957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17832_ (.A1(_08668_),
    .A2(_08957_),
    .A3(_08945_),
    .ZN(_08958_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17833_ (.A1(_08566_),
    .A2(_08849_),
    .B(_08826_),
    .C(_08659_),
    .ZN(_08959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17834_ (.A1(_08782_),
    .A2(_08877_),
    .Z(_08960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17835_ (.A1(_08740_),
    .A2(net30),
    .ZN(_08961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17836_ (.A1(_08960_),
    .A2(_08731_),
    .A3(_08961_),
    .ZN(_08962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17837_ (.A1(_08959_),
    .A2(_08597_),
    .A3(_08962_),
    .ZN(_08963_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17838_ (.A1(_08701_),
    .A2(_08627_),
    .B(_07640_),
    .ZN(_08964_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17839_ (.I(_08964_),
    .ZN(_08965_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17840_ (.A1(_08783_),
    .A2(_08706_),
    .ZN(_08966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17841_ (.A1(_08965_),
    .A2(_08966_),
    .B(_08596_),
    .ZN(_08967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17842_ (.A1(_08592_),
    .A2(_08656_),
    .ZN(_08968_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17843_ (.A1(_08968_),
    .A2(_08661_),
    .Z(_08969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17844_ (.A1(_08651_),
    .A2(_08683_),
    .A3(_08969_),
    .ZN(_08970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17845_ (.A1(_08967_),
    .A2(_08970_),
    .B(_08698_),
    .ZN(_08971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17846_ (.A1(_08971_),
    .A2(_08963_),
    .ZN(_08972_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17847_ (.A1(_08686_),
    .A2(_08634_),
    .A3(_08580_),
    .ZN(_08973_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17848_ (.A1(_08936_),
    .A2(_08757_),
    .A3(_08973_),
    .Z(_08974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17849_ (.A1(_08770_),
    .A2(_08840_),
    .B(_08659_),
    .ZN(_08975_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17850_ (.A1(_08974_),
    .A2(_08975_),
    .B(_08664_),
    .ZN(_08976_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17851_ (.A1(_08625_),
    .A2(_15603_),
    .B(_08649_),
    .ZN(_08977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17852_ (.A1(_08772_),
    .A2(_08977_),
    .A3(_08651_),
    .ZN(_08978_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17853_ (.A1(_08569_),
    .A2(_08877_),
    .ZN(_08979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17854_ (.A1(_08979_),
    .A2(_08680_),
    .B(_08596_),
    .ZN(_08980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17855_ (.A1(_08978_),
    .A2(_08980_),
    .B(_08642_),
    .ZN(_08981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17856_ (.A1(_08976_),
    .A2(_08981_),
    .ZN(_08982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17857_ (.A1(_08972_),
    .A2(_08982_),
    .A3(_00389_),
    .ZN(_08983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17858_ (.A1(_08983_),
    .A2(_08958_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17859_ (.A1(_08965_),
    .A2(_08600_),
    .B(_08698_),
    .ZN(_08984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17860_ (.A1(_08621_),
    .A2(_08627_),
    .ZN(_08985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17861_ (.A1(_08985_),
    .A2(_08894_),
    .ZN(_08986_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17862_ (.A1(_08789_),
    .A2(_08986_),
    .Z(_08987_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17863_ (.A1(_08984_),
    .A2(_08987_),
    .B(_00389_),
    .ZN(_08988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17864_ (.A1(_08610_),
    .A2(net79),
    .ZN(_08989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17865_ (.A1(_08888_),
    .A2(_08588_),
    .ZN(_08990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17866_ (.A1(_08989_),
    .A2(_08990_),
    .B(_08696_),
    .ZN(_08991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17867_ (.A1(_00385_),
    .A2(net77),
    .ZN(_08992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17868_ (.A1(_08624_),
    .A2(_08992_),
    .B(_08659_),
    .ZN(_08993_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17869_ (.A1(_08991_),
    .A2(_08993_),
    .B(_08698_),
    .ZN(_08994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17870_ (.A1(_08988_),
    .A2(_08994_),
    .B(_08597_),
    .ZN(_08995_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17871_ (.A1(_08601_),
    .A2(_08612_),
    .Z(_08996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17872_ (.A1(_08996_),
    .A2(_08571_),
    .B(_08696_),
    .ZN(_08997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17873_ (.A1(_08751_),
    .A2(_08621_),
    .Z(_08998_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17874_ (.A1(_08682_),
    .A2(_08679_),
    .A3(_08656_),
    .Z(_08999_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17875_ (.A1(_08998_),
    .A2(_08999_),
    .B(_08757_),
    .ZN(_09000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17876_ (.A1(_08997_),
    .A2(_09000_),
    .A3(_08698_),
    .ZN(_09001_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17877_ (.A1(_08579_),
    .A2(_08645_),
    .A3(_08656_),
    .Z(_09002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17878_ (.A1(_08616_),
    .A2(_08934_),
    .ZN(_09003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17879_ (.A1(_09002_),
    .A2(_09003_),
    .A3(_08757_),
    .ZN(_09004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17880_ (.A1(_08615_),
    .A2(net77),
    .ZN(_09005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17881_ (.A1(_09005_),
    .A2(net30),
    .ZN(_09006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17882_ (.A1(_08568_),
    .A2(_09006_),
    .ZN(_09007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17883_ (.A1(_09007_),
    .A2(_08696_),
    .ZN(_09008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17884_ (.A1(_09004_),
    .A2(_08642_),
    .A3(_09008_),
    .ZN(_09009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17885_ (.A1(_09001_),
    .A2(_09009_),
    .ZN(_09010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17886_ (.A1(_09010_),
    .A2(_00389_),
    .ZN(_09011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17887_ (.A1(_08995_),
    .A2(_09011_),
    .ZN(_09012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17888_ (.A1(_07639_),
    .A2(_08894_),
    .ZN(_09013_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17889_ (.A1(_08734_),
    .A2(_09013_),
    .Z(_09014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17890_ (.A1(_09014_),
    .A2(_07654_),
    .Z(_09015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17891_ (.A1(_08604_),
    .A2(_08671_),
    .ZN(_09016_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17892_ (.A1(_08926_),
    .A2(_08614_),
    .A3(_09016_),
    .ZN(_09017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17893_ (.A1(_09015_),
    .A2(_09017_),
    .B(_08667_),
    .ZN(_09018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17894_ (.A1(_08654_),
    .A2(_07631_),
    .Z(_09019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17895_ (.A1(_09019_),
    .A2(_08648_),
    .ZN(_09020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17896_ (.A1(_08814_),
    .A2(_08657_),
    .ZN(_09021_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17897_ (.A1(_09020_),
    .A2(_08614_),
    .A3(_09021_),
    .ZN(_09022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17898_ (.A1(_08796_),
    .A2(_08686_),
    .ZN(_09023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17899_ (.A1(_08842_),
    .A2(_09023_),
    .ZN(_09024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17900_ (.A1(_09022_),
    .A2(_09024_),
    .A3(_08643_),
    .ZN(_09025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17901_ (.A1(_09025_),
    .A2(_09018_),
    .B(_00387_),
    .ZN(_09026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17902_ (.A1(_08746_),
    .A2(_08726_),
    .ZN(_09027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17903_ (.A1(_09027_),
    .A2(_08581_),
    .A3(_08574_),
    .ZN(_09028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17904_ (.A1(_08645_),
    .A2(_00385_),
    .ZN(_09029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17905_ (.A1(_08815_),
    .A2(_08764_),
    .A3(_09029_),
    .ZN(_09030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17906_ (.A1(_09028_),
    .A2(_00388_),
    .A3(_09030_),
    .ZN(_09031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17907_ (.A1(_08736_),
    .A2(_08690_),
    .ZN(_09032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17908_ (.I(_08904_),
    .ZN(_09033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17909_ (.A1(_09032_),
    .A2(_08815_),
    .A3(_09033_),
    .ZN(_09034_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17910_ (.A1(net84),
    .A2(_08577_),
    .B(_08693_),
    .ZN(_09035_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17911_ (.A1(_15583_),
    .A2(_08657_),
    .B(_09035_),
    .C(_08696_),
    .ZN(_09036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17912_ (.A1(_09034_),
    .A2(_09036_),
    .A3(_08643_),
    .ZN(_09037_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17913_ (.A1(_09031_),
    .A2(_09037_),
    .A3(_08668_),
    .ZN(_09038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17914_ (.A1(_09026_),
    .A2(_09038_),
    .ZN(_09039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17915_ (.A1(_09012_),
    .A2(_09039_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17916_ (.I(_08654_),
    .ZN(_09040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17917_ (.A1(_09040_),
    .A2(_08671_),
    .ZN(_09041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17918_ (.A1(_08926_),
    .A2(_08877_),
    .A3(_09041_),
    .ZN(_09042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17919_ (.A1(_08725_),
    .A2(_08607_),
    .ZN(_09043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17920_ (.A1(_09042_),
    .A2(_09043_),
    .ZN(_09044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17921_ (.A1(_09044_),
    .A2(_08664_),
    .ZN(_09045_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17922_ (.A1(_08576_),
    .A2(_08656_),
    .A3(_08626_),
    .Z(_09046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17923_ (.A1(_08588_),
    .A2(_08894_),
    .A3(_08693_),
    .ZN(_09047_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17924_ (.A1(_09046_),
    .A2(_08696_),
    .A3(_09047_),
    .ZN(_09048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17925_ (.A1(_08623_),
    .A2(_08627_),
    .ZN(_09049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17926_ (.A1(_09049_),
    .A2(_08968_),
    .ZN(_09050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17927_ (.A1(_07640_),
    .A2(_08575_),
    .Z(_09051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17928_ (.A1(_09050_),
    .A2(_09051_),
    .B(_08595_),
    .ZN(_09052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17929_ (.A1(_09048_),
    .A2(_09052_),
    .ZN(_09053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17930_ (.A1(_09045_),
    .A2(_09053_),
    .A3(_00388_),
    .ZN(_09054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17931_ (.A1(_08690_),
    .A2(_08671_),
    .ZN(_09055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17932_ (.A1(_08942_),
    .A2(_09055_),
    .ZN(_09056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17933_ (.A1(_09056_),
    .A2(_08659_),
    .ZN(_09057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17934_ (.A1(_08823_),
    .A2(_08595_),
    .Z(_09058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17935_ (.A1(_09057_),
    .A2(_09058_),
    .B(_08698_),
    .ZN(_09059_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17936_ (.A1(_09040_),
    .A2(_08600_),
    .B(_08749_),
    .ZN(_09060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17937_ (.A1(_08567_),
    .A2(_15593_),
    .Z(_09061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17938_ (.A1(_08990_),
    .A2(_08877_),
    .A3(_09061_),
    .ZN(_09062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17939_ (.A1(_09060_),
    .A2(_09062_),
    .ZN(_09063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17940_ (.A1(_09063_),
    .A2(_08728_),
    .ZN(_09064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17941_ (.A1(_09059_),
    .A2(_09064_),
    .ZN(_09065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17942_ (.A1(_09065_),
    .A2(_09054_),
    .ZN(_09066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17943_ (.A1(_09066_),
    .A2(_08668_),
    .ZN(_09067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17944_ (.A1(_08888_),
    .A2(_08592_),
    .ZN(_09068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17945_ (.A1(net84),
    .A2(_08577_),
    .ZN(_09069_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17946_ (.A1(_09069_),
    .A2(_08671_),
    .ZN(_09070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17947_ (.I(_09070_),
    .ZN(_09071_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17948_ (.A1(_09068_),
    .A2(_08651_),
    .A3(_08670_),
    .A4(_09071_),
    .Z(_09072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17949_ (.A1(_08622_),
    .A2(_08688_),
    .ZN(_09073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17950_ (.A1(_09073_),
    .A2(_08708_),
    .A3(_08926_),
    .ZN(_09074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17951_ (.A1(_09074_),
    .A2(_08597_),
    .ZN(_09075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17952_ (.A1(_08833_),
    .A2(_00385_),
    .ZN(_09076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17953_ (.A1(_08949_),
    .A2(_08915_),
    .A3(_09076_),
    .ZN(_09077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17954_ (.A1(_08935_),
    .A2(_08649_),
    .ZN(_09078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17955_ (.A1(net78),
    .A2(_08656_),
    .ZN(_09079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17956_ (.A1(_09079_),
    .A2(_08573_),
    .Z(_09080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17957_ (.A1(_09078_),
    .A2(_09080_),
    .B(_08596_),
    .ZN(_09081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17958_ (.A1(_09077_),
    .A2(_09081_),
    .ZN(_09082_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17959_ (.A1(_09072_),
    .A2(_09075_),
    .B(_00388_),
    .C(_09082_),
    .ZN(_09083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17960_ (.A1(_08586_),
    .A2(net79),
    .ZN(_09084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17961_ (.A1(_08855_),
    .A2(_07640_),
    .ZN(_09085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17962_ (.I(_09085_),
    .ZN(_09086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17963_ (.A1(_09084_),
    .A2(_09086_),
    .B(_08596_),
    .ZN(_09087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17964_ (.A1(_08610_),
    .A2(_08588_),
    .ZN(_09088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17965_ (.A1(_08796_),
    .A2(_08654_),
    .ZN(_09089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17966_ (.A1(_09088_),
    .A2(_09089_),
    .A3(_08696_),
    .ZN(_09090_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17967_ (.A1(_09087_),
    .A2(_09090_),
    .B(_08698_),
    .ZN(_09091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17968_ (.A1(_08672_),
    .A2(_08757_),
    .Z(_09092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17969_ (.I(_08849_),
    .ZN(_09093_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17970_ (.A1(_09093_),
    .A2(_08653_),
    .ZN(_09094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17971_ (.A1(_09092_),
    .A2(_09094_),
    .B(_08728_),
    .ZN(_09095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17972_ (.A1(_09093_),
    .A2(_08575_),
    .ZN(_09096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17973_ (.A1(_09073_),
    .A2(_09096_),
    .A3(_08614_),
    .ZN(_09097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17974_ (.A1(_09095_),
    .A2(_09097_),
    .ZN(_09098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17975_ (.A1(_09091_),
    .A2(_09098_),
    .B(_08668_),
    .ZN(_09099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17976_ (.A1(_09083_),
    .A2(_09099_),
    .ZN(_09100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17977_ (.A1(_09067_),
    .A2(_09100_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17978_ (.A1(_08637_),
    .A2(_08671_),
    .ZN(_09101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17979_ (.A1(_08849_),
    .A2(_09101_),
    .ZN(_09102_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17980_ (.A1(_09102_),
    .A2(_08757_),
    .A3(_09041_),
    .Z(_09103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17981_ (.A1(_08578_),
    .A2(_08580_),
    .ZN(_09104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17982_ (.A1(_09016_),
    .A2(_09104_),
    .A3(_08877_),
    .Z(_09105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17983_ (.A1(_09103_),
    .A2(_09105_),
    .B(_08597_),
    .ZN(_09106_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17984_ (.A1(_08985_),
    .A2(_08566_),
    .B(_08659_),
    .C(_09005_),
    .ZN(_09107_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17985_ (.A1(_08588_),
    .A2(_08637_),
    .A3(_08638_),
    .ZN(_09108_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17986_ (.A1(_08840_),
    .A2(_09108_),
    .A3(_08651_),
    .ZN(_09109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17987_ (.A1(_09107_),
    .A2(_09109_),
    .A3(_08728_),
    .ZN(_09110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17988_ (.A1(_09106_),
    .A2(_08668_),
    .A3(_09110_),
    .ZN(_09111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17989_ (.I(_08817_),
    .ZN(_09112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17990_ (.A1(_08627_),
    .A2(_15603_),
    .ZN(_09113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17991_ (.A1(_09113_),
    .A2(_08573_),
    .ZN(_09114_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17992_ (.A1(_09112_),
    .A2(_09114_),
    .ZN(_09115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17993_ (.A1(_08661_),
    .A2(_08657_),
    .ZN(_09116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17994_ (.A1(_09115_),
    .A2(_09116_),
    .B(_08728_),
    .ZN(_09117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17995_ (.A1(_09019_),
    .A2(_08660_),
    .ZN(_09118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17996_ (.A1(_08749_),
    .A2(_09118_),
    .A3(_08851_),
    .ZN(_09119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17997_ (.A1(_09117_),
    .A2(_09119_),
    .ZN(_09120_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17998_ (.A1(_08832_),
    .A2(_07631_),
    .B(_07638_),
    .ZN(_09121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17999_ (.A1(_07631_),
    .A2(_08577_),
    .Z(_09122_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18000_ (.A1(_09121_),
    .A2(_09122_),
    .Z(_09123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18001_ (.A1(_09123_),
    .A2(_07647_),
    .Z(_09124_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18002_ (.A1(_08769_),
    .A2(_08676_),
    .A3(_08568_),
    .ZN(_09125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18003_ (.A1(_09124_),
    .A2(_09125_),
    .ZN(_09126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18004_ (.A1(_09120_),
    .A2(_09126_),
    .A3(_00389_),
    .ZN(_09127_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18005_ (.A1(_09111_),
    .A2(_09127_),
    .A3(_08643_),
    .ZN(_09128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18006_ (.A1(_08687_),
    .A2(_08637_),
    .ZN(_09129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18007_ (.A1(_08933_),
    .A2(_09129_),
    .A3(_08708_),
    .ZN(_09130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18008_ (.A1(_09019_),
    .A2(_08690_),
    .ZN(_09131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18009_ (.A1(_15596_),
    .A2(_08633_),
    .ZN(_09132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18010_ (.A1(_09132_),
    .A2(_09069_),
    .ZN(_09133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18011_ (.A1(_09133_),
    .A2(_08657_),
    .ZN(_09134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18012_ (.A1(_09131_),
    .A2(_08614_),
    .A3(_09134_),
    .ZN(_09135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18013_ (.A1(_09130_),
    .A2(_09135_),
    .A3(_00387_),
    .ZN(_09136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18014_ (.A1(_08657_),
    .A2(_15580_),
    .ZN(_09137_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18015_ (.A1(_09078_),
    .A2(_08708_),
    .A3(_09137_),
    .ZN(_09138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18016_ (.A1(_08565_),
    .A2(_08693_),
    .B(_09132_),
    .ZN(_09139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18017_ (.A1(_09139_),
    .A2(_09121_),
    .Z(_09140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18018_ (.A1(_09138_),
    .A2(_09140_),
    .A3(_08664_),
    .ZN(_09141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18019_ (.A1(_09136_),
    .A2(_09141_),
    .A3(_00389_),
    .ZN(_09142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18020_ (.A1(_08968_),
    .A2(_08877_),
    .Z(_09143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18021_ (.A1(_09143_),
    .A2(_08942_),
    .B(_08596_),
    .ZN(_09144_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18022_ (.A1(_08616_),
    .A2(_09070_),
    .B(_08682_),
    .ZN(_09145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18023_ (.A1(_09145_),
    .A2(_08878_),
    .ZN(_09146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18024_ (.A1(_09144_),
    .A2(_09146_),
    .B(_00389_),
    .ZN(_09147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18025_ (.A1(_08847_),
    .A2(_09068_),
    .A3(_08614_),
    .ZN(_09148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18026_ (.A1(_08659_),
    .A2(_08730_),
    .A3(_08913_),
    .ZN(_09149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18027_ (.A1(_09148_),
    .A2(_08664_),
    .A3(_09149_),
    .ZN(_09150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18028_ (.A1(_09150_),
    .A2(_09147_),
    .ZN(_09151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18029_ (.A1(_09142_),
    .A2(_09151_),
    .A3(_00388_),
    .ZN(_09152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18030_ (.A1(_09152_),
    .A2(_09128_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18031_ (.A1(_07550_),
    .A2(_07542_),
    .B(_07553_),
    .ZN(_15605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18032_ (.A1(_07559_),
    .A2(_07467_),
    .B(_07561_),
    .ZN(_09153_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _18033_ (.I(_09153_),
    .Z(_09154_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _18034_ (.I(_09154_),
    .Z(_15625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18035_ (.A1(_07468_),
    .A2(_07541_),
    .B(_07545_),
    .ZN(_15606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18036_ (.A1(_15616_),
    .A2(_09153_),
    .ZN(_09155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18037_ (.I(_09155_),
    .ZN(_09156_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18038_ (.I(_07570_),
    .Z(_09157_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18039_ (.I(_09157_),
    .Z(_09158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18040_ (.A1(_09156_),
    .A2(_09158_),
    .ZN(_09159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18041_ (.I(_15608_),
    .ZN(_09160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18042_ (.A1(_09160_),
    .A2(_07563_),
    .ZN(_09161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18043_ (.I(_09161_),
    .ZN(_09162_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18044_ (.I(_09157_),
    .Z(_09163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18045_ (.A1(_09162_),
    .A2(_09163_),
    .ZN(_09164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18046_ (.A1(_09154_),
    .A2(_09160_),
    .ZN(_09165_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18047_ (.I(_07571_),
    .Z(_09166_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18048_ (.I(_09166_),
    .Z(_09167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18049_ (.A1(_09165_),
    .A2(_09167_),
    .ZN(_09168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18050_ (.A1(_09159_),
    .A2(_09164_),
    .A3(_09168_),
    .ZN(_09169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18051_ (.A1(_09169_),
    .A2(_00401_),
    .ZN(_09170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18052_ (.I(_15621_),
    .ZN(_09171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18053_ (.A1(_15630_),
    .A2(_09171_),
    .Z(_09172_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18054_ (.I(_15617_),
    .ZN(_09173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18055_ (.A1(_09154_),
    .A2(_09173_),
    .ZN(_09174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18056_ (.I(_09174_),
    .ZN(_09175_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18057_ (.I(_09163_),
    .Z(_09176_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18058_ (.A1(_09172_),
    .A2(_09175_),
    .B(_09176_),
    .ZN(_09177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18059_ (.A1(_07571_),
    .A2(_09161_),
    .ZN(_09178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18060_ (.I(_09178_),
    .ZN(_09179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18061_ (.A1(_15625_),
    .A2(_15621_),
    .ZN(_09180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18062_ (.A1(_09179_),
    .A2(_09180_),
    .ZN(_09181_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _18063_ (.I(_07578_),
    .ZN(_09182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18064_ (.I(_09182_),
    .Z(_09183_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18065_ (.I(_09183_),
    .Z(_09184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18066_ (.A1(_09177_),
    .A2(_09181_),
    .A3(_09184_),
    .ZN(_09185_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _18067_ (.I(_07586_),
    .ZN(_09186_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18068_ (.I(_09186_),
    .Z(_09187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18069_ (.A1(_09170_),
    .A2(_09185_),
    .A3(_09187_),
    .ZN(_09188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18070_ (.A1(_15630_),
    .A2(_09173_),
    .ZN(_09189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18071_ (.I(_09189_),
    .ZN(_09190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18072_ (.A1(_15625_),
    .A2(_09171_),
    .ZN(_09191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18073_ (.I(_09191_),
    .ZN(_09192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18074_ (.A1(_09190_),
    .A2(_09192_),
    .B(_00400_),
    .ZN(_09193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18075_ (.A1(_09161_),
    .A2(_09157_),
    .Z(_09194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18076_ (.A1(_09153_),
    .A2(_15607_),
    .ZN(_09195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18077_ (.A1(_09194_),
    .A2(_09195_),
    .ZN(_09196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18078_ (.A1(_09193_),
    .A2(_09196_),
    .A3(_09184_),
    .ZN(_09197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18079_ (.A1(_07563_),
    .A2(_15606_),
    .ZN(_09198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18080_ (.A1(_09198_),
    .A2(_09157_),
    .ZN(_09199_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18081_ (.I(_09199_),
    .ZN(_09200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18082_ (.A1(net88),
    .A2(net89),
    .ZN(_09201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18083_ (.A1(_09200_),
    .A2(_09201_),
    .ZN(_09202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18084_ (.A1(_09154_),
    .A2(net87),
    .ZN(_09203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18085_ (.A1(net88),
    .A2(net86),
    .ZN(_09204_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18086_ (.I(_09166_),
    .Z(_09205_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18087_ (.A1(_09203_),
    .A2(_09204_),
    .A3(_09205_),
    .ZN(_09206_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18088_ (.I(_07579_),
    .Z(_09207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18089_ (.A1(_09202_),
    .A2(_09206_),
    .A3(_09207_),
    .ZN(_09208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18090_ (.A1(_09197_),
    .A2(_09208_),
    .A3(_00402_),
    .ZN(_09209_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18091_ (.I(_00403_),
    .ZN(_09210_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18092_ (.I(_09210_),
    .Z(_09211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18093_ (.A1(_09188_),
    .A2(_09209_),
    .A3(_09211_),
    .ZN(_09212_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18094_ (.I(_00404_),
    .ZN(_09213_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18095_ (.I(_09213_),
    .Z(_09214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18096_ (.A1(_15611_),
    .A2(_09154_),
    .ZN(_09215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18097_ (.A1(_09215_),
    .A2(_09158_),
    .Z(_09216_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18098_ (.I(_07578_),
    .Z(_09217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18099_ (.A1(_09216_),
    .A2(_09217_),
    .ZN(_09218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18100_ (.A1(_09154_),
    .A2(_15612_),
    .ZN(_09219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18101_ (.A1(_09219_),
    .A2(_07572_),
    .ZN(_09220_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18102_ (.I(_09220_),
    .ZN(_09221_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _18103_ (.I(_07563_),
    .Z(_09222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18104_ (.I(_15614_),
    .ZN(_09223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18105_ (.A1(_09222_),
    .A2(_09223_),
    .ZN(_09224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18106_ (.A1(_09221_),
    .A2(_09224_),
    .ZN(_09225_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18107_ (.I(_09186_),
    .Z(_09226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18108_ (.A1(_09218_),
    .A2(_09225_),
    .B(_09226_),
    .ZN(_09227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18109_ (.A1(net88),
    .A2(_15630_),
    .B(_09166_),
    .ZN(_09228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18110_ (.A1(_09228_),
    .A2(_09219_),
    .ZN(_09229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18111_ (.I(_15609_),
    .ZN(_09230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18112_ (.A1(_09154_),
    .A2(_09230_),
    .ZN(_09231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18113_ (.A1(_09231_),
    .A2(_09166_),
    .ZN(_09232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18114_ (.I(_09232_),
    .ZN(_09233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18115_ (.A1(_09233_),
    .A2(_09161_),
    .ZN(_09234_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18116_ (.I(_07578_),
    .Z(_09235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18117_ (.A1(_09229_),
    .A2(_09234_),
    .A3(_09235_),
    .ZN(_09236_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18118_ (.I(_09210_),
    .Z(_09237_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18119_ (.A1(_09227_),
    .A2(_09236_),
    .B(_09237_),
    .ZN(_09238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18120_ (.A1(_09222_),
    .A2(_15623_),
    .Z(_09239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18121_ (.A1(_09239_),
    .A2(_09163_),
    .ZN(_09240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18122_ (.A1(_09159_),
    .A2(_09240_),
    .Z(_09241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18123_ (.A1(_09166_),
    .A2(net87),
    .Z(_09242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18124_ (.A1(_09242_),
    .A2(_15625_),
    .ZN(_09243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18125_ (.I(_15607_),
    .ZN(_09244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18126_ (.A1(_09222_),
    .A2(_09244_),
    .ZN(_09245_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18127_ (.I(_09245_),
    .ZN(_09246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18128_ (.A1(_09246_),
    .A2(_09205_),
    .B(_07578_),
    .ZN(_09247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18129_ (.A1(_09241_),
    .A2(_09243_),
    .A3(_09247_),
    .ZN(_09248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18130_ (.A1(net89),
    .A2(_09222_),
    .ZN(_09249_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18131_ (.A1(_09249_),
    .A2(_09157_),
    .Z(_09250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18132_ (.A1(_09250_),
    .A2(_09219_),
    .ZN(_09251_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18133_ (.I(_09166_),
    .Z(_09252_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18134_ (.A1(_09215_),
    .A2(_09252_),
    .Z(_09253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18135_ (.A1(_09222_),
    .A2(_09230_),
    .ZN(_09254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18136_ (.A1(_09253_),
    .A2(_09254_),
    .ZN(_09255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18137_ (.A1(_09251_),
    .A2(_09255_),
    .A3(_09207_),
    .ZN(_09256_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18138_ (.I(_09186_),
    .Z(_09257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18139_ (.A1(_09248_),
    .A2(_09256_),
    .A3(_09257_),
    .ZN(_09258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18140_ (.A1(_09238_),
    .A2(_09258_),
    .ZN(_09259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18141_ (.A1(_09212_),
    .A2(_09214_),
    .A3(_09259_),
    .ZN(_09260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18142_ (.A1(_09154_),
    .A2(_15614_),
    .ZN(_09261_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18143_ (.A1(_09261_),
    .A2(_09166_),
    .Z(_09262_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18144_ (.A1(_09247_),
    .A2(_09243_),
    .A3(_09262_),
    .ZN(_09263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18145_ (.A1(_09262_),
    .A2(_07579_),
    .Z(_09264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18146_ (.A1(_09222_),
    .A2(_15619_),
    .ZN(_09265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18147_ (.I(_09265_),
    .ZN(_09266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18148_ (.A1(_09266_),
    .A2(_09158_),
    .ZN(_09267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18149_ (.A1(_09267_),
    .A2(_09178_),
    .Z(_09268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18150_ (.A1(_09264_),
    .A2(_09268_),
    .ZN(_09269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18151_ (.A1(_09263_),
    .A2(_09269_),
    .A3(_09257_),
    .ZN(_09270_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18152_ (.I(_09163_),
    .Z(_09271_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18153_ (.A1(_09239_),
    .A2(_09192_),
    .B(_09271_),
    .ZN(_09272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18154_ (.A1(_09224_),
    .A2(_07572_),
    .ZN(_09273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18155_ (.A1(_09272_),
    .A2(_09207_),
    .A3(_09273_),
    .ZN(_09274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18156_ (.A1(net88),
    .A2(_15630_),
    .ZN(_09275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18157_ (.A1(_15625_),
    .A2(_15617_),
    .ZN(_09276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18158_ (.A1(_09275_),
    .A2(_09276_),
    .A3(_09167_),
    .ZN(_09277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18159_ (.A1(_09222_),
    .A2(net86),
    .ZN(_09278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18160_ (.A1(_15608_),
    .A2(_09153_),
    .ZN(_09279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18161_ (.A1(_09278_),
    .A2(_09279_),
    .A3(_09158_),
    .ZN(_09280_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18162_ (.I(_09182_),
    .Z(_09281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18163_ (.A1(_09277_),
    .A2(_09280_),
    .A3(_09281_),
    .ZN(_09282_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18164_ (.I(_07586_),
    .Z(_09283_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18165_ (.A1(_09274_),
    .A2(_09282_),
    .A3(_09283_),
    .ZN(_09284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18166_ (.A1(_09270_),
    .A2(_09284_),
    .A3(_00403_),
    .ZN(_09285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18167_ (.I(_15619_),
    .ZN(_09286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18168_ (.A1(_09154_),
    .A2(_09286_),
    .ZN(_09287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18169_ (.A1(_09287_),
    .A2(_09166_),
    .ZN(_09288_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18170_ (.I(_09288_),
    .ZN(_09289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18171_ (.A1(_09222_),
    .A2(_15612_),
    .ZN(_09290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18172_ (.A1(_09289_),
    .A2(_09290_),
    .ZN(_09291_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18173_ (.A1(_09291_),
    .A2(_09281_),
    .A3(_09240_),
    .ZN(_09292_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18174_ (.I(_15612_),
    .ZN(_09293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18175_ (.A1(_09222_),
    .A2(_09293_),
    .ZN(_09294_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18176_ (.A1(_09294_),
    .A2(_09166_),
    .Z(_09295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18177_ (.A1(_09295_),
    .A2(_07578_),
    .Z(_09296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18178_ (.A1(_09239_),
    .A2(_09252_),
    .ZN(_09297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18179_ (.A1(_09175_),
    .A2(_09158_),
    .ZN(_09298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18180_ (.A1(_09297_),
    .A2(_09298_),
    .Z(_09299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18181_ (.A1(_09296_),
    .A2(_09299_),
    .ZN(_09300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18182_ (.A1(_09292_),
    .A2(_09300_),
    .A3(_09283_),
    .ZN(_09301_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18183_ (.A1(_09203_),
    .A2(_09290_),
    .A3(_09271_),
    .Z(_09302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18184_ (.A1(_09172_),
    .A2(_09167_),
    .B(_07578_),
    .ZN(_09303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18185_ (.A1(_09303_),
    .A2(_09243_),
    .ZN(_09304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18186_ (.I(_09279_),
    .ZN(_09305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18187_ (.A1(_09305_),
    .A2(_09271_),
    .ZN(_09306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18188_ (.I(_15633_),
    .ZN(_09307_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18189_ (.A1(_09158_),
    .A2(_09307_),
    .B(_07578_),
    .ZN(_09308_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18190_ (.I(_09308_),
    .ZN(_09309_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18191_ (.I(_07586_),
    .Z(_09310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18192_ (.A1(_09306_),
    .A2(_09309_),
    .B(_09310_),
    .ZN(_09311_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18193_ (.A1(_09302_),
    .A2(_09304_),
    .B(_09311_),
    .ZN(_09312_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18194_ (.A1(_09301_),
    .A2(_09211_),
    .A3(_09312_),
    .ZN(_09313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18195_ (.A1(_09285_),
    .A2(_09313_),
    .A3(_00404_),
    .ZN(_09314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18196_ (.A1(_09260_),
    .A2(_09314_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18197_ (.A1(_09295_),
    .A2(_09262_),
    .Z(_09315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18198_ (.A1(_09254_),
    .A2(_09165_),
    .A3(_09167_),
    .ZN(_09316_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18199_ (.I(_09183_),
    .Z(_09317_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18200_ (.A1(_09315_),
    .A2(_09316_),
    .A3(_09317_),
    .ZN(_09318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18201_ (.A1(_09278_),
    .A2(_09163_),
    .Z(_09319_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18202_ (.A1(_07560_),
    .A2(_07562_),
    .A3(_09223_),
    .ZN(_09320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18203_ (.A1(_09319_),
    .A2(_09320_),
    .ZN(_09321_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18204_ (.A1(_09157_),
    .A2(_15626_),
    .Z(_09322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18205_ (.A1(_09322_),
    .A2(_09217_),
    .ZN(_09323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18206_ (.I(_09323_),
    .ZN(_09324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18207_ (.A1(_09321_),
    .A2(_09324_),
    .B(_09310_),
    .ZN(_09325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18208_ (.A1(_09318_),
    .A2(_09325_),
    .B(_00403_),
    .ZN(_09326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18209_ (.A1(_09224_),
    .A2(_09163_),
    .ZN(_09327_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18210_ (.I(_09327_),
    .ZN(_09328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18211_ (.A1(_09328_),
    .A2(_09203_),
    .ZN(_09329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18212_ (.A1(_09179_),
    .A2(_09215_),
    .ZN(_09330_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18213_ (.A1(_09329_),
    .A2(_09330_),
    .A3(_00401_),
    .ZN(_09331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18214_ (.A1(_09319_),
    .A2(_09201_),
    .ZN(_09332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18215_ (.A1(_15625_),
    .A2(_09293_),
    .ZN(_09333_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18216_ (.I(_09157_),
    .Z(_09334_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18217_ (.A1(_09333_),
    .A2(_09334_),
    .Z(_09335_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18218_ (.A1(_09332_),
    .A2(_09317_),
    .A3(_09335_),
    .ZN(_09336_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18219_ (.A1(_09331_),
    .A2(_09336_),
    .A3(_00402_),
    .ZN(_09337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18220_ (.A1(_09326_),
    .A2(_09337_),
    .ZN(_09338_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18221_ (.A1(_15630_),
    .A2(_15614_),
    .Z(_09339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18222_ (.A1(_09339_),
    .A2(_09176_),
    .B(_09217_),
    .ZN(_09340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18223_ (.A1(_09195_),
    .A2(_09166_),
    .ZN(_09341_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18224_ (.I(_09341_),
    .ZN(_09342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18225_ (.A1(_09222_),
    .A2(_15608_),
    .ZN(_09343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18226_ (.A1(_09342_),
    .A2(_09343_),
    .ZN(_09344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18227_ (.A1(_09340_),
    .A2(_09344_),
    .B(_09226_),
    .ZN(_09345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18228_ (.A1(_09233_),
    .A2(_09249_),
    .ZN(_09346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18229_ (.A1(_09246_),
    .A2(_09163_),
    .ZN(_09347_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18230_ (.A1(_09346_),
    .A2(_00401_),
    .A3(_09347_),
    .ZN(_09348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18231_ (.A1(_09345_),
    .A2(_09348_),
    .B(_09237_),
    .ZN(_09349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18232_ (.A1(_09228_),
    .A2(_09279_),
    .ZN(_09350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18233_ (.A1(net89),
    .A2(net87),
    .ZN(_09351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18234_ (.A1(_09253_),
    .A2(_09351_),
    .ZN(_09352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18235_ (.A1(_09350_),
    .A2(_09352_),
    .A3(_09317_),
    .ZN(_09353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18236_ (.I(_09203_),
    .ZN(_09354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18237_ (.A1(_09354_),
    .A2(_09334_),
    .B(_09182_),
    .ZN(_09355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18238_ (.A1(_09320_),
    .A2(_09252_),
    .ZN(_09356_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18239_ (.I(_09343_),
    .ZN(_09357_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18240_ (.A1(_09356_),
    .A2(_09357_),
    .Z(_09358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18241_ (.A1(_09172_),
    .A2(_09271_),
    .ZN(_09359_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18242_ (.A1(_09355_),
    .A2(_09358_),
    .A3(_09359_),
    .ZN(_09360_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18243_ (.A1(_09353_),
    .A2(_09360_),
    .A3(_09187_),
    .ZN(_09361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18244_ (.A1(_09349_),
    .A2(_09361_),
    .ZN(_09362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18245_ (.A1(_09338_),
    .A2(_09362_),
    .A3(_00404_),
    .ZN(_09363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18246_ (.A1(_09246_),
    .A2(_09252_),
    .ZN(_09364_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18247_ (.A1(_09364_),
    .A2(_07586_),
    .Z(_09365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18248_ (.A1(_09228_),
    .A2(_09180_),
    .ZN(_09366_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18249_ (.A1(_09365_),
    .A2(_09366_),
    .A3(_09335_),
    .ZN(_09367_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18250_ (.A1(_09273_),
    .A2(_09156_),
    .Z(_09368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18251_ (.A1(_15625_),
    .A2(net86),
    .ZN(_09369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18252_ (.A1(_09200_),
    .A2(_09369_),
    .ZN(_09370_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18253_ (.A1(_09368_),
    .A2(_09370_),
    .A3(_09226_),
    .ZN(_09371_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18254_ (.A1(_09367_),
    .A2(_09371_),
    .A3(_00401_),
    .ZN(_09372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18255_ (.A1(_09245_),
    .A2(_09174_),
    .B(_09252_),
    .ZN(_09373_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18256_ (.A1(_07586_),
    .A2(_15635_),
    .A3(_09334_),
    .ZN(_09374_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18257_ (.A1(_09373_),
    .A2(_09374_),
    .Z(_09375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18258_ (.A1(_09375_),
    .A2(_09317_),
    .B(_00403_),
    .ZN(_09376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18259_ (.A1(_09372_),
    .A2(_09376_),
    .B(_00404_),
    .ZN(_09377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18260_ (.A1(_09172_),
    .A2(_09252_),
    .ZN(_09378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18261_ (.A1(_07572_),
    .A2(_09305_),
    .ZN(_09379_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18262_ (.A1(_09378_),
    .A2(_09355_),
    .A3(_09240_),
    .A4(_09379_),
    .ZN(_09380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18263_ (.A1(_09200_),
    .A2(_09180_),
    .ZN(_09381_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18264_ (.A1(_09368_),
    .A2(_09381_),
    .A3(_09184_),
    .ZN(_09382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18265_ (.A1(_09380_),
    .A2(_00402_),
    .A3(_09382_),
    .ZN(_09383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18266_ (.A1(_09347_),
    .A2(_09183_),
    .Z(_09384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18267_ (.A1(_09178_),
    .A2(_09203_),
    .Z(_09385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18268_ (.A1(_09384_),
    .A2(_09385_),
    .B(_09310_),
    .ZN(_09386_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18269_ (.A1(_15630_),
    .A2(_15623_),
    .B(_09157_),
    .ZN(_09387_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18270_ (.I(_09387_),
    .ZN(_09388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18271_ (.A1(_09388_),
    .A2(_09254_),
    .ZN(_09389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18272_ (.A1(_09389_),
    .A2(_09344_),
    .A3(_09207_),
    .ZN(_09390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18273_ (.A1(_09386_),
    .A2(_09390_),
    .B(_09237_),
    .ZN(_09391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18274_ (.A1(_09383_),
    .A2(_09391_),
    .ZN(_09392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18275_ (.A1(_09377_),
    .A2(_09392_),
    .ZN(_09393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18276_ (.A1(_09363_),
    .A2(_09393_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18277_ (.A1(_09278_),
    .A2(_09219_),
    .A3(_09252_),
    .Z(_09394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18278_ (.I(_09231_),
    .ZN(_09395_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18279_ (.A1(_09327_),
    .A2(_09395_),
    .ZN(_09396_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18280_ (.A1(_09394_),
    .A2(_09396_),
    .B(_09235_),
    .ZN(_09397_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18281_ (.A1(_09294_),
    .A2(_09261_),
    .A3(_09205_),
    .ZN(_09398_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18282_ (.I(_09182_),
    .Z(_09399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18283_ (.A1(_09280_),
    .A2(_09398_),
    .A3(_09399_),
    .ZN(_09400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18284_ (.A1(_09397_),
    .A2(_09257_),
    .A3(_09400_),
    .ZN(_09401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18285_ (.A1(_09254_),
    .A2(_09195_),
    .A3(_09205_),
    .ZN(_09402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18286_ (.A1(_09219_),
    .A2(_09163_),
    .ZN(_09403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18287_ (.A1(_09402_),
    .A2(_09403_),
    .ZN(_09404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18288_ (.A1(_09404_),
    .A2(_09399_),
    .ZN(_09405_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18289_ (.A1(_09155_),
    .A2(_09343_),
    .A3(_09334_),
    .ZN(_09406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18290_ (.A1(_15625_),
    .A2(_15623_),
    .ZN(_09407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18291_ (.A1(_09198_),
    .A2(_09407_),
    .A3(_09167_),
    .ZN(_09408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18292_ (.A1(_09406_),
    .A2(_09408_),
    .A3(_09217_),
    .ZN(_09409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18293_ (.A1(_09405_),
    .A2(_09409_),
    .A3(_09283_),
    .ZN(_09410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18294_ (.A1(_09401_),
    .A2(_09410_),
    .A3(_09237_),
    .ZN(_09411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18295_ (.A1(_09262_),
    .A2(_09356_),
    .ZN(_09412_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18296_ (.A1(_09249_),
    .A2(_09182_),
    .Z(_09413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18297_ (.A1(_09267_),
    .A2(_09186_),
    .ZN(_09414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18298_ (.A1(_09412_),
    .A2(_09413_),
    .B(_09414_),
    .ZN(_09415_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18299_ (.A1(_09275_),
    .A2(_09252_),
    .A3(_09320_),
    .Z(_09416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18300_ (.A1(_09154_),
    .A2(_15609_),
    .ZN(_09417_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18301_ (.I(_09417_),
    .ZN(_09418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18302_ (.A1(_09418_),
    .A2(_09158_),
    .ZN(_09419_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18303_ (.I(_09419_),
    .ZN(_09420_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18304_ (.A1(_09416_),
    .A2(_09420_),
    .B(_09217_),
    .ZN(_09421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18305_ (.A1(_09415_),
    .A2(_09421_),
    .B(_09210_),
    .ZN(_09422_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18306_ (.A1(_09179_),
    .A2(_09279_),
    .Z(_09423_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18307_ (.A1(_09275_),
    .A2(_09158_),
    .A3(_09287_),
    .Z(_09424_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18308_ (.A1(_09423_),
    .A2(_09424_),
    .B(_09399_),
    .ZN(_09425_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18309_ (.A1(_09199_),
    .A2(_09418_),
    .B(_07578_),
    .ZN(_09426_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18310_ (.A1(_09155_),
    .A2(_09265_),
    .A3(_07572_),
    .Z(_09427_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18311_ (.A1(_09426_),
    .A2(_09427_),
    .Z(_09428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18312_ (.A1(_09283_),
    .A2(_09428_),
    .A3(_09425_),
    .ZN(_09429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18313_ (.A1(_09429_),
    .A2(_09422_),
    .ZN(_09430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18314_ (.A1(_09430_),
    .A2(_09411_),
    .ZN(_09431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18315_ (.A1(_09431_),
    .A2(_09214_),
    .ZN(_09432_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18316_ (.A1(_09157_),
    .A2(_15631_),
    .Z(_09433_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18317_ (.A1(_09403_),
    .A2(_09183_),
    .A3(_09433_),
    .Z(_09434_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18318_ (.A1(_09434_),
    .A2(_09283_),
    .ZN(_09435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18319_ (.A1(_09158_),
    .A2(_15628_),
    .ZN(_09436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18320_ (.A1(_09436_),
    .A2(_09217_),
    .ZN(_09437_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18321_ (.A1(_09394_),
    .A2(_09437_),
    .Z(_09438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18322_ (.A1(_09435_),
    .A2(_09438_),
    .B(_00403_),
    .ZN(_09439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18323_ (.A1(_09342_),
    .A2(_09198_),
    .Z(_09440_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18324_ (.A1(_09440_),
    .A2(_09399_),
    .A3(_09373_),
    .Z(_09441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18325_ (.A1(_09179_),
    .A2(_09320_),
    .ZN(_09442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18326_ (.A1(_09172_),
    .A2(_09271_),
    .B(_07579_),
    .ZN(_09443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18327_ (.A1(_09442_),
    .A2(_09443_),
    .B(_09226_),
    .ZN(_09444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18328_ (.A1(_09441_),
    .A2(_09444_),
    .ZN(_09445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18329_ (.A1(_09439_),
    .A2(_09445_),
    .B(_09214_),
    .ZN(_09446_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18330_ (.A1(_09201_),
    .A2(_09278_),
    .A3(_09205_),
    .ZN(_09447_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18331_ (.A1(_15635_),
    .A2(_00400_),
    .B(_09447_),
    .C(_09281_),
    .ZN(_09448_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18332_ (.A1(_09379_),
    .A2(_07579_),
    .Z(_09449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18333_ (.A1(_09250_),
    .A2(_09180_),
    .ZN(_09450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18334_ (.A1(_09190_),
    .A2(_00400_),
    .ZN(_09451_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18335_ (.A1(_09449_),
    .A2(_09450_),
    .A3(_09451_),
    .ZN(_09452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18336_ (.A1(_09448_),
    .A2(_09452_),
    .A3(_09187_),
    .ZN(_09453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18337_ (.A1(_09290_),
    .A2(_07572_),
    .Z(_09454_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18338_ (.I(_09454_),
    .ZN(_09455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18339_ (.I(_09165_),
    .ZN(_09456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18340_ (.A1(_09271_),
    .A2(_15633_),
    .ZN(_09457_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18341_ (.A1(_09455_),
    .A2(_09456_),
    .B(_09399_),
    .C(_09457_),
    .ZN(_09458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18342_ (.I(_09198_),
    .ZN(_09459_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18343_ (.A1(_09459_),
    .A2(_15628_),
    .B(_09167_),
    .ZN(_09460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18344_ (.A1(_09460_),
    .A2(_09235_),
    .A3(_09280_),
    .ZN(_09461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18345_ (.A1(_09458_),
    .A2(_09283_),
    .A3(_09461_),
    .ZN(_09462_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18346_ (.A1(_09453_),
    .A2(_09462_),
    .A3(_00403_),
    .ZN(_09463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18347_ (.A1(_09446_),
    .A2(_09463_),
    .ZN(_09464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18348_ (.A1(_09432_),
    .A2(_09464_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18349_ (.A1(_09200_),
    .A2(_09204_),
    .ZN(_09465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18350_ (.A1(_09155_),
    .A2(_09161_),
    .A3(_00400_),
    .ZN(_09466_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18351_ (.A1(_09465_),
    .A2(_09184_),
    .A3(_09466_),
    .ZN(_09467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18352_ (.I(_15628_),
    .ZN(_09468_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18353_ (.A1(_09198_),
    .A2(_09468_),
    .A3(_09334_),
    .ZN(_09469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18354_ (.A1(_09456_),
    .A2(_09252_),
    .ZN(_09470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18355_ (.A1(_09469_),
    .A2(_09470_),
    .ZN(_09471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18356_ (.A1(_09471_),
    .A2(_00401_),
    .ZN(_09472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18357_ (.A1(_09467_),
    .A2(_09187_),
    .A3(_09472_),
    .ZN(_09473_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18358_ (.A1(_09203_),
    .A2(_09189_),
    .A3(_09334_),
    .ZN(_09474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18359_ (.A1(_09474_),
    .A2(_09168_),
    .ZN(_09475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18360_ (.A1(_09378_),
    .A2(_07579_),
    .Z(_09476_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18361_ (.A1(_09475_),
    .A2(_09476_),
    .ZN(_09477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18362_ (.A1(_09254_),
    .A2(_09320_),
    .A3(_09167_),
    .ZN(_09478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18363_ (.A1(_09406_),
    .A2(_09478_),
    .A3(_09281_),
    .ZN(_09479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18364_ (.A1(_09477_),
    .A2(_09283_),
    .A3(_09479_),
    .ZN(_09480_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18365_ (.A1(_09473_),
    .A2(_09480_),
    .A3(_09211_),
    .ZN(_09481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18366_ (.A1(_09220_),
    .A2(_09183_),
    .Z(_09482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18367_ (.A1(_09465_),
    .A2(_09482_),
    .B(_09310_),
    .ZN(_09483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18368_ (.A1(_09287_),
    .A2(_09157_),
    .ZN(_09484_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18369_ (.I(_09484_),
    .ZN(_09485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18370_ (.A1(_09485_),
    .A2(_09343_),
    .ZN(_09486_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18371_ (.A1(_09346_),
    .A2(_09486_),
    .A3(_09235_),
    .ZN(_09487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18372_ (.A1(_09483_),
    .A2(_09487_),
    .B(_09237_),
    .ZN(_09488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18373_ (.A1(_09189_),
    .A2(_09333_),
    .B(_09334_),
    .ZN(_09489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18374_ (.A1(_09245_),
    .A2(_09279_),
    .B(_09205_),
    .ZN(_09490_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18375_ (.A1(_09489_),
    .A2(_09490_),
    .B(_09399_),
    .ZN(_09491_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18376_ (.A1(_09161_),
    .A2(_09174_),
    .A3(_09334_),
    .ZN(_09492_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18377_ (.A1(_09206_),
    .A2(_09492_),
    .A3(_09217_),
    .ZN(_09493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18378_ (.A1(_09491_),
    .A2(_09493_),
    .ZN(_09494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18379_ (.A1(_09494_),
    .A2(_00402_),
    .ZN(_09495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18380_ (.A1(_09488_),
    .A2(_09495_),
    .ZN(_09496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18381_ (.A1(_09481_),
    .A2(_09496_),
    .B(_09214_),
    .ZN(_09497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18382_ (.A1(_09194_),
    .A2(_09215_),
    .ZN(_09498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18383_ (.A1(_09233_),
    .A2(_09198_),
    .ZN(_09499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18384_ (.A1(_09498_),
    .A2(_09499_),
    .A3(_09226_),
    .ZN(_09500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18385_ (.A1(_09266_),
    .A2(_09252_),
    .ZN(_09501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18386_ (.A1(_09501_),
    .A2(_07586_),
    .ZN(_09502_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18387_ (.A1(_09424_),
    .A2(_09502_),
    .Z(_09503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18388_ (.A1(_09500_),
    .A2(_09503_),
    .B(_00401_),
    .ZN(_09504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18389_ (.A1(_09249_),
    .A2(_09174_),
    .B(_09205_),
    .ZN(_09505_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18390_ (.I(_09470_),
    .ZN(_09506_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18391_ (.A1(_09505_),
    .A2(_09506_),
    .B(_09186_),
    .ZN(_09507_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18392_ (.A1(_09164_),
    .A2(_09186_),
    .ZN(_09508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18393_ (.A1(_09297_),
    .A2(_07579_),
    .ZN(_09509_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18394_ (.A1(_09508_),
    .A2(_09509_),
    .ZN(_09510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18395_ (.A1(_09507_),
    .A2(_09510_),
    .ZN(_09511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18396_ (.A1(_09511_),
    .A2(_09237_),
    .ZN(_09512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18397_ (.A1(_09504_),
    .A2(_09512_),
    .B(_09214_),
    .ZN(_09513_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18398_ (.A1(_09288_),
    .A2(_09459_),
    .ZN(_09514_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18399_ (.A1(_09514_),
    .A2(_09373_),
    .B(_09399_),
    .ZN(_09515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18400_ (.A1(_09515_),
    .A2(_09426_),
    .ZN(_09516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18401_ (.A1(_09516_),
    .A2(_09187_),
    .ZN(_09517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18402_ (.A1(_09332_),
    .A2(_09303_),
    .A3(_09243_),
    .ZN(_09518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18403_ (.A1(_09194_),
    .A2(_09231_),
    .ZN(_09519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18404_ (.A1(_09215_),
    .A2(_09265_),
    .ZN(_09520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18405_ (.A1(_09520_),
    .A2(_09205_),
    .ZN(_09521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18406_ (.A1(_09519_),
    .A2(_09235_),
    .A3(_09521_),
    .ZN(_09522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18407_ (.A1(_09518_),
    .A2(_09522_),
    .A3(_09283_),
    .ZN(_09523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18408_ (.A1(_09517_),
    .A2(_09523_),
    .B(_09237_),
    .ZN(_09524_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18409_ (.A1(_09513_),
    .A2(_09524_),
    .ZN(_09525_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18410_ (.A1(_09497_),
    .A2(_09525_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18411_ (.A1(_09396_),
    .A2(_09399_),
    .ZN(_09526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18412_ (.A1(_09156_),
    .A2(_09455_),
    .B(_09526_),
    .ZN(_09527_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18413_ (.A1(_09369_),
    .A2(_09334_),
    .Z(_09528_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18414_ (.A1(_09315_),
    .A2(_09303_),
    .A3(_09528_),
    .ZN(_09529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18415_ (.A1(_09527_),
    .A2(_09529_),
    .A3(_09187_),
    .ZN(_09530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18416_ (.A1(_09379_),
    .A2(_09265_),
    .Z(_09531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18417_ (.A1(_09264_),
    .A2(_09531_),
    .B(_09226_),
    .ZN(_09532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18418_ (.A1(_09254_),
    .A2(_09163_),
    .Z(_09533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18419_ (.A1(_09533_),
    .A2(_09165_),
    .ZN(_09534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18420_ (.A1(_09534_),
    .A2(_09291_),
    .A3(_09184_),
    .ZN(_09535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18421_ (.A1(_09532_),
    .A2(_09535_),
    .B(_09213_),
    .ZN(_09536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18422_ (.A1(_09530_),
    .A2(_09536_),
    .ZN(_09537_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18423_ (.I(_09514_),
    .ZN(_09538_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18424_ (.A1(_09155_),
    .A2(_09204_),
    .Z(_09539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18425_ (.A1(_09539_),
    .A2(_09176_),
    .ZN(_09540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18426_ (.A1(_09538_),
    .A2(_09540_),
    .A3(_09207_),
    .ZN(_09541_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18427_ (.A1(_09272_),
    .A2(_09281_),
    .A3(_09206_),
    .ZN(_09542_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18428_ (.A1(_09541_),
    .A2(_09542_),
    .A3(_09257_),
    .ZN(_09543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18429_ (.A1(_09289_),
    .A2(_09249_),
    .ZN(_09544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18430_ (.A1(_09296_),
    .A2(_09544_),
    .Z(_09545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18431_ (.A1(_09163_),
    .A2(_15607_),
    .ZN(_09546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18432_ (.A1(_09379_),
    .A2(_09546_),
    .ZN(_09547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18433_ (.A1(_09547_),
    .A2(_09183_),
    .ZN(_09548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18434_ (.A1(_09548_),
    .A2(_09310_),
    .ZN(_09549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18435_ (.A1(_09545_),
    .A2(_09549_),
    .Z(_09550_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18436_ (.A1(_09543_),
    .A2(_09550_),
    .A3(_09214_),
    .ZN(_09551_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18437_ (.A1(_09537_),
    .A2(_09551_),
    .A3(_09211_),
    .ZN(_09552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18438_ (.A1(_09249_),
    .A2(_09180_),
    .A3(_09167_),
    .ZN(_09553_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18439_ (.A1(_00400_),
    .A2(_09539_),
    .B(_09553_),
    .C(_09235_),
    .ZN(_09554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18440_ (.A1(_09370_),
    .A2(_09317_),
    .A3(_09447_),
    .ZN(_09555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18441_ (.A1(_09554_),
    .A2(_09555_),
    .A3(_09187_),
    .ZN(_09556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18442_ (.A1(_07572_),
    .A2(_15637_),
    .ZN(_09557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18443_ (.A1(_09557_),
    .A2(_09182_),
    .ZN(_09558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18444_ (.A1(_15630_),
    .A2(_09242_),
    .B(_09558_),
    .ZN(_09559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18445_ (.A1(_09559_),
    .A2(_09366_),
    .ZN(_09560_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18446_ (.A1(_09239_),
    .A2(_09399_),
    .ZN(_09561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18447_ (.A1(_09561_),
    .A2(_09288_),
    .B(_09186_),
    .ZN(_09562_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18448_ (.A1(_09560_),
    .A2(_09562_),
    .B(_09213_),
    .ZN(_09563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18449_ (.A1(_09556_),
    .A2(_09563_),
    .ZN(_09564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18450_ (.A1(_09159_),
    .A2(_07579_),
    .Z(_09565_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18451_ (.A1(_09565_),
    .A2(_09359_),
    .A3(_09368_),
    .ZN(_09566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18452_ (.A1(_09200_),
    .A2(_09231_),
    .ZN(_09567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18453_ (.A1(_00400_),
    .A2(_15625_),
    .B(_09217_),
    .ZN(_09568_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18454_ (.A1(_09567_),
    .A2(_09568_),
    .B(_09310_),
    .ZN(_09569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18455_ (.A1(_09566_),
    .A2(_09569_),
    .ZN(_09570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18456_ (.A1(_09341_),
    .A2(_07579_),
    .Z(_09571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18457_ (.A1(_09571_),
    .A2(_09387_),
    .B(_09226_),
    .ZN(_09572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18458_ (.A1(_09328_),
    .A2(_09279_),
    .ZN(_09573_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18459_ (.A1(_09573_),
    .A2(_09247_),
    .A3(_09243_),
    .ZN(_09574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18460_ (.A1(_09572_),
    .A2(_09574_),
    .ZN(_09575_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18461_ (.A1(_09570_),
    .A2(_09575_),
    .A3(_09213_),
    .ZN(_09576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18462_ (.A1(_09564_),
    .A2(_09576_),
    .A3(_00403_),
    .ZN(_09577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18463_ (.A1(_09552_),
    .A2(_09577_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18464_ (.A1(_09198_),
    .A2(_07572_),
    .ZN(_09578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18465_ (.A1(_09384_),
    .A2(_09333_),
    .A3(_09578_),
    .ZN(_09579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18466_ (.A1(_09264_),
    .A2(_09232_),
    .ZN(_09580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18467_ (.A1(_09579_),
    .A2(_00402_),
    .A3(_09580_),
    .ZN(_09581_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18468_ (.A1(_09164_),
    .A2(_09419_),
    .A3(_09217_),
    .Z(_09582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18469_ (.A1(_09179_),
    .A2(_09276_),
    .ZN(_09583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18470_ (.A1(_09582_),
    .A2(_09583_),
    .ZN(_09584_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18471_ (.A1(_09546_),
    .A2(_15625_),
    .B1(_09173_),
    .B2(_09271_),
    .ZN(_09585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18472_ (.A1(_09585_),
    .A2(_09317_),
    .B(_09310_),
    .ZN(_09586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18473_ (.A1(_09584_),
    .A2(_09586_),
    .ZN(_09587_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18474_ (.A1(_09581_),
    .A2(_09587_),
    .A3(_09211_),
    .ZN(_09588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18475_ (.A1(_09347_),
    .A2(_09419_),
    .Z(_09589_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18476_ (.A1(_09175_),
    .A2(_09167_),
    .B(_09183_),
    .ZN(_09590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18477_ (.A1(_09589_),
    .A2(_09590_),
    .B(_09310_),
    .ZN(_09591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18478_ (.A1(_09228_),
    .A2(_09320_),
    .ZN(_09592_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18479_ (.A1(_09592_),
    .A2(_09247_),
    .A3(_09243_),
    .ZN(_09593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18480_ (.A1(_09591_),
    .A2(_09593_),
    .B(_09237_),
    .ZN(_09594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18481_ (.A1(_09221_),
    .A2(_09161_),
    .ZN(_09595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18482_ (.A1(_09485_),
    .A2(_09249_),
    .ZN(_09596_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18483_ (.A1(_09595_),
    .A2(_09596_),
    .A3(_00401_),
    .ZN(_09597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18484_ (.I(_09242_),
    .ZN(_09598_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18485_ (.A1(_09202_),
    .A2(_09184_),
    .A3(_09598_),
    .ZN(_09599_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18486_ (.A1(_09597_),
    .A2(_09599_),
    .A3(_00402_),
    .ZN(_09600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18487_ (.A1(_09594_),
    .A2(_09600_),
    .ZN(_09601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18488_ (.A1(_09588_),
    .A2(_09601_),
    .A3(_09214_),
    .ZN(_09602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18489_ (.A1(_09327_),
    .A2(_09333_),
    .Z(_09603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18490_ (.A1(_09603_),
    .A2(_09207_),
    .B(_09310_),
    .ZN(_09604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18491_ (.I(_09194_),
    .ZN(_09605_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18492_ (.A1(_09521_),
    .A2(_09605_),
    .A3(_09281_),
    .ZN(_09606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18493_ (.A1(_09604_),
    .A2(_09606_),
    .B(_09237_),
    .ZN(_09607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18494_ (.A1(_09233_),
    .A2(_09224_),
    .ZN(_09608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18495_ (.A1(_09241_),
    .A2(_09184_),
    .A3(_09608_),
    .ZN(_09609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18496_ (.I(_09578_),
    .ZN(_09610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18497_ (.A1(_09610_),
    .A2(_09320_),
    .ZN(_09611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18498_ (.A1(_09485_),
    .A2(_09290_),
    .ZN(_09612_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18499_ (.A1(_09611_),
    .A2(_09612_),
    .A3(_09235_),
    .ZN(_09613_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18500_ (.A1(_09609_),
    .A2(_09613_),
    .A3(_09283_),
    .ZN(_09614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18501_ (.A1(_09607_),
    .A2(_09614_),
    .B(_09213_),
    .ZN(_09615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18502_ (.A1(_09158_),
    .A2(net87),
    .ZN(_09616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18503_ (.A1(_09156_),
    .A2(_09176_),
    .B1(_09616_),
    .B2(net86),
    .ZN(_09617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18504_ (.A1(_09617_),
    .A2(_09317_),
    .ZN(_09618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18505_ (.A1(_09228_),
    .A2(_09351_),
    .ZN(_09619_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18506_ (.A1(_09619_),
    .A2(_09590_),
    .A3(_09364_),
    .ZN(_09620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18507_ (.A1(_09618_),
    .A2(_09620_),
    .A3(_00402_),
    .ZN(_09621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18508_ (.A1(_09343_),
    .A2(_07572_),
    .Z(_09622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18509_ (.A1(_09622_),
    .A2(_09180_),
    .ZN(_09623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18510_ (.A1(_09623_),
    .A2(_09184_),
    .A3(_09419_),
    .ZN(_09624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18511_ (.A1(_09388_),
    .A2(_09278_),
    .ZN(_09625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18512_ (.A1(_09449_),
    .A2(_09625_),
    .ZN(_09626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18513_ (.A1(_09624_),
    .A2(_09626_),
    .A3(_09257_),
    .ZN(_09627_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18514_ (.A1(_09621_),
    .A2(_09627_),
    .A3(_09211_),
    .ZN(_09628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18515_ (.A1(_09615_),
    .A2(_09628_),
    .ZN(_09629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18516_ (.A1(_09602_),
    .A2(_09629_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18517_ (.A1(_09200_),
    .A2(_09279_),
    .ZN(_09630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18518_ (.A1(_09454_),
    .A2(_09203_),
    .ZN(_09631_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18519_ (.A1(_09630_),
    .A2(_09631_),
    .A3(_09317_),
    .ZN(_09632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18520_ (.A1(_09454_),
    .A2(_09369_),
    .ZN(_09633_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18521_ (.A1(_09633_),
    .A2(_00401_),
    .A3(_09298_),
    .ZN(_09634_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18522_ (.A1(_09632_),
    .A2(_09634_),
    .A3(_09187_),
    .ZN(_09635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18523_ (.A1(_09388_),
    .A2(_09343_),
    .ZN(_09636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18524_ (.A1(_09221_),
    .A2(_09249_),
    .ZN(_09637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18525_ (.A1(_09636_),
    .A2(_09637_),
    .A3(_09184_),
    .ZN(_09638_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18526_ (.A1(_09403_),
    .A2(_09162_),
    .B(_09235_),
    .C(_09433_),
    .ZN(_09639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18527_ (.A1(_09638_),
    .A2(_00402_),
    .A3(_09639_),
    .ZN(_09640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18528_ (.A1(_09635_),
    .A2(_09640_),
    .A3(_00404_),
    .ZN(_09641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18529_ (.A1(_09276_),
    .A2(_09176_),
    .ZN(_09642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18530_ (.A1(_09544_),
    .A2(_09642_),
    .B(_09281_),
    .ZN(_09643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18531_ (.A1(_09398_),
    .A2(_09399_),
    .ZN(_09644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18532_ (.A1(_09644_),
    .A2(_09257_),
    .ZN(_09645_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18533_ (.A1(_09643_),
    .A2(_09645_),
    .ZN(_09646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18534_ (.A1(_09622_),
    .A2(_09231_),
    .ZN(_09647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18535_ (.A1(_09355_),
    .A2(_09647_),
    .ZN(_09648_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18536_ (.A1(_15627_),
    .A2(_09334_),
    .B(_09182_),
    .ZN(_09649_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18537_ (.I(_09649_),
    .ZN(_09650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18538_ (.A1(_09596_),
    .A2(_09650_),
    .ZN(_09651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18539_ (.A1(_09648_),
    .A2(_09651_),
    .B(_09257_),
    .ZN(_09652_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18540_ (.A1(_09646_),
    .A2(_09652_),
    .B(_09214_),
    .ZN(_09653_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18541_ (.A1(_09641_),
    .A2(_09653_),
    .A3(_09211_),
    .ZN(_09654_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18542_ (.I(_09407_),
    .ZN(_09655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18543_ (.A1(_09266_),
    .A2(_09655_),
    .B(_09167_),
    .ZN(_09656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18544_ (.A1(_09172_),
    .A2(_09271_),
    .B(_09183_),
    .ZN(_09657_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18545_ (.A1(_09656_),
    .A2(_09657_),
    .B(_09226_),
    .ZN(_09658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18546_ (.A1(_09539_),
    .A2(_00400_),
    .ZN(_09659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18547_ (.A1(net89),
    .A2(_09176_),
    .ZN(_09660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18548_ (.A1(_09659_),
    .A2(_09281_),
    .A3(_09660_),
    .ZN(_09661_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18549_ (.A1(_09658_),
    .A2(_09661_),
    .B(_09213_),
    .ZN(_09662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18550_ (.A1(_09297_),
    .A2(_09183_),
    .Z(_09663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18551_ (.A1(_09485_),
    .A2(_09254_),
    .ZN(_09664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18552_ (.A1(_07572_),
    .A2(_09244_),
    .ZN(_09665_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18553_ (.A1(_09665_),
    .A2(_15630_),
    .Z(_09666_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18554_ (.A1(_09663_),
    .A2(_09664_),
    .A3(_09666_),
    .ZN(_09667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18555_ (.A1(_09630_),
    .A2(_09521_),
    .A3(_09235_),
    .ZN(_09668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18556_ (.A1(_09667_),
    .A2(_09668_),
    .A3(_09257_),
    .ZN(_09669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18557_ (.A1(_09662_),
    .A2(_09669_),
    .B(_09211_),
    .ZN(_09670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18558_ (.A1(_09250_),
    .A2(_09333_),
    .ZN(_09671_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18559_ (.A1(_09201_),
    .A2(_09203_),
    .A3(_09205_),
    .ZN(_09672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18560_ (.A1(_09671_),
    .A2(_09672_),
    .ZN(_09673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18561_ (.A1(_09673_),
    .A2(_09317_),
    .ZN(_09674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18562_ (.A1(_09533_),
    .A2(_09203_),
    .ZN(_09675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18563_ (.A1(_09675_),
    .A2(_09207_),
    .A3(_09672_),
    .ZN(_09676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18564_ (.A1(_09674_),
    .A2(_09676_),
    .A3(_00402_),
    .ZN(_09677_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18565_ (.A1(_09229_),
    .A2(_09207_),
    .A3(_09322_),
    .ZN(_09678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18566_ (.A1(_09357_),
    .A2(_09271_),
    .ZN(_09679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18567_ (.A1(_09521_),
    .A2(_09281_),
    .A3(_09679_),
    .ZN(_09680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18568_ (.A1(_09678_),
    .A2(_09257_),
    .A3(_09680_),
    .ZN(_09681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18569_ (.A1(_09677_),
    .A2(_09681_),
    .A3(_09214_),
    .ZN(_09682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18570_ (.A1(_09670_),
    .A2(_09682_),
    .ZN(_09683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18571_ (.A1(_09654_),
    .A2(_09683_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18572_ (.A1(_09176_),
    .A2(_09655_),
    .B(_09172_),
    .ZN(_09684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18573_ (.A1(_09156_),
    .A2(_00400_),
    .ZN(_09685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18574_ (.A1(_09684_),
    .A2(_09317_),
    .A3(_09685_),
    .ZN(_09686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18575_ (.A1(_09176_),
    .A2(_15614_),
    .ZN(_09687_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18576_ (.A1(_09659_),
    .A2(_00401_),
    .A3(_09687_),
    .ZN(_09688_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18577_ (.A1(_09686_),
    .A2(_09688_),
    .A3(_09187_),
    .ZN(_09689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18578_ (.A1(_09319_),
    .A2(_09195_),
    .ZN(_09690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18579_ (.A1(_09538_),
    .A2(_09690_),
    .A3(_09207_),
    .ZN(_09691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18580_ (.A1(_09343_),
    .A2(_09276_),
    .A3(_00400_),
    .ZN(_09692_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18581_ (.A1(_09205_),
    .A2(_15607_),
    .A3(_15630_),
    .Z(_09693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18582_ (.A1(_09443_),
    .A2(_09692_),
    .A3(_09693_),
    .ZN(_09694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18583_ (.A1(_09691_),
    .A2(_09694_),
    .A3(_09283_),
    .ZN(_09695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18584_ (.A1(_09689_),
    .A2(_09695_),
    .A3(_00403_),
    .ZN(_09696_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18585_ (.I(_09267_),
    .ZN(_09697_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18586_ (.A1(_09697_),
    .A2(_09558_),
    .ZN(_09698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18587_ (.A1(_09456_),
    .A2(_09176_),
    .ZN(_09699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18588_ (.A1(_09698_),
    .A2(_09699_),
    .B(_09310_),
    .ZN(_09700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18589_ (.A1(_09622_),
    .A2(_09165_),
    .ZN(_09701_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18590_ (.A1(_09355_),
    .A2(_09701_),
    .A3(_09457_),
    .ZN(_09702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18591_ (.A1(_09700_),
    .A2(_09702_),
    .ZN(_09703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18592_ (.A1(_09565_),
    .A2(_09295_),
    .A3(_09368_),
    .ZN(_09704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18593_ (.A1(_09665_),
    .A2(_09183_),
    .ZN(_09705_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18594_ (.I(_09705_),
    .ZN(_09706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18595_ (.A1(_09655_),
    .A2(_09176_),
    .ZN(_09707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18596_ (.A1(_09706_),
    .A2(_09707_),
    .B(_09186_),
    .ZN(_09708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18597_ (.A1(_09704_),
    .A2(_09708_),
    .ZN(_09709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18598_ (.A1(_09703_),
    .A2(_09211_),
    .A3(_09709_),
    .ZN(_09710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18599_ (.A1(_09696_),
    .A2(_09710_),
    .A3(_00404_),
    .ZN(_09711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18600_ (.A1(_09216_),
    .A2(_09290_),
    .ZN(_09712_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18601_ (.A1(_09476_),
    .A2(_09666_),
    .A3(_09712_),
    .ZN(_09713_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18602_ (.A1(_09533_),
    .A2(_09217_),
    .ZN(_09714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18603_ (.A1(_09714_),
    .A2(_09544_),
    .B(_09226_),
    .ZN(_09715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18604_ (.A1(_09713_),
    .A2(_09715_),
    .B(_09237_),
    .ZN(_09716_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18605_ (.A1(_09460_),
    .A2(_09664_),
    .A3(_09184_),
    .ZN(_09717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18606_ (.A1(_09498_),
    .A2(_09207_),
    .A3(_09316_),
    .ZN(_09718_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18607_ (.A1(_09717_),
    .A2(_09718_),
    .A3(_09187_),
    .ZN(_09719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18608_ (.A1(_09716_),
    .A2(_09719_),
    .ZN(_09720_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18609_ (.A1(_09343_),
    .A2(_09195_),
    .A3(_09271_),
    .ZN(_09721_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18610_ (.A1(_09455_),
    .A2(_09721_),
    .A3(_09235_),
    .ZN(_09722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18611_ (.A1(_09247_),
    .A2(_09164_),
    .ZN(_09723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18612_ (.A1(_09722_),
    .A2(_09723_),
    .A3(_09257_),
    .ZN(_09724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18613_ (.A1(_09610_),
    .A2(_09155_),
    .ZN(_09725_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18614_ (.A1(_09616_),
    .A2(_07579_),
    .Z(_09726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18615_ (.A1(_09725_),
    .A2(_09726_),
    .B(_09226_),
    .ZN(_09727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18616_ (.A1(_09250_),
    .A2(_09195_),
    .ZN(_09728_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18617_ (.A1(_09728_),
    .A2(_09281_),
    .A3(_09447_),
    .ZN(_09729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18618_ (.A1(_09727_),
    .A2(_09729_),
    .ZN(_09730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18619_ (.A1(_09724_),
    .A2(_09730_),
    .A3(_09211_),
    .ZN(_09731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18620_ (.A1(_09720_),
    .A2(_09731_),
    .A3(_09214_),
    .ZN(_09732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18621_ (.A1(_09711_),
    .A2(_09732_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _18622_ (.I(_15650_),
    .ZN(_15639_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18623_ (.A1(_07437_),
    .A2(net134),
    .ZN(_09733_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18624_ (.A1(_07437_),
    .A2(_07694_),
    .B(_09733_),
    .ZN(_09734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _18625_ (.I(_09734_),
    .Z(_15659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18626_ (.A1(_07404_),
    .A2(_07679_),
    .ZN(_09735_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18627_ (.I(_07680_),
    .ZN(_09736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18628_ (.A1(_09735_),
    .A2(_09736_),
    .ZN(_15640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18629_ (.A1(net825),
    .A2(net706),
    .ZN(_09737_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18630_ (.I(_09737_),
    .ZN(_09738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18631_ (.A1(_09738_),
    .A2(net25),
    .Z(_09739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18632_ (.I(_15641_),
    .ZN(_09740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18633_ (.A1(net832),
    .A2(_09740_),
    .ZN(_09741_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _18634_ (.I(_07706_),
    .ZN(_09742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18635_ (.A1(_09741_),
    .A2(_09742_),
    .B(_07716_),
    .ZN(_09743_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18636_ (.A1(_09739_),
    .A2(_09743_),
    .ZN(_09744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18637_ (.I(_09744_),
    .ZN(_09745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18638_ (.A1(_15659_),
    .A2(_15653_),
    .ZN(_09746_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18639_ (.I(_09746_),
    .ZN(_09747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18640_ (.I(_09742_),
    .Z(_09748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18641_ (.A1(_09747_),
    .A2(_09748_),
    .ZN(_09749_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18642_ (.I(_07717_),
    .Z(_09750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18643_ (.I(_15642_),
    .ZN(_09751_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18644_ (.A1(_07695_),
    .A2(_09751_),
    .A3(_07696_),
    .ZN(_09752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18645_ (.A1(_09752_),
    .A2(net824),
    .ZN(_09753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18646_ (.A1(_09749_),
    .A2(_09750_),
    .A3(_09753_),
    .ZN(_09754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18647_ (.A1(_09745_),
    .A2(_09754_),
    .ZN(_09755_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _18648_ (.I(_07697_),
    .Z(_09756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18649_ (.A1(_09756_),
    .A2(_15648_),
    .ZN(_09757_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18650_ (.I(_09757_),
    .ZN(_09758_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18651_ (.I(_09742_),
    .Z(_09759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18652_ (.A1(_09758_),
    .A2(_09759_),
    .ZN(_09760_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18653_ (.A1(_09760_),
    .A2(_07726_),
    .Z(_09761_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18654_ (.I(_07735_),
    .ZN(_09762_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18655_ (.I(_09762_),
    .Z(_09763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18656_ (.A1(_09755_),
    .A2(_09761_),
    .B(_09763_),
    .ZN(_09764_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18657_ (.I(_15655_),
    .ZN(_09765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18658_ (.A1(_09756_),
    .A2(_09765_),
    .ZN(_09766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18659_ (.I(_09766_),
    .ZN(_09767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18660_ (.A1(_15659_),
    .A2(_15657_),
    .Z(_09768_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18661_ (.I(_09742_),
    .Z(_09769_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18662_ (.A1(_09767_),
    .A2(_09768_),
    .B(_09769_),
    .ZN(_09770_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18663_ (.I(_15648_),
    .ZN(_09771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18664_ (.A1(_09771_),
    .A2(_15659_),
    .ZN(_09772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18665_ (.I(_07706_),
    .Z(_09773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18666_ (.A1(_09772_),
    .A2(_09773_),
    .ZN(_09774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18667_ (.A1(_09770_),
    .A2(_09774_),
    .ZN(_09775_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18668_ (.I(_07717_),
    .Z(_09776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18669_ (.A1(_09775_),
    .A2(_09776_),
    .ZN(_09777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18670_ (.A1(net37),
    .A2(_15659_),
    .ZN(_09778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18671_ (.A1(net707),
    .A2(net711),
    .ZN(_09779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18672_ (.A1(_09778_),
    .A2(_09779_),
    .A3(_09759_),
    .ZN(_09780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18673_ (.I(_09780_),
    .ZN(_09781_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18674_ (.I(_15651_),
    .ZN(_09782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18675_ (.A1(_09756_),
    .A2(_09782_),
    .ZN(_09783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18676_ (.A1(net838),
    .A2(_15640_),
    .ZN(_09784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18677_ (.A1(_09783_),
    .A2(_09784_),
    .B(_09748_),
    .ZN(_09785_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18678_ (.I(_07716_),
    .Z(_09786_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18679_ (.I(_09786_),
    .Z(_09787_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18680_ (.A1(_09781_),
    .A2(_09785_),
    .B(_09787_),
    .ZN(_09788_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18681_ (.I(_07727_),
    .Z(_09789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18682_ (.A1(_09777_),
    .A2(_09788_),
    .A3(_09789_),
    .ZN(_09790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18683_ (.A1(_09764_),
    .A2(_09790_),
    .ZN(_09791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18684_ (.I(_15653_),
    .ZN(_09792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18685_ (.A1(_09792_),
    .A2(_09756_),
    .ZN(_09793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18686_ (.A1(_15659_),
    .A2(_15646_),
    .ZN(_09794_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18687_ (.I(_09773_),
    .Z(_09795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18688_ (.A1(_09793_),
    .A2(_09794_),
    .A3(_09795_),
    .ZN(_09796_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18689_ (.I(_09786_),
    .Z(_09797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18690_ (.A1(_09768_),
    .A2(_09759_),
    .ZN(_09798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18691_ (.A1(_09796_),
    .A2(_09797_),
    .A3(_09798_),
    .ZN(_09799_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18692_ (.I(_09783_),
    .ZN(_09800_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18693_ (.I(_15646_),
    .ZN(_09801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18694_ (.A1(_15659_),
    .A2(_09801_),
    .ZN(_09802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18695_ (.I(_09802_),
    .ZN(_09803_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18696_ (.A1(_09800_),
    .A2(_09803_),
    .B(_09748_),
    .ZN(_09804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18697_ (.A1(_09768_),
    .A2(_09795_),
    .B(_09786_),
    .ZN(_09805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18698_ (.A1(_09804_),
    .A2(_09805_),
    .ZN(_09806_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18699_ (.I(_07727_),
    .Z(_09807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18700_ (.A1(_09799_),
    .A2(_09806_),
    .A3(_09807_),
    .ZN(_09808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18701_ (.A1(_09765_),
    .A2(net833),
    .ZN(_09809_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18702_ (.I(_09742_),
    .Z(_09810_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18703_ (.A1(_09809_),
    .A2(_09810_),
    .B(_09786_),
    .ZN(_09811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18704_ (.A1(_09739_),
    .A2(_09811_),
    .ZN(_09812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18705_ (.A1(_09756_),
    .A2(net25),
    .ZN(_09813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18706_ (.A1(_09813_),
    .A2(_09742_),
    .Z(_09814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18707_ (.A1(_09814_),
    .A2(_09794_),
    .ZN(_09815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18708_ (.A1(_09812_),
    .A2(_09815_),
    .ZN(_09816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18709_ (.I(_09779_),
    .ZN(_09817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18710_ (.A1(_09817_),
    .A2(_09748_),
    .ZN(_09818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18711_ (.A1(_09795_),
    .A2(_15662_),
    .B(_09786_),
    .ZN(_09819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18712_ (.A1(_09818_),
    .A2(_09819_),
    .B(_07727_),
    .ZN(_09820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18713_ (.A1(_09816_),
    .A2(_09820_),
    .ZN(_09821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18714_ (.A1(_09808_),
    .A2(_09821_),
    .ZN(_09822_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18715_ (.I(_09762_),
    .Z(_09823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18716_ (.A1(_09822_),
    .A2(_09823_),
    .ZN(_09824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18717_ (.A1(_09791_),
    .A2(_09824_),
    .ZN(_09825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18718_ (.A1(_09825_),
    .A2(_00399_),
    .ZN(_09826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18719_ (.A1(_09756_),
    .A2(net759),
    .ZN(_09827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18720_ (.A1(_09827_),
    .A2(_09810_),
    .Z(_09828_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18721_ (.I(_07717_),
    .Z(_09829_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18722_ (.A1(_09828_),
    .A2(_09829_),
    .ZN(_09830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18723_ (.A1(_09756_),
    .A2(_15646_),
    .ZN(_09831_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18724_ (.I(_09773_),
    .Z(_09832_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18725_ (.A1(_09831_),
    .A2(_09772_),
    .A3(_09832_),
    .ZN(_09833_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18726_ (.I(_07726_),
    .Z(_09834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18727_ (.A1(_09830_),
    .A2(_09833_),
    .B(_09834_),
    .ZN(_09835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18728_ (.A1(_09831_),
    .A2(_09810_),
    .ZN(_09836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18729_ (.I(_09836_),
    .ZN(_09837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18730_ (.A1(net832),
    .A2(net962),
    .ZN(_09838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18731_ (.A1(_09837_),
    .A2(_09838_),
    .ZN(_09839_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _18732_ (.I(_09753_),
    .ZN(_09840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18733_ (.I(_15643_),
    .ZN(_09841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18734_ (.A1(_09841_),
    .A2(_09756_),
    .ZN(_09842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18735_ (.A1(_09840_),
    .A2(_09842_),
    .ZN(_09843_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18736_ (.I(_09750_),
    .Z(_09844_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18737_ (.A1(_09839_),
    .A2(_09843_),
    .A3(_09844_),
    .ZN(_09845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18738_ (.A1(_09835_),
    .A2(_09845_),
    .B(_09763_),
    .ZN(_09846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18739_ (.A1(net832),
    .A2(net11),
    .ZN(_09847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18740_ (.A1(_09837_),
    .A2(_09847_),
    .ZN(_09848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18741_ (.A1(_09841_),
    .A2(net839),
    .ZN(_09849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18742_ (.A1(_09849_),
    .A2(_09773_),
    .ZN(_09850_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18743_ (.I(_09850_),
    .ZN(_09851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18744_ (.A1(_09851_),
    .A2(_09827_),
    .ZN(_09852_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18745_ (.A1(_09848_),
    .A2(_09852_),
    .A3(_09844_),
    .ZN(_09853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18746_ (.A1(net706),
    .A2(net481),
    .ZN(_09854_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18747_ (.I(_09854_),
    .ZN(_09855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18748_ (.A1(_09855_),
    .A2(_09759_),
    .ZN(_09856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18749_ (.A1(_09856_),
    .A2(_09798_),
    .Z(_09857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18750_ (.A1(_09744_),
    .A2(_09857_),
    .ZN(_09858_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18751_ (.I(_07726_),
    .Z(_09859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18752_ (.A1(_09853_),
    .A2(_09858_),
    .A3(_09859_),
    .ZN(_09860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18753_ (.A1(_09846_),
    .A2(_09860_),
    .B(_00399_),
    .ZN(_09861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18754_ (.A1(_09856_),
    .A2(_09750_),
    .ZN(_09862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18755_ (.A1(_09756_),
    .A2(_09751_),
    .ZN(_09863_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18756_ (.A1(_09863_),
    .A2(_09773_),
    .Z(_09864_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18757_ (.A1(_09752_),
    .A2(_07707_),
    .ZN(_09865_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18758_ (.A1(_09862_),
    .A2(_09864_),
    .A3(_09865_),
    .ZN(_09866_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _18759_ (.I(_09809_),
    .ZN(_09867_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18760_ (.I(_09810_),
    .Z(_09868_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18761_ (.A1(_09800_),
    .A2(_09867_),
    .B(_09868_),
    .ZN(_09869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18762_ (.A1(_15664_),
    .A2(_15655_),
    .ZN(_09870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18763_ (.A1(_09840_),
    .A2(_09870_),
    .ZN(_09871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18764_ (.A1(_09869_),
    .A2(_09871_),
    .B(_09776_),
    .ZN(_09872_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18765_ (.A1(_09866_),
    .A2(_09872_),
    .B(_09859_),
    .ZN(_09873_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18766_ (.A1(_09784_),
    .A2(_09742_),
    .Z(_09874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18767_ (.A1(net757),
    .A2(net11),
    .ZN(_09875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18768_ (.A1(_09874_),
    .A2(_09875_),
    .ZN(_09876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18769_ (.I(_09784_),
    .ZN(_09877_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18770_ (.I(_09875_),
    .ZN(_09878_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18771_ (.I(_09773_),
    .Z(_09879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18772_ (.A1(_09877_),
    .A2(_09878_),
    .B(_09879_),
    .ZN(_09880_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18773_ (.A1(_09876_),
    .A2(_09880_),
    .A3(_09844_),
    .ZN(_09881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18774_ (.A1(_09767_),
    .A2(_09832_),
    .B(_09750_),
    .ZN(_09882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18775_ (.A1(_09742_),
    .A2(_09752_),
    .ZN(_09883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18776_ (.I(_09883_),
    .ZN(_09884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18777_ (.A1(_09756_),
    .A2(_15641_),
    .ZN(_09885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18778_ (.A1(_09884_),
    .A2(_09885_),
    .ZN(_09886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18779_ (.A1(_15659_),
    .A2(_09782_),
    .Z(_09887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18780_ (.A1(_09887_),
    .A2(_09795_),
    .ZN(_09888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18781_ (.A1(_09882_),
    .A2(_09886_),
    .A3(_09888_),
    .ZN(_09889_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18782_ (.A1(_09881_),
    .A2(_09889_),
    .A3(_00397_),
    .ZN(_09890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18783_ (.A1(_09873_),
    .A2(_09890_),
    .A3(_09823_),
    .ZN(_09891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18784_ (.A1(_09861_),
    .A2(_09891_),
    .ZN(_09892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18785_ (.A1(_09826_),
    .A2(_09892_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18786_ (.A1(_09774_),
    .A2(_09855_),
    .Z(_09893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18787_ (.A1(_09874_),
    .A2(_09870_),
    .ZN(_09894_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18788_ (.I(_09786_),
    .Z(_09895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18789_ (.A1(_09893_),
    .A2(_09894_),
    .A3(_09895_),
    .ZN(_09896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18790_ (.A1(net761),
    .A2(_09748_),
    .B(_09750_),
    .ZN(_09897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18791_ (.I(_09798_),
    .ZN(_09898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18792_ (.A1(_09897_),
    .A2(_09898_),
    .ZN(_09899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18793_ (.I(_09813_),
    .ZN(_09900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18794_ (.A1(_09900_),
    .A2(_09810_),
    .ZN(_09901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18795_ (.A1(_09817_),
    .A2(_09795_),
    .ZN(_09902_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18796_ (.A1(_09901_),
    .A2(_09902_),
    .Z(_09903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18797_ (.A1(_09899_),
    .A2(_09903_),
    .ZN(_09904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18798_ (.A1(_09896_),
    .A2(_09904_),
    .A3(_00397_),
    .ZN(_09905_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18799_ (.A1(_09741_),
    .A2(_09773_),
    .Z(_09906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18800_ (.A1(_09906_),
    .A2(_09901_),
    .Z(_09907_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18801_ (.I(_07716_),
    .Z(_09908_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18802_ (.A1(net760),
    .A2(_09908_),
    .Z(_09909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18803_ (.A1(_09909_),
    .A2(_09907_),
    .B(_09807_),
    .ZN(_09910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18804_ (.A1(_09885_),
    .A2(_07707_),
    .Z(_09911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18805_ (.A1(net832),
    .A2(net711),
    .ZN(_09912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18806_ (.A1(_09911_),
    .A2(net823),
    .ZN(_09913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18807_ (.A1(_09849_),
    .A2(_09810_),
    .ZN(_09914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18808_ (.I(_09914_),
    .ZN(_09915_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18809_ (.I(_15657_),
    .ZN(_09916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18810_ (.A1(_15664_),
    .A2(_09916_),
    .ZN(_09917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18811_ (.A1(_09915_),
    .A2(_09917_),
    .ZN(_09918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18812_ (.A1(_09913_),
    .A2(_09918_),
    .A3(_00396_),
    .ZN(_09919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18813_ (.A1(_09910_),
    .A2(_09919_),
    .ZN(_09920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18814_ (.A1(_09905_),
    .A2(_09920_),
    .A3(_00398_),
    .ZN(_09921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18815_ (.A1(_09870_),
    .A2(_09838_),
    .A3(_09759_),
    .ZN(_09922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18816_ (.A1(_15659_),
    .A2(_15641_),
    .ZN(_09923_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18817_ (.I(_07707_),
    .Z(_09924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18818_ (.A1(_09831_),
    .A2(_09923_),
    .A3(_09924_),
    .ZN(_09925_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18819_ (.A1(_09922_),
    .A2(_09925_),
    .A3(_09807_),
    .ZN(_09926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18820_ (.A1(_09926_),
    .A2(_00396_),
    .ZN(_09927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18821_ (.A1(_15664_),
    .A2(net37),
    .ZN(_09928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18822_ (.A1(_09874_),
    .A2(_09928_),
    .ZN(_09929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18823_ (.A1(_09893_),
    .A2(_09929_),
    .ZN(_09930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18824_ (.A1(_09930_),
    .A2(_09789_),
    .ZN(_09931_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18825_ (.A1(_09748_),
    .A2(_15669_),
    .A3(_07727_),
    .Z(_09932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18826_ (.A1(_09783_),
    .A2(_09741_),
    .ZN(_09933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18827_ (.A1(_09933_),
    .A2(_09769_),
    .ZN(_09934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18828_ (.A1(_09932_),
    .A2(_09934_),
    .ZN(_09935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18829_ (.A1(_09935_),
    .A2(_09895_),
    .ZN(_09936_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18830_ (.A1(_09927_),
    .A2(_09931_),
    .B(_09823_),
    .C(_09936_),
    .ZN(_09937_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18831_ (.I(_07744_),
    .Z(_09938_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18832_ (.A1(_09921_),
    .A2(_09937_),
    .A3(_09938_),
    .ZN(_09939_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18833_ (.I(_09810_),
    .Z(_09940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18834_ (.A1(_09758_),
    .A2(_09940_),
    .B(_09908_),
    .ZN(_09941_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18835_ (.I(_09847_),
    .ZN(_09942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18836_ (.A1(_07704_),
    .A2(_07705_),
    .B(_15665_),
    .ZN(_09943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18837_ (.A1(_09942_),
    .A2(_09868_),
    .B(_09943_),
    .ZN(_09944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18838_ (.A1(_09941_),
    .A2(_09944_),
    .B(_09807_),
    .ZN(_09945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18839_ (.A1(_09851_),
    .A2(_09863_),
    .ZN(_09946_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _18840_ (.I(_09786_),
    .Z(_09947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18841_ (.A1(_09757_),
    .A2(_09802_),
    .ZN(_09948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18842_ (.A1(_09948_),
    .A2(_09940_),
    .ZN(_09949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18843_ (.A1(_09946_),
    .A2(_09947_),
    .A3(_09949_),
    .ZN(_09950_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18844_ (.I(_07735_),
    .Z(_09951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18845_ (.A1(_09945_),
    .A2(_09950_),
    .B(_09951_),
    .ZN(_09952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18846_ (.A1(_09772_),
    .A2(_09759_),
    .ZN(_09953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18847_ (.I(_09953_),
    .ZN(_09954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18848_ (.A1(_09954_),
    .A2(_09813_),
    .ZN(_09955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18849_ (.A1(_09840_),
    .A2(_09827_),
    .ZN(_09956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18850_ (.A1(_09955_),
    .A2(_09956_),
    .A3(_09844_),
    .ZN(_09957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18851_ (.A1(_09778_),
    .A2(_09940_),
    .A3(_09875_),
    .ZN(_09958_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18852_ (.A1(_15664_),
    .A2(_09801_),
    .Z(_09959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18853_ (.A1(_09959_),
    .A2(_09795_),
    .ZN(_09960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18854_ (.A1(_09958_),
    .A2(_09960_),
    .A3(_09947_),
    .ZN(_09961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18855_ (.A1(_09957_),
    .A2(_00397_),
    .A3(_09961_),
    .ZN(_09962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18856_ (.A1(_09952_),
    .A2(_09962_),
    .B(_09938_),
    .ZN(_09963_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18857_ (.A1(_09779_),
    .A2(_09838_),
    .A3(_09769_),
    .Z(_09964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18858_ (.A1(net37),
    .A2(net25),
    .ZN(_09965_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18859_ (.A1(_09965_),
    .A2(_09838_),
    .B(_09748_),
    .ZN(_09966_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18860_ (.A1(_09964_),
    .A2(_09966_),
    .B(_09787_),
    .ZN(_09967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18861_ (.A1(_09814_),
    .A2(_09809_),
    .ZN(_09968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18862_ (.A1(_09840_),
    .A2(_09757_),
    .ZN(_09969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18863_ (.A1(_09968_),
    .A2(_09969_),
    .A3(_09829_),
    .ZN(_09970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18864_ (.A1(_09967_),
    .A2(_09970_),
    .ZN(_09971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18865_ (.A1(_09971_),
    .A2(_09859_),
    .ZN(_09972_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18866_ (.A1(_09842_),
    .A2(_07707_),
    .Z(_09973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18867_ (.A1(_09973_),
    .A2(_09847_),
    .ZN(_09974_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18868_ (.A1(_09974_),
    .A2(_00396_),
    .A3(_09906_),
    .ZN(_09975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18869_ (.A1(_09759_),
    .A2(_15648_),
    .ZN(_09976_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18870_ (.A1(_09976_),
    .A2(_15664_),
    .Z(_09977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18871_ (.A1(_09913_),
    .A2(_09947_),
    .A3(_09977_),
    .ZN(_09978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18872_ (.A1(_09975_),
    .A2(_09978_),
    .A3(_09789_),
    .ZN(_09979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18873_ (.A1(_09972_),
    .A2(_09979_),
    .A3(_00398_),
    .ZN(_09980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18874_ (.A1(_09963_),
    .A2(_09980_),
    .ZN(_09981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18875_ (.A1(_09939_),
    .A2(_09981_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18876_ (.A1(_09757_),
    .A2(_09802_),
    .A3(_09879_),
    .ZN(_09982_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18877_ (.A1(_09780_),
    .A2(_09982_),
    .A3(_09787_),
    .Z(_09983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18878_ (.A1(_09778_),
    .A2(_09831_),
    .A3(_07707_),
    .ZN(_09984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18879_ (.A1(_09842_),
    .A2(_09772_),
    .A3(_09940_),
    .ZN(_09985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18880_ (.A1(_09984_),
    .A2(_09985_),
    .B(_09947_),
    .ZN(_09986_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18881_ (.A1(_09983_),
    .A2(_09986_),
    .B(_09823_),
    .ZN(_09987_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _18882_ (.I(_09759_),
    .Z(_09988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18883_ (.A1(_09747_),
    .A2(_09988_),
    .B(_09797_),
    .ZN(_09989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18884_ (.A1(_15664_),
    .A2(_09771_),
    .ZN(_09990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18885_ (.A1(_09990_),
    .A2(_09838_),
    .A3(_00395_),
    .ZN(_09991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18886_ (.A1(_15664_),
    .A2(_15643_),
    .ZN(_09992_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18887_ (.A1(_09992_),
    .A2(_09832_),
    .Z(_09993_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18888_ (.A1(_09989_),
    .A2(_09991_),
    .A3(_09993_),
    .ZN(_09994_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18889_ (.A1(_09746_),
    .A2(_09879_),
    .B(_09786_),
    .ZN(_09995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18890_ (.I(_09995_),
    .ZN(_09996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18891_ (.A1(_09990_),
    .A2(_09847_),
    .A3(_09832_),
    .ZN(_09997_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18892_ (.A1(_09996_),
    .A2(_09760_),
    .A3(_09997_),
    .ZN(_09998_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18893_ (.A1(_09994_),
    .A2(_09998_),
    .A3(_00398_),
    .ZN(_09999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18894_ (.A1(_09987_),
    .A2(_09999_),
    .A3(_09859_),
    .ZN(_10000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18895_ (.A1(_09992_),
    .A2(_09769_),
    .ZN(_10001_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18896_ (.A1(_10001_),
    .A2(_09877_),
    .B(_09829_),
    .ZN(_10002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18897_ (.A1(_09854_),
    .A2(_09746_),
    .A3(_09879_),
    .Z(_10003_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18898_ (.A1(_10002_),
    .A2(_10003_),
    .ZN(_10004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18899_ (.A1(_09793_),
    .A2(_09838_),
    .A3(_09940_),
    .ZN(_10005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18900_ (.A1(net765),
    .A2(net624),
    .A3(_09832_),
    .ZN(_10006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18901_ (.A1(_10005_),
    .A2(_10006_),
    .B(_09776_),
    .ZN(_10007_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18902_ (.A1(_10004_),
    .A2(_10007_),
    .B(_00398_),
    .ZN(_10008_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18903_ (.A1(_09836_),
    .A2(_09908_),
    .Z(_10009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18904_ (.A1(_09911_),
    .A2(_09849_),
    .ZN(_10010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18905_ (.A1(_10009_),
    .A2(_10010_),
    .B(_09951_),
    .ZN(_10011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18906_ (.A1(_15664_),
    .A2(_15657_),
    .ZN(_10012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18907_ (.I(_10012_),
    .ZN(_10013_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18908_ (.A1(_10013_),
    .A2(_09877_),
    .B(_09924_),
    .ZN(_10014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18909_ (.A1(_09928_),
    .A2(_09988_),
    .A3(net624),
    .ZN(_10015_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18910_ (.A1(_10014_),
    .A2(_00396_),
    .A3(_10015_),
    .ZN(_10016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18911_ (.A1(_10011_),
    .A2(_10016_),
    .ZN(_10017_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18912_ (.A1(_10008_),
    .A2(_00397_),
    .A3(_10017_),
    .ZN(_10018_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18913_ (.A1(_10000_),
    .A2(_10018_),
    .A3(_09938_),
    .ZN(_10019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18914_ (.A1(_09867_),
    .A2(_09748_),
    .B(_07717_),
    .ZN(_10020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18915_ (.A1(_09840_),
    .A2(_09990_),
    .ZN(_10021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18916_ (.A1(_10021_),
    .A2(_10020_),
    .B(_07726_),
    .ZN(_10022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18917_ (.A1(_09784_),
    .A2(_09773_),
    .Z(_10023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18918_ (.A1(_10023_),
    .A2(_09885_),
    .ZN(_10024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18919_ (.A1(_10024_),
    .A2(_09750_),
    .A3(_09934_),
    .ZN(_10025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18920_ (.A1(_10025_),
    .A2(_10022_),
    .ZN(_10026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18921_ (.A1(_09810_),
    .A2(_15667_),
    .ZN(_10027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18922_ (.A1(_10027_),
    .A2(_07717_),
    .ZN(_10028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18923_ (.I(_10028_),
    .ZN(_10029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18924_ (.A1(_10029_),
    .A2(_09984_),
    .ZN(_10030_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18925_ (.A1(_09810_),
    .A2(_15660_),
    .Z(_10031_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18926_ (.A1(_09908_),
    .A2(_09836_),
    .A3(_10031_),
    .ZN(_10032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18927_ (.A1(_10030_),
    .A2(_10032_),
    .A3(_07726_),
    .ZN(_10033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18928_ (.A1(_10033_),
    .A2(_09763_),
    .A3(_10026_),
    .ZN(_10034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18929_ (.A1(_00399_),
    .A2(_10034_),
    .ZN(_10035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18930_ (.I(_10035_),
    .ZN(_10036_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18931_ (.A1(_09817_),
    .A2(_09887_),
    .B(_09924_),
    .ZN(_10037_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18932_ (.A1(_09870_),
    .A2(_09847_),
    .A3(_09868_),
    .ZN(_10038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18933_ (.A1(_10037_),
    .A2(_10038_),
    .B(_09947_),
    .ZN(_10039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18934_ (.A1(_09778_),
    .A2(_07707_),
    .A3(_09875_),
    .ZN(_10040_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18935_ (.A1(_09879_),
    .A2(_15669_),
    .Z(_10041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18936_ (.A1(_10040_),
    .A2(_10041_),
    .B(_09776_),
    .ZN(_10042_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18937_ (.A1(_10039_),
    .A2(_10042_),
    .B(_09859_),
    .ZN(_10043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18938_ (.A1(_09854_),
    .A2(_09838_),
    .A3(_09832_),
    .ZN(_10044_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18939_ (.A1(_09780_),
    .A2(_10044_),
    .A3(_09844_),
    .ZN(_10045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18940_ (.A1(_09794_),
    .A2(_09773_),
    .ZN(_10046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18941_ (.I(_09863_),
    .ZN(_10047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18942_ (.A1(_09940_),
    .A2(_15662_),
    .ZN(_10048_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18943_ (.A1(_10046_),
    .A2(_10047_),
    .B(_10048_),
    .C(_09787_),
    .ZN(_10049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18944_ (.A1(_10045_),
    .A2(_10049_),
    .A3(_09789_),
    .ZN(_10050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18945_ (.A1(_10043_),
    .A2(_00398_),
    .A3(_10050_),
    .ZN(_10051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18946_ (.A1(_10036_),
    .A2(_10051_),
    .ZN(_10052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18947_ (.A1(_10052_),
    .A2(_10019_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18948_ (.A1(_09851_),
    .A2(_09990_),
    .Z(_10053_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18949_ (.A1(_09854_),
    .A2(net822),
    .A3(_09769_),
    .Z(_10054_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18950_ (.A1(_10053_),
    .A2(_10054_),
    .B(_09787_),
    .ZN(_10055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18951_ (.I(_09887_),
    .ZN(_10056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18952_ (.A1(_09814_),
    .A2(_10056_),
    .ZN(_10057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18953_ (.A1(_09864_),
    .A2(net761),
    .ZN(_10058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18954_ (.A1(_10057_),
    .A2(_10058_),
    .A3(_09776_),
    .ZN(_10059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18955_ (.A1(_10055_),
    .A2(_10059_),
    .A3(_09763_),
    .ZN(_10060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18956_ (.A1(_09923_),
    .A2(_09810_),
    .ZN(_10061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18957_ (.I(_10061_),
    .ZN(_10062_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18958_ (.A1(_10062_),
    .A2(_09863_),
    .Z(_10063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18959_ (.A1(_09960_),
    .A2(_09888_),
    .ZN(_10064_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18960_ (.A1(_10063_),
    .A2(_10064_),
    .B(_09787_),
    .ZN(_10065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18961_ (.A1(_09884_),
    .A2(_09783_),
    .ZN(_10066_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18962_ (.A1(_09880_),
    .A2(_10066_),
    .A3(_09829_),
    .ZN(_10067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18963_ (.A1(_10065_),
    .A2(_10067_),
    .A3(_09951_),
    .ZN(_10068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18964_ (.A1(_10060_),
    .A2(_10068_),
    .ZN(_10069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18965_ (.A1(_10069_),
    .A2(_00397_),
    .ZN(_10070_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18966_ (.A1(_09900_),
    .A2(_09878_),
    .B(_09940_),
    .ZN(_10071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18967_ (.A1(_09840_),
    .A2(_09854_),
    .ZN(_10072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18968_ (.A1(_10071_),
    .A2(_10072_),
    .A3(_09895_),
    .ZN(_10073_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18969_ (.A1(_09863_),
    .A2(_09924_),
    .B(_09797_),
    .ZN(_10074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18970_ (.A1(_09854_),
    .A2(_09838_),
    .A3(_09868_),
    .ZN(_10075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18971_ (.A1(_10074_),
    .A2(_10075_),
    .B(_07735_),
    .ZN(_10076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18972_ (.A1(_10073_),
    .A2(_10076_),
    .B(_09789_),
    .ZN(_10077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18973_ (.A1(_09793_),
    .A2(_09769_),
    .Z(_10078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18974_ (.A1(_10078_),
    .A2(net823),
    .ZN(_10079_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18975_ (.A1(_09974_),
    .A2(_10079_),
    .A3(_00396_),
    .ZN(_10080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18976_ (.A1(_09831_),
    .A2(_07707_),
    .ZN(_10081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18977_ (.A1(_10071_),
    .A2(_09895_),
    .A3(_10081_),
    .ZN(_10082_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18978_ (.A1(_10080_),
    .A2(_10082_),
    .A3(_00398_),
    .ZN(_10083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18979_ (.A1(_10077_),
    .A2(_10083_),
    .B(_09938_),
    .ZN(_10084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18980_ (.A1(_10070_),
    .A2(_10084_),
    .ZN(_10085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18981_ (.A1(_09793_),
    .A2(_09784_),
    .A3(_09879_),
    .ZN(_10086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18982_ (.A1(_09934_),
    .A2(_10086_),
    .B(_09776_),
    .ZN(_10087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18983_ (.I(_10002_),
    .ZN(_10088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18984_ (.A1(_10087_),
    .A2(_10088_),
    .B(_09859_),
    .ZN(_10089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18985_ (.A1(_09812_),
    .A2(_09958_),
    .ZN(_10090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18986_ (.A1(_09884_),
    .A2(_09842_),
    .ZN(_10091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18987_ (.A1(_09827_),
    .A2(_09746_),
    .ZN(_10092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18988_ (.A1(_10092_),
    .A2(_09879_),
    .ZN(_10093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18989_ (.A1(_10091_),
    .A2(_10093_),
    .A3(_09776_),
    .ZN(_10094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18990_ (.A1(_10090_),
    .A2(_10094_),
    .A3(_09789_),
    .ZN(_10095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18991_ (.A1(_10089_),
    .A2(_10095_),
    .A3(_00398_),
    .ZN(_10096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18992_ (.A1(_09842_),
    .A2(_09784_),
    .A3(_09832_),
    .ZN(_10097_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18993_ (.A1(_09827_),
    .A2(_09940_),
    .A3(_09752_),
    .ZN(_10098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18994_ (.A1(_10097_),
    .A2(_10098_),
    .A3(_09834_),
    .ZN(_10099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18995_ (.A1(_09747_),
    .A2(_09832_),
    .ZN(_10100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18996_ (.A1(_10005_),
    .A2(_09807_),
    .A3(_10100_),
    .ZN(_10101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18997_ (.A1(_10099_),
    .A2(_10101_),
    .B(_00396_),
    .ZN(_10102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18998_ (.A1(_15664_),
    .A2(_15651_),
    .ZN(_10103_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18999_ (.A1(_09778_),
    .A2(_10103_),
    .A3(_09868_),
    .ZN(_10104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19000_ (.A1(_10047_),
    .A2(_09924_),
    .ZN(_10105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19001_ (.A1(_10104_),
    .A2(_10105_),
    .ZN(_10106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19002_ (.A1(_09865_),
    .A2(_07727_),
    .ZN(_10107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19003_ (.A1(_09805_),
    .A2(_10107_),
    .ZN(_10108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19004_ (.A1(_09834_),
    .A2(_10106_),
    .B(_10108_),
    .ZN(_10109_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19005_ (.A1(_10102_),
    .A2(_10109_),
    .B(_09823_),
    .ZN(_10110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19006_ (.A1(_10096_),
    .A2(_10110_),
    .A3(_09938_),
    .ZN(_10111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19007_ (.A1(_10085_),
    .A2(_10111_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19008_ (.A1(_00395_),
    .A2(net761),
    .B(_09893_),
    .ZN(_10112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19009_ (.A1(_09874_),
    .A2(_09842_),
    .ZN(_10113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19010_ (.A1(_09737_),
    .A2(_09908_),
    .Z(_10114_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19011_ (.A1(_10113_),
    .A2(_10114_),
    .B(_09807_),
    .ZN(_10115_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19012_ (.A1(_10112_),
    .A2(_09862_),
    .B(_10115_),
    .ZN(_10116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19013_ (.A1(_09954_),
    .A2(net765),
    .ZN(_10117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19014_ (.A1(_09744_),
    .A2(_10117_),
    .ZN(_10118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19015_ (.A1(_09885_),
    .A2(_09924_),
    .B(_09908_),
    .ZN(_10119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19016_ (.A1(_09917_),
    .A2(_09769_),
    .ZN(_10120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19017_ (.A1(_10119_),
    .A2(_10120_),
    .B(_09834_),
    .ZN(_10121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19018_ (.A1(_10118_),
    .A2(_10121_),
    .B(_09763_),
    .ZN(_10122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19019_ (.A1(_10116_),
    .A2(_10122_),
    .ZN(_10123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19020_ (.A1(_09793_),
    .A2(_07707_),
    .ZN(_10124_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19021_ (.A1(_10124_),
    .A2(_09942_),
    .Z(_10125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19022_ (.A1(_09803_),
    .A2(_09868_),
    .ZN(_10126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19023_ (.A1(_10125_),
    .A2(_00396_),
    .A3(_10126_),
    .ZN(_10127_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19024_ (.A1(_09879_),
    .A2(_15641_),
    .B(_09786_),
    .ZN(_10128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19025_ (.I(_10128_),
    .ZN(_10129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19026_ (.A1(_09779_),
    .A2(_00395_),
    .ZN(_10130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19027_ (.A1(_10129_),
    .A2(_10130_),
    .B(_09834_),
    .ZN(_10131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19028_ (.A1(_10127_),
    .A2(_10131_),
    .B(_09951_),
    .ZN(_10132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19029_ (.A1(_09770_),
    .A2(_09880_),
    .A3(_09895_),
    .ZN(_10133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19030_ (.A1(_09965_),
    .A2(_09847_),
    .ZN(_10134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19031_ (.A1(_10134_),
    .A2(_09748_),
    .ZN(_10135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19032_ (.A1(_10135_),
    .A2(_10086_),
    .A3(_09844_),
    .ZN(_10136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19033_ (.A1(_10133_),
    .A2(_10136_),
    .A3(_09859_),
    .ZN(_10137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19034_ (.A1(_10132_),
    .A2(_10137_),
    .ZN(_10138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19035_ (.A1(_10123_),
    .A2(_10138_),
    .B(_00399_),
    .ZN(_10139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19036_ (.A1(_09929_),
    .A2(_10040_),
    .ZN(_10140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19037_ (.A1(_10140_),
    .A2(_07726_),
    .ZN(_10141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19038_ (.A1(_09928_),
    .A2(_09838_),
    .A3(_07707_),
    .ZN(_10142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19039_ (.A1(_10142_),
    .A2(_09922_),
    .ZN(_10143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19040_ (.A1(_10143_),
    .A2(_09807_),
    .ZN(_10144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19041_ (.A1(_10141_),
    .A2(_09895_),
    .A3(_10144_),
    .ZN(_10145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19042_ (.I(_09768_),
    .ZN(_10146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19043_ (.A1(_10124_),
    .A2(_10146_),
    .ZN(_10147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19044_ (.A1(_10147_),
    .A2(_09807_),
    .B(_09797_),
    .ZN(_10148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19045_ (.A1(_09778_),
    .A2(_09766_),
    .A3(_09879_),
    .ZN(_10149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19046_ (.A1(_10135_),
    .A2(_10149_),
    .A3(_07726_),
    .ZN(_10150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19047_ (.A1(_10148_),
    .A2(_10150_),
    .B(_09762_),
    .ZN(_10151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19048_ (.A1(_10145_),
    .A2(_10151_),
    .ZN(_10152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19049_ (.A1(_10152_),
    .A2(_00399_),
    .ZN(_10153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19050_ (.I(_10046_),
    .ZN(_10154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19051_ (.A1(_10154_),
    .A2(_09854_),
    .ZN(_10155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19052_ (.A1(_10155_),
    .A2(_09844_),
    .A3(_09985_),
    .ZN(_10156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19053_ (.I(_09811_),
    .ZN(_10157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19054_ (.A1(_09738_),
    .A2(net37),
    .ZN(_10158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19055_ (.A1(_10157_),
    .A2(_09949_),
    .A3(_10158_),
    .ZN(_10159_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19056_ (.A1(_10156_),
    .A2(_10159_),
    .A3(_09834_),
    .ZN(_10160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19057_ (.A1(_09915_),
    .A2(_09863_),
    .ZN(_10161_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19058_ (.A1(_10161_),
    .A2(_09947_),
    .A3(_09796_),
    .ZN(_10162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19059_ (.A1(_09902_),
    .A2(_09750_),
    .Z(_10163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19060_ (.A1(_09760_),
    .A2(_09746_),
    .Z(_10164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19061_ (.A1(_10163_),
    .A2(_10164_),
    .ZN(_10165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19062_ (.A1(_10162_),
    .A2(_10165_),
    .A3(_09789_),
    .ZN(_10166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19063_ (.A1(_10166_),
    .A2(_10160_),
    .B(_00398_),
    .ZN(_10167_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19064_ (.A1(_10167_),
    .A2(_10153_),
    .ZN(_10168_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19065_ (.A1(_10139_),
    .A2(_10168_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19066_ (.A1(_09831_),
    .A2(_09840_),
    .Z(_10169_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19067_ (.A1(_09793_),
    .A2(_09847_),
    .A3(_09759_),
    .Z(_10170_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _19068_ (.A1(_10169_),
    .A2(_10170_),
    .A3(_09787_),
    .Z(_10171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19069_ (.A1(_00395_),
    .A2(net25),
    .B(_09829_),
    .ZN(_10172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19070_ (.A1(_09876_),
    .A2(_10172_),
    .B(_09762_),
    .ZN(_10173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19071_ (.A1(_10171_),
    .A2(_10173_),
    .ZN(_10174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19072_ (.A1(_09831_),
    .A2(_09923_),
    .A3(_09988_),
    .ZN(_10175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19073_ (.I(_10023_),
    .ZN(_10176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19074_ (.A1(_10175_),
    .A2(_10176_),
    .A3(_09895_),
    .ZN(_10177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19075_ (.I(_09973_),
    .ZN(_10178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19076_ (.A1(_09941_),
    .A2(_10178_),
    .ZN(_10179_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19077_ (.A1(_10177_),
    .A2(_10179_),
    .A3(_09763_),
    .ZN(_10180_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19078_ (.A1(_10174_),
    .A2(_00397_),
    .A3(_10180_),
    .ZN(_10181_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19079_ (.A1(_09990_),
    .A2(_09838_),
    .A3(_09988_),
    .Z(_10182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19080_ (.A1(_09800_),
    .A2(_09924_),
    .B(_09797_),
    .ZN(_10183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19081_ (.A1(_10062_),
    .A2(net840),
    .ZN(_10184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19082_ (.A1(_10183_),
    .A2(_10184_),
    .ZN(_10185_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19083_ (.A1(_09745_),
    .A2(_10182_),
    .B(_10185_),
    .C(_09951_),
    .ZN(_10186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19084_ (.A1(_09795_),
    .A2(_09782_),
    .ZN(_10187_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19085_ (.A1(_10061_),
    .A2(_09908_),
    .A3(_10187_),
    .Z(_10188_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19086_ (.A1(_10188_),
    .A2(_09951_),
    .ZN(_10189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19087_ (.A1(_09840_),
    .A2(_10103_),
    .ZN(_10190_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19088_ (.A1(net840),
    .A2(net822),
    .A3(_09868_),
    .ZN(_10191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19089_ (.A1(_10190_),
    .A2(_10191_),
    .A3(_09844_),
    .ZN(_10192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19090_ (.A1(_10189_),
    .A2(_10192_),
    .B(_09789_),
    .ZN(_10193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19091_ (.A1(_10186_),
    .A2(_10193_),
    .ZN(_10194_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19092_ (.A1(_09938_),
    .A2(_10181_),
    .A3(_10194_),
    .ZN(_10195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19093_ (.A1(_10001_),
    .A2(net760),
    .ZN(_10196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19094_ (.A1(_09882_),
    .A2(_10196_),
    .B(_09951_),
    .ZN(_10197_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19095_ (.A1(_09778_),
    .A2(_09917_),
    .A3(_09988_),
    .ZN(_10198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19096_ (.A1(_10163_),
    .A2(_10198_),
    .ZN(_10199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19097_ (.A1(_10197_),
    .A2(_10199_),
    .B(_09789_),
    .ZN(_10200_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19098_ (.A1(_09954_),
    .A2(_09797_),
    .A3(_09959_),
    .Z(_10201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19099_ (.A1(_10093_),
    .A2(_09947_),
    .A3(_09883_),
    .ZN(_10202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19100_ (.A1(_10201_),
    .A2(_10202_),
    .A3(_09951_),
    .ZN(_10203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19101_ (.A1(_10200_),
    .A2(_10203_),
    .B(_09938_),
    .ZN(_10204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19102_ (.A1(_09832_),
    .A2(net11),
    .ZN(_10205_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19103_ (.A1(_10135_),
    .A2(_09797_),
    .A3(_10205_),
    .Z(_10206_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19104_ (.A1(_09933_),
    .A2(_09988_),
    .B(_09829_),
    .ZN(_10207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19105_ (.A1(_09828_),
    .A2(_09965_),
    .Z(_10208_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19106_ (.A1(_10207_),
    .A2(_10208_),
    .ZN(_10209_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19107_ (.A1(_10206_),
    .A2(_10209_),
    .B(_09823_),
    .ZN(_10210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19108_ (.A1(_09973_),
    .A2(_09772_),
    .ZN(_10211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19109_ (.A1(_09857_),
    .A2(_09895_),
    .A3(_10211_),
    .ZN(_10212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19110_ (.A1(_10078_),
    .A2(_09794_),
    .ZN(_10213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19111_ (.A1(_10023_),
    .A2(_09990_),
    .ZN(_10214_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19112_ (.A1(_10213_),
    .A2(_10214_),
    .A3(_09844_),
    .ZN(_10215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19113_ (.A1(_10212_),
    .A2(_10215_),
    .A3(_09951_),
    .ZN(_10216_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19114_ (.A1(_10210_),
    .A2(_10216_),
    .A3(_00397_),
    .ZN(_10217_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19115_ (.A1(_10204_),
    .A2(_10217_),
    .ZN(_10218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19116_ (.A1(_10195_),
    .A2(_10218_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19117_ (.A1(net765),
    .A2(_09784_),
    .A3(_09940_),
    .ZN(_10219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19118_ (.A1(_10093_),
    .A2(_10219_),
    .A3(_00396_),
    .ZN(_10220_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19119_ (.A1(_15659_),
    .A2(_15641_),
    .ZN(_10221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19120_ (.A1(_10221_),
    .A2(_00395_),
    .B(_09829_),
    .ZN(_10222_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19121_ (.A1(_09793_),
    .A2(_09849_),
    .A3(_09940_),
    .ZN(_10223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19122_ (.A1(_09768_),
    .A2(_00395_),
    .ZN(_10224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19123_ (.A1(_10222_),
    .A2(_10223_),
    .A3(_10224_),
    .ZN(_10225_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19124_ (.A1(_10220_),
    .A2(_10225_),
    .A3(_00398_),
    .ZN(_10226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19125_ (.A1(_09813_),
    .A2(_09794_),
    .A3(_09924_),
    .ZN(_10227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19126_ (.A1(_10219_),
    .A2(_10227_),
    .A3(_09895_),
    .ZN(_10228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19127_ (.A1(_09800_),
    .A2(_09988_),
    .B(_09797_),
    .ZN(_10229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19128_ (.A1(_10154_),
    .A2(_09928_),
    .ZN(_10230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19129_ (.A1(_10229_),
    .A2(_10230_),
    .ZN(_10231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19130_ (.A1(_10228_),
    .A2(_10231_),
    .A3(_09763_),
    .ZN(_10232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19131_ (.A1(_10226_),
    .A2(_10232_),
    .A3(_09859_),
    .ZN(_10233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19132_ (.A1(_09867_),
    .A2(_09988_),
    .B(_09797_),
    .ZN(_10234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19133_ (.A1(_10012_),
    .A2(_09746_),
    .ZN(_10235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19134_ (.A1(_10235_),
    .A2(_00395_),
    .ZN(_10236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19135_ (.A1(_10234_),
    .A2(_10236_),
    .B(_09762_),
    .ZN(_10237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19136_ (.A1(_10134_),
    .A2(_09924_),
    .ZN(_10238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19137_ (.A1(_09988_),
    .A2(net11),
    .B(_09829_),
    .ZN(_10239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19138_ (.A1(_10238_),
    .A2(_10239_),
    .ZN(_10240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19139_ (.A1(_10237_),
    .A2(_10240_),
    .B(_09834_),
    .ZN(_10241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19140_ (.I(net822),
    .ZN(_10242_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19141_ (.A1(_10120_),
    .A2(_10242_),
    .ZN(_10243_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19142_ (.A1(_10081_),
    .A2(_09942_),
    .ZN(_10244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19143_ (.A1(_10243_),
    .A2(_10244_),
    .B(_09787_),
    .ZN(_10245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19144_ (.A1(_09884_),
    .A2(_09831_),
    .ZN(_10246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19145_ (.A1(_10246_),
    .A2(_10031_),
    .ZN(_10247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19146_ (.A1(_10247_),
    .A2(_09776_),
    .ZN(_10248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19147_ (.A1(_10248_),
    .A2(_10245_),
    .ZN(_10249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19148_ (.A1(_10249_),
    .A2(_09823_),
    .ZN(_10250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19149_ (.A1(_10250_),
    .A2(_10241_),
    .ZN(_10251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19150_ (.A1(_10233_),
    .A2(_10251_),
    .B(_09938_),
    .ZN(_10252_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19151_ (.A1(_09959_),
    .A2(_09942_),
    .A3(_09795_),
    .Z(_10253_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19152_ (.A1(_09900_),
    .A2(_09759_),
    .A3(_09878_),
    .Z(_10254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19153_ (.A1(_10253_),
    .A2(_10254_),
    .A3(_09787_),
    .ZN(_10255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19154_ (.A1(_10255_),
    .A2(_09951_),
    .ZN(_10256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19155_ (.A1(_09915_),
    .A2(_09813_),
    .ZN(_10257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19156_ (.A1(_10254_),
    .A2(_10257_),
    .B(_09947_),
    .ZN(_10258_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19157_ (.A1(_10256_),
    .A2(_10258_),
    .ZN(_10259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19158_ (.A1(_09912_),
    .A2(_09773_),
    .ZN(_10260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19159_ (.I(_10260_),
    .ZN(_10261_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19160_ (.A1(_10261_),
    .A2(_09842_),
    .Z(_10262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19161_ (.A1(_09901_),
    .A2(_09750_),
    .ZN(_10263_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19162_ (.A1(_10262_),
    .A2(_10263_),
    .ZN(_10264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19163_ (.A1(_09795_),
    .A2(_15661_),
    .ZN(_10265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19164_ (.A1(_10265_),
    .A2(_09908_),
    .ZN(_10266_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19165_ (.A1(_10170_),
    .A2(_10266_),
    .ZN(_10267_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19166_ (.A1(_10264_),
    .A2(_10267_),
    .B(_09763_),
    .ZN(_10268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19167_ (.A1(_10268_),
    .A2(_00397_),
    .ZN(_10269_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19168_ (.A1(_10259_),
    .A2(_10269_),
    .ZN(_10270_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19169_ (.I(_09943_),
    .ZN(_10271_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19170_ (.A1(_09839_),
    .A2(_09776_),
    .A3(_10271_),
    .ZN(_10272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19171_ (.A1(_10242_),
    .A2(_09868_),
    .ZN(_10273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19172_ (.A1(_10093_),
    .A2(_09947_),
    .A3(_10273_),
    .ZN(_10274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19173_ (.A1(_10272_),
    .A2(_10274_),
    .B(_09763_),
    .ZN(_10275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19174_ (.A1(_10103_),
    .A2(_09769_),
    .ZN(_10276_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19175_ (.A1(_10124_),
    .A2(_09942_),
    .B(_10276_),
    .ZN(_10277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19176_ (.A1(_10277_),
    .A2(_09829_),
    .ZN(_10278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19177_ (.A1(_09982_),
    .A2(_09797_),
    .B(_07735_),
    .ZN(_10279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19178_ (.A1(_10278_),
    .A2(_10279_),
    .ZN(_10280_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19179_ (.A1(_10280_),
    .A2(_09859_),
    .ZN(_10281_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19180_ (.A1(_10275_),
    .A2(_10281_),
    .B(_09938_),
    .ZN(_10282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19181_ (.A1(_10270_),
    .A2(_10282_),
    .ZN(_10283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19182_ (.A1(_10283_),
    .A2(_10252_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19183_ (.A1(_10098_),
    .A2(_00396_),
    .A3(_09946_),
    .ZN(_10284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19184_ (.A1(_10044_),
    .A2(_10223_),
    .A3(_09947_),
    .ZN(_10285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19185_ (.A1(_10284_),
    .A2(_10285_),
    .A3(_09859_),
    .ZN(_10286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19186_ (.A1(_09914_),
    .A2(_09908_),
    .Z(_10287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19187_ (.A1(_10125_),
    .A2(_10287_),
    .B(_09834_),
    .ZN(_10288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19188_ (.A1(_09828_),
    .A2(_09794_),
    .ZN(_10289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19189_ (.A1(_09867_),
    .A2(_00395_),
    .ZN(_10290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19190_ (.A1(_10221_),
    .A2(_09832_),
    .B(_09908_),
    .ZN(_10291_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19191_ (.A1(_10289_),
    .A2(_10290_),
    .A3(_10291_),
    .ZN(_10292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19192_ (.A1(_10288_),
    .A2(_10292_),
    .ZN(_10293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19193_ (.A1(_10293_),
    .A2(_10286_),
    .B(_09823_),
    .ZN(_10294_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19194_ (.A1(_09885_),
    .A2(_09912_),
    .A3(_09769_),
    .Z(_10295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19195_ (.A1(_10046_),
    .A2(_09750_),
    .ZN(_10296_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19196_ (.A1(_10295_),
    .A2(_10296_),
    .ZN(_10297_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19197_ (.A1(_09865_),
    .A2(_09743_),
    .ZN(_10298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19198_ (.A1(_10297_),
    .A2(_10298_),
    .B(_09834_),
    .ZN(_10299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19199_ (.A1(_10299_),
    .A2(_09823_),
    .ZN(_10300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19200_ (.A1(_09885_),
    .A2(_09847_),
    .A3(_09769_),
    .ZN(_10301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19201_ (.A1(_10301_),
    .A2(_10040_),
    .ZN(_10302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19202_ (.A1(_10302_),
    .A2(_09787_),
    .ZN(_10303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19203_ (.A1(_09748_),
    .A2(net758),
    .ZN(_10304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19204_ (.A1(_10142_),
    .A2(_09829_),
    .A3(_10304_),
    .ZN(_10305_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19205_ (.A1(_10303_),
    .A2(_09789_),
    .A3(_10305_),
    .Z(_10306_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19206_ (.A1(_10300_),
    .A2(_10306_),
    .ZN(_10307_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19207_ (.A1(_10294_),
    .A2(_10307_),
    .B(_09938_),
    .ZN(_10308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19208_ (.A1(_09795_),
    .A2(_15671_),
    .Z(_10309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19209_ (.A1(_09988_),
    .A2(_10047_),
    .B(_10309_),
    .ZN(_10310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19210_ (.A1(_10310_),
    .A2(_09996_),
    .B(_09807_),
    .ZN(_10311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19211_ (.I(_10263_),
    .ZN(_10312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19212_ (.A1(_10261_),
    .A2(_09863_),
    .ZN(_10313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19213_ (.A1(_10312_),
    .A2(_10048_),
    .A3(_10313_),
    .ZN(_10314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19214_ (.A1(_10311_),
    .A2(_10314_),
    .ZN(_10315_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19215_ (.I(_09862_),
    .ZN(_10316_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19216_ (.A1(_10316_),
    .A2(_10126_),
    .A3(_09893_),
    .ZN(_10317_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19217_ (.A1(_10012_),
    .A2(_09879_),
    .ZN(_10318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19218_ (.I(_10318_),
    .ZN(_10319_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19219_ (.A1(_09924_),
    .A2(_09740_),
    .B(_09750_),
    .ZN(_10320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19220_ (.A1(_10319_),
    .A2(_10320_),
    .B(_09834_),
    .ZN(_10321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19221_ (.A1(_10317_),
    .A2(_10321_),
    .ZN(_10322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19222_ (.A1(_10315_),
    .A2(_10322_),
    .A3(_09823_),
    .ZN(_10323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19223_ (.A1(net761),
    .A2(_09786_),
    .ZN(_10324_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19224_ (.A1(_10318_),
    .A2(_10324_),
    .ZN(_10325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19225_ (.A1(_09855_),
    .A2(_00395_),
    .ZN(_10326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19226_ (.A1(_10325_),
    .A2(_10326_),
    .B(_09807_),
    .ZN(_10327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19227_ (.A1(_10238_),
    .A2(_09844_),
    .A3(_09976_),
    .ZN(_10328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19228_ (.A1(_10327_),
    .A2(_10328_),
    .B(_09763_),
    .ZN(_10329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19229_ (.A1(_10261_),
    .A2(_10103_),
    .ZN(_10330_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19230_ (.A1(_09867_),
    .A2(_10221_),
    .B(_09868_),
    .ZN(_10331_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19231_ (.A1(_10330_),
    .A2(_10331_),
    .A3(_09895_),
    .ZN(_10332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19232_ (.A1(_09778_),
    .A2(_09885_),
    .A3(_09868_),
    .ZN(_10333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19233_ (.A1(_10333_),
    .A2(_10086_),
    .A3(_09776_),
    .ZN(_10334_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19234_ (.A1(_10332_),
    .A2(_00397_),
    .A3(_10334_),
    .ZN(_10335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19235_ (.A1(_10329_),
    .A2(_10335_),
    .ZN(_10336_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19236_ (.A1(_10323_),
    .A2(_10336_),
    .A3(_00399_),
    .ZN(_10337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19237_ (.A1(_10308_),
    .A2(_10337_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19238_ (.I(\sa00_sr[7] ),
    .ZN(_10338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19239_ (.I(\sa00_sr[0] ),
    .ZN(_10339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19240_ (.A1(_10338_),
    .A2(_10339_),
    .ZN(_10340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19241_ (.A1(\sa00_sr[7] ),
    .A2(net695),
    .ZN(_10341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19242_ (.A1(_10341_),
    .A2(_10340_),
    .ZN(_10342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19243_ (.I(net688),
    .ZN(_10343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19244_ (.A1(_10343_),
    .A2(\sa20_sr[1] ),
    .ZN(_10344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19245_ (.I(net875),
    .ZN(_10345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19246_ (.A1(_10345_),
    .A2(net687),
    .ZN(_10346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19247_ (.A1(_10344_),
    .A2(_10346_),
    .ZN(_10347_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19248_ (.A1(_10342_),
    .A2(_10347_),
    .ZN(_10348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19249_ (.A1(_10339_),
    .A2(\sa00_sr[7] ),
    .ZN(_10349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19250_ (.A1(_10338_),
    .A2(net695),
    .ZN(_10350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19251_ (.A1(_10350_),
    .A2(_10349_),
    .ZN(_10351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19252_ (.A1(_10345_),
    .A2(_10343_),
    .ZN(_10352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19253_ (.A1(net874),
    .A2(net1078),
    .ZN(_10353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19254_ (.A1(_10353_),
    .A2(_10352_),
    .ZN(_10354_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19255_ (.A1(_10354_),
    .A2(_10351_),
    .ZN(_10355_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19256_ (.A1(_10348_),
    .A2(_10355_),
    .ZN(_10356_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19257_ (.I(\sa10_sr[0] ),
    .ZN(_10357_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19258_ (.I(\sa10_sr[7] ),
    .Z(_10358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19259_ (.A1(_10358_),
    .A2(_10357_),
    .ZN(_10359_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19260_ (.I(\sa10_sr[7] ),
    .ZN(_10360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19261_ (.A1(_10360_),
    .A2(\sa10_sr[0] ),
    .ZN(_10361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19262_ (.A1(_10359_),
    .A2(_10361_),
    .ZN(_10362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19263_ (.A1(net866),
    .A2(net492),
    .ZN(_10363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19264_ (.A1(_10357_),
    .A2(_10360_),
    .ZN(_10364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19265_ (.A1(\sa10_sr[7] ),
    .A2(\sa10_sr[0] ),
    .ZN(_10365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19266_ (.A1(_10365_),
    .A2(_10364_),
    .ZN(_10366_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19267_ (.I(\sa10_sr[1] ),
    .ZN(_10367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19268_ (.A1(_10366_),
    .A2(_10367_),
    .ZN(_10368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19269_ (.A1(_10363_),
    .A2(_10368_),
    .ZN(_10369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19270_ (.A1(_10369_),
    .A2(_10356_),
    .ZN(_10370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19271_ (.A1(_10354_),
    .A2(_10351_),
    .ZN(_10371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19272_ (.A1(_10342_),
    .A2(_10347_),
    .ZN(_10372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19273_ (.A1(_10371_),
    .A2(_10372_),
    .ZN(_10373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19274_ (.A1(_10366_),
    .A2(net492),
    .ZN(_10374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19275_ (.A1(_10362_),
    .A2(_10367_),
    .ZN(_10375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19276_ (.A1(_10374_),
    .A2(_10375_),
    .ZN(_10376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19277_ (.A1(_10373_),
    .A2(_10376_),
    .ZN(_10377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _19278_ (.I(net477),
    .ZN(_10378_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _19279_ (.I(_10378_),
    .Z(_10379_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19280_ (.A1(net811),
    .A2(_10377_),
    .A3(_10370_),
    .ZN(_10380_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19281_ (.I(net477),
    .Z(_10381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19282_ (.A1(\text_in_r[121] ),
    .A2(_10381_),
    .ZN(_10382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19283_ (.A1(_10380_),
    .A2(_10382_),
    .ZN(_10383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19284_ (.I(net630),
    .ZN(_10384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19285_ (.A1(_10383_),
    .A2(_10384_),
    .ZN(_10385_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19286_ (.A1(net827),
    .A2(net630),
    .A3(_10382_),
    .ZN(_10386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19287_ (.A1(_10386_),
    .A2(_10385_),
    .ZN(_15679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19288_ (.A1(_10338_),
    .A2(_10360_),
    .ZN(_10387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19289_ (.A1(\sa00_sr[7] ),
    .A2(_10358_),
    .ZN(_10388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19290_ (.A1(_10387_),
    .A2(_10388_),
    .ZN(_10389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19291_ (.A1(_10389_),
    .A2(net583),
    .ZN(_10390_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19292_ (.I(\sa30_sr[0] ),
    .ZN(_10391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19293_ (.A1(_10387_),
    .A2(_10391_),
    .A3(_10388_),
    .ZN(_10392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19294_ (.A1(_10390_),
    .A2(_10392_),
    .ZN(_10393_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19295_ (.I(\sa20_sr[0] ),
    .ZN(_10394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19296_ (.A1(_10357_),
    .A2(_10394_),
    .ZN(_10395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19297_ (.A1(net679),
    .A2(net577),
    .ZN(_10396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19298_ (.A1(_10395_),
    .A2(_10396_),
    .ZN(_10397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19299_ (.I(_10397_),
    .ZN(_10398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19300_ (.A1(_10393_),
    .A2(_10398_),
    .ZN(_10399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19301_ (.A1(_10390_),
    .A2(_10392_),
    .A3(_10397_),
    .ZN(_10400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19302_ (.A1(_10399_),
    .A2(_10400_),
    .ZN(_10401_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19303_ (.I(_10378_),
    .Z(_10402_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _19304_ (.I(_10402_),
    .Z(_10403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19305_ (.A1(_10401_),
    .A2(_10403_),
    .ZN(_10404_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19306_ (.I(_10379_),
    .Z(_10405_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19307_ (.A1(_10405_),
    .A2(\text_in_r[120] ),
    .Z(_10406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19308_ (.A1(_10404_),
    .A2(_07672_),
    .A3(_10406_),
    .ZN(_10407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19309_ (.A1(_10399_),
    .A2(_10400_),
    .A3(_10403_),
    .ZN(_10408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19310_ (.I(net475),
    .Z(_10409_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _19311_ (.I(_10409_),
    .Z(_10410_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _19312_ (.I(_10410_),
    .Z(_10411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19313_ (.A1(_10411_),
    .A2(\text_in_r[120] ),
    .ZN(_10412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19314_ (.A1(_10408_),
    .A2(\u0.w[0][24] ),
    .A3(_10412_),
    .ZN(_10413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19315_ (.A1(_10407_),
    .A2(_10413_),
    .ZN(_15682_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19316_ (.I(\sa00_sr[1] ),
    .ZN(_10414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19317_ (.A1(_10414_),
    .A2(\sa10_sr[1] ),
    .ZN(_10415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19318_ (.A1(_10367_),
    .A2(net618),
    .ZN(_10416_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _19319_ (.I(\sa20_sr[2] ),
    .ZN(_10417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19320_ (.A1(_10415_),
    .A2(_10416_),
    .A3(_10417_),
    .ZN(_10418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19321_ (.A1(_10367_),
    .A2(_10414_),
    .ZN(_10419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19322_ (.A1(\sa10_sr[1] ),
    .A2(net618),
    .ZN(_10420_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19323_ (.A1(_10419_),
    .A2(\sa20_sr[2] ),
    .A3(_10420_),
    .ZN(_10421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19324_ (.A1(_10418_),
    .A2(_10421_),
    .ZN(_10422_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19325_ (.I(\sa30_sr[2] ),
    .ZN(_10423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19326_ (.A1(_10423_),
    .A2(net861),
    .ZN(_10424_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19327_ (.I(\sa10_sr[2] ),
    .ZN(_10425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19328_ (.A1(_10425_),
    .A2(\sa30_sr[2] ),
    .ZN(_10426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19329_ (.A1(_10424_),
    .A2(_10426_),
    .ZN(_10427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19330_ (.I(_10427_),
    .ZN(_10428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19331_ (.A1(_10422_),
    .A2(_10428_),
    .ZN(_10429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19332_ (.A1(_10418_),
    .A2(_10421_),
    .A3(_10427_),
    .ZN(_10430_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _19333_ (.I(net475),
    .Z(_10431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _19334_ (.A1(_10429_),
    .A2(_10430_),
    .B(_10431_),
    .ZN(_10432_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19335_ (.I(\text_in_r[122] ),
    .ZN(_10433_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19336_ (.A1(_10433_),
    .A2(net594),
    .Z(_10434_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19337_ (.A1(_10432_),
    .A2(_10434_),
    .B(_07689_),
    .ZN(_10435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19338_ (.A1(_10429_),
    .A2(_10430_),
    .ZN(_10436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19339_ (.A1(_10436_),
    .A2(net811),
    .ZN(_10437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19340_ (.I(_10434_),
    .ZN(_10438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19341_ (.A1(_10437_),
    .A2(\u0.w[0][26] ),
    .A3(_10438_),
    .ZN(_10439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19342_ (.A1(_10435_),
    .A2(_10439_),
    .ZN(_10440_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19343_ (.I(_10440_),
    .Z(_15698_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19344_ (.A1(_10404_),
    .A2(\u0.w[0][24] ),
    .A3(_10406_),
    .ZN(_10441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19345_ (.A1(_10408_),
    .A2(_07672_),
    .A3(_10412_),
    .ZN(_10442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19346_ (.A1(_10441_),
    .A2(_10442_),
    .ZN(_15673_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _19347_ (.A1(_10432_),
    .A2(_10434_),
    .B(\u0.w[0][26] ),
    .ZN(_10443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19348_ (.A1(_10437_),
    .A2(_10438_),
    .A3(_07689_),
    .ZN(_10444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19349_ (.A1(_10443_),
    .A2(_10444_),
    .ZN(_10445_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _19350_ (.I(_10445_),
    .Z(_15691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19351_ (.A1(net599),
    .A2(_10445_),
    .ZN(_10446_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19352_ (.I(_10446_),
    .ZN(_10447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19353_ (.A1(_10447_),
    .A2(net33),
    .ZN(_10448_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19354_ (.A1(\sa20_sr[3] ),
    .A2(\sa30_sr[3] ),
    .Z(_10449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19355_ (.I(\sa00_sr[2] ),
    .ZN(_10450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19356_ (.A1(_10338_),
    .A2(_10450_),
    .ZN(_10451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19357_ (.A1(net76),
    .A2(\sa00_sr[2] ),
    .ZN(_10452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19358_ (.A1(_10451_),
    .A2(_10452_),
    .ZN(_10453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19359_ (.A1(_10449_),
    .A2(_10453_),
    .ZN(_10454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19360_ (.A1(_10450_),
    .A2(net76),
    .ZN(_10455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19361_ (.A1(_10338_),
    .A2(\sa00_sr[2] ),
    .ZN(_10456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19362_ (.A1(_10455_),
    .A2(_10456_),
    .ZN(_10457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19363_ (.I(\sa20_sr[3] ),
    .ZN(_10458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19364_ (.I(\sa30_sr[3] ),
    .ZN(_10459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19365_ (.A1(_10458_),
    .A2(_10459_),
    .ZN(_10460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19366_ (.A1(\sa20_sr[3] ),
    .A2(\sa30_sr[3] ),
    .ZN(_10461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19367_ (.A1(_10460_),
    .A2(_10461_),
    .ZN(_10462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19368_ (.A1(_10457_),
    .A2(_10462_),
    .ZN(_10463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19369_ (.A1(_10454_),
    .A2(_10463_),
    .ZN(_10464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19370_ (.I(_10464_),
    .ZN(_10465_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19371_ (.I(\sa10_sr[3] ),
    .ZN(_10466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19372_ (.A1(_10466_),
    .A2(net46),
    .ZN(_10467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19373_ (.A1(net683),
    .A2(\sa10_sr[3] ),
    .ZN(_10468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19374_ (.A1(_10467_),
    .A2(_10468_),
    .ZN(_10469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19375_ (.A1(_10469_),
    .A2(\sa10_sr[2] ),
    .ZN(_10470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19376_ (.A1(net683),
    .A2(_10466_),
    .ZN(_10471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19377_ (.A1(net46),
    .A2(\sa10_sr[3] ),
    .ZN(_10472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19378_ (.A1(_10471_),
    .A2(_10472_),
    .ZN(_10473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19379_ (.A1(_10473_),
    .A2(_10425_),
    .ZN(_10474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19380_ (.A1(_10470_),
    .A2(_10474_),
    .ZN(_10475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19381_ (.A1(_10465_),
    .A2(_10475_),
    .ZN(_10476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19382_ (.I(_10475_),
    .ZN(_10477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19383_ (.A1(_10477_),
    .A2(_10464_),
    .ZN(_10478_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19384_ (.I(_10402_),
    .Z(_10479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19385_ (.A1(_10476_),
    .A2(_10478_),
    .A3(_10479_),
    .ZN(_10480_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19386_ (.I(\u0.w[0][27] ),
    .ZN(_10481_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _19387_ (.I(_10409_),
    .Z(_10482_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _19388_ (.I(_10482_),
    .Z(_10483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19389_ (.A1(_10483_),
    .A2(\text_in_r[123] ),
    .ZN(_10484_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19390_ (.A1(_10480_),
    .A2(_10481_),
    .A3(_10484_),
    .ZN(_10485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19391_ (.A1(_10465_),
    .A2(_10477_),
    .ZN(_10486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19392_ (.A1(_10464_),
    .A2(_10475_),
    .ZN(_10487_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19393_ (.A1(_10486_),
    .A2(_10479_),
    .A3(_10487_),
    .ZN(_10488_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19394_ (.I(_10379_),
    .Z(_10489_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19395_ (.A1(_10489_),
    .A2(\text_in_r[123] ),
    .Z(_10490_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19396_ (.A1(_10488_),
    .A2(\u0.w[0][27] ),
    .A3(_10490_),
    .ZN(_10491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19397_ (.A1(_10485_),
    .A2(_10491_),
    .ZN(_10492_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19398_ (.I(_10492_),
    .Z(_10493_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19399_ (.I(_15680_),
    .ZN(_10494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19400_ (.A1(_10440_),
    .A2(_10494_),
    .ZN(_10495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19401_ (.A1(_10448_),
    .A2(_10493_),
    .A3(_10495_),
    .ZN(_10496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19402_ (.A1(_10440_),
    .A2(net829),
    .ZN(_10497_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19403_ (.I(_15675_),
    .ZN(_10498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19404_ (.A1(_10445_),
    .A2(_10498_),
    .ZN(_10499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19405_ (.A1(_10497_),
    .A2(_10499_),
    .ZN(_10500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19406_ (.A1(_10480_),
    .A2(\u0.w[0][27] ),
    .A3(_10484_),
    .ZN(_10501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19407_ (.A1(_10488_),
    .A2(_10481_),
    .A3(_10490_),
    .ZN(_10502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19408_ (.A1(_10501_),
    .A2(_10502_),
    .ZN(_10503_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19409_ (.I(_10503_),
    .Z(_10504_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19410_ (.I(_10504_),
    .Z(_10505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19411_ (.A1(_10500_),
    .A2(_10505_),
    .ZN(_10506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19412_ (.A1(_10443_),
    .A2(_10444_),
    .A3(_15677_),
    .ZN(_10507_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19413_ (.I(_10507_),
    .ZN(_10508_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19414_ (.I(_10492_),
    .Z(_10509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19415_ (.A1(_10508_),
    .A2(_10509_),
    .ZN(_10510_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19416_ (.A1(\sa00_sr[7] ),
    .A2(\sa00_sr[3] ),
    .Z(_10511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19417_ (.I(\sa20_sr[4] ),
    .ZN(_10512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19418_ (.A1(_10511_),
    .A2(_10512_),
    .Z(_10513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19419_ (.A1(_10511_),
    .A2(_10512_),
    .ZN(_10514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19420_ (.A1(_10513_),
    .A2(_10514_),
    .ZN(_10515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19421_ (.I(_10515_),
    .ZN(_10516_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19422_ (.A1(\sa10_sr[4] ),
    .A2(\sa30_sr[4] ),
    .Z(_10517_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19423_ (.A1(_10473_),
    .A2(_10517_),
    .Z(_10518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19424_ (.A1(_10516_),
    .A2(_10518_),
    .ZN(_10519_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19425_ (.A1(_10469_),
    .A2(_10517_),
    .Z(_10520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19426_ (.A1(_10520_),
    .A2(_10515_),
    .ZN(_10521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19427_ (.I(_10379_),
    .Z(_10522_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _19428_ (.I(_10522_),
    .Z(_10523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19429_ (.A1(_10519_),
    .A2(_10521_),
    .A3(_10523_),
    .ZN(_10524_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _19430_ (.I(_10431_),
    .Z(_10525_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _19431_ (.I(_10525_),
    .Z(_10526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19432_ (.A1(_10526_),
    .A2(\text_in_r[124] ),
    .ZN(_10527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19433_ (.A1(_10524_),
    .A2(_10527_),
    .ZN(_10528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19434_ (.A1(_10528_),
    .A2(\u0.w[0][28] ),
    .ZN(_10529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19435_ (.I(\u0.w[0][28] ),
    .ZN(_10530_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19436_ (.A1(_10524_),
    .A2(_10530_),
    .A3(_10527_),
    .ZN(_10531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19437_ (.A1(_10529_),
    .A2(_10531_),
    .ZN(_10532_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19438_ (.I(_10532_),
    .Z(_10533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19439_ (.A1(_10510_),
    .A2(_10533_),
    .Z(_10534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19440_ (.A1(_10496_),
    .A2(_10506_),
    .A3(_10534_),
    .ZN(_10535_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19441_ (.A1(_10443_),
    .A2(net608),
    .A3(net604),
    .ZN(_10536_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19442_ (.I(_10536_),
    .ZN(_10537_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19443_ (.I(_10532_),
    .Z(_10538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19444_ (.A1(_10537_),
    .A2(_10493_),
    .B(_10538_),
    .ZN(_10539_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19445_ (.I(_10504_),
    .Z(_10540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19446_ (.A1(_10540_),
    .A2(_15696_),
    .ZN(_10541_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19447_ (.A1(\sa10_sr[4] ),
    .A2(\sa00_sr[4] ),
    .Z(_10542_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19448_ (.A1(\sa20_sr[5] ),
    .A2(\sa30_sr[5] ),
    .Z(_10543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19449_ (.A1(\sa20_sr[5] ),
    .A2(\sa30_sr[5] ),
    .ZN(_10544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19450_ (.A1(_10543_),
    .A2(_10544_),
    .ZN(_10545_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19451_ (.A1(\sa10_sr[5] ),
    .A2(_10545_),
    .Z(_10546_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19452_ (.A1(_10542_),
    .A2(_10546_),
    .Z(_10547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19453_ (.A1(_10547_),
    .A2(_10523_),
    .ZN(_10548_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _19454_ (.I(_10379_),
    .Z(_10549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19455_ (.A1(_10549_),
    .A2(\text_in_r[125] ),
    .Z(_10550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19456_ (.A1(_10548_),
    .A2(_10550_),
    .ZN(_10551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19457_ (.I(\u0.w[0][29] ),
    .ZN(_10552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19458_ (.A1(_10551_),
    .A2(_10552_),
    .ZN(_10553_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19459_ (.A1(_10548_),
    .A2(\u0.w[0][29] ),
    .A3(_10550_),
    .ZN(_10554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19460_ (.A1(_10553_),
    .A2(_10554_),
    .ZN(_10555_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19461_ (.I(_10555_),
    .ZN(_10556_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19462_ (.I(_10556_),
    .Z(_10557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19463_ (.A1(_10539_),
    .A2(_10541_),
    .B(_10557_),
    .ZN(_10558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19464_ (.A1(_10535_),
    .A2(_10558_),
    .ZN(_10559_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19465_ (.I(_15685_),
    .ZN(_10560_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19466_ (.A1(_10443_),
    .A2(_10444_),
    .A3(_10560_),
    .ZN(_10561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19467_ (.A1(_10503_),
    .A2(_10561_),
    .Z(_10562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19468_ (.A1(_10448_),
    .A2(_10562_),
    .ZN(_10563_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19469_ (.I(_10538_),
    .Z(_10564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19470_ (.A1(_10445_),
    .A2(_15677_),
    .Z(_10565_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _19471_ (.I(_10492_),
    .Z(_10566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19472_ (.A1(_10565_),
    .A2(_10566_),
    .ZN(_10567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19473_ (.A1(_10563_),
    .A2(_10564_),
    .A3(_10567_),
    .ZN(_10568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19474_ (.A1(_10565_),
    .A2(_10504_),
    .ZN(_10569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19475_ (.A1(_10528_),
    .A2(_10530_),
    .ZN(_10570_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19476_ (.A1(_10524_),
    .A2(\u0.w[0][28] ),
    .A3(_10527_),
    .ZN(_10571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19477_ (.A1(_10570_),
    .A2(_10571_),
    .ZN(_10572_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19478_ (.I(_10572_),
    .Z(_10573_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19479_ (.A1(_10569_),
    .A2(_10573_),
    .Z(_10574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19480_ (.A1(_10440_),
    .A2(_15683_),
    .ZN(_10575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19481_ (.A1(_10575_),
    .A2(_10492_),
    .Z(_10576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19482_ (.A1(_10448_),
    .A2(_10576_),
    .ZN(_10577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19483_ (.A1(_10574_),
    .A2(_10577_),
    .ZN(_10578_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19484_ (.I(_10556_),
    .Z(_10579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19485_ (.A1(_10568_),
    .A2(_10578_),
    .A3(_10579_),
    .ZN(_10580_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _19486_ (.A1(\sa10_sr[5] ),
    .A2(\sa00_sr[5] ),
    .ZN(_10581_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _19487_ (.A1(\sa20_sr[6] ),
    .A2(\sa30_sr[6] ),
    .ZN(_10582_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19488_ (.A1(\sa10_sr[6] ),
    .A2(_10582_),
    .Z(_10583_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19489_ (.A1(_10581_),
    .A2(_10583_),
    .Z(_10584_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _19490_ (.I(_10403_),
    .Z(_10585_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _19491_ (.I(_10431_),
    .Z(_10586_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _19492_ (.I(_10586_),
    .Z(_10587_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19493_ (.A1(_10587_),
    .A2(\text_in_r[126] ),
    .Z(_10588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19494_ (.A1(_10584_),
    .A2(_10585_),
    .B(_10588_),
    .ZN(_10589_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _19495_ (.A1(\u0.w[0][30] ),
    .A2(_10589_),
    .Z(_10590_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19496_ (.I(_10590_),
    .Z(_10591_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19497_ (.A1(_10559_),
    .A2(_10580_),
    .A3(_10591_),
    .ZN(_10592_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19498_ (.I(_10492_),
    .Z(_10593_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19499_ (.I(_10593_),
    .Z(_10594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19500_ (.A1(_10445_),
    .A2(net830),
    .ZN(_10595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19501_ (.I(_15683_),
    .ZN(_10596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19502_ (.A1(_15698_),
    .A2(_10596_),
    .ZN(_10597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19503_ (.A1(_10595_),
    .A2(_10597_),
    .Z(_10598_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19504_ (.A1(_10446_),
    .A2(_10509_),
    .A3(_10536_),
    .ZN(_10599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19505_ (.I(_10538_),
    .Z(_10600_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19506_ (.A1(_10594_),
    .A2(_10598_),
    .B(_10599_),
    .C(_10600_),
    .ZN(_10601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19507_ (.A1(_10494_),
    .A2(_15691_),
    .ZN(_10602_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19508_ (.I(_10503_),
    .Z(_10603_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19509_ (.A1(_10603_),
    .A2(_10602_),
    .Z(_10604_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19510_ (.I(_10538_),
    .Z(_10605_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19511_ (.A1(_10604_),
    .A2(_10605_),
    .ZN(_10606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19512_ (.A1(_15698_),
    .A2(_10498_),
    .ZN(_10607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19513_ (.I(_10607_),
    .ZN(_10608_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19514_ (.A1(_10565_),
    .A2(_10608_),
    .B(_10493_),
    .ZN(_10609_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19515_ (.I(_10555_),
    .Z(_10610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19516_ (.A1(_10606_),
    .A2(_10609_),
    .B(_10610_),
    .ZN(_10611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19517_ (.A1(_10601_),
    .A2(_10611_),
    .ZN(_10612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19518_ (.A1(net80),
    .A2(_10447_),
    .ZN(_10613_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19519_ (.I(_10603_),
    .Z(_10614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19520_ (.A1(_10440_),
    .A2(net597),
    .ZN(_10615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19521_ (.A1(_10613_),
    .A2(_10614_),
    .A3(_10615_),
    .ZN(_10616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19522_ (.A1(_15698_),
    .A2(_15680_),
    .ZN(_10617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19523_ (.I(_10617_),
    .ZN(_10618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19524_ (.A1(_10618_),
    .A2(_10493_),
    .B(_10573_),
    .ZN(_10619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19525_ (.A1(_10616_),
    .A2(_10619_),
    .ZN(_10620_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19526_ (.I(_15676_),
    .ZN(_10621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19527_ (.A1(_10445_),
    .A2(_10621_),
    .ZN(_10622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19528_ (.A1(_10622_),
    .A2(_10603_),
    .ZN(_10623_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19529_ (.A1(_10623_),
    .A2(_10573_),
    .Z(_10624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19530_ (.A1(_10445_),
    .A2(_15685_),
    .ZN(_10625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19531_ (.A1(_10617_),
    .A2(_10625_),
    .ZN(_10626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19532_ (.A1(_10626_),
    .A2(_10594_),
    .ZN(_10627_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19533_ (.I(_10556_),
    .Z(_10628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19534_ (.A1(_10624_),
    .A2(_10627_),
    .B(_10628_),
    .ZN(_10629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19535_ (.A1(_10620_),
    .A2(_10629_),
    .ZN(_10630_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19536_ (.I(_10590_),
    .ZN(_10631_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19537_ (.I(_10631_),
    .Z(_10632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19538_ (.A1(_10612_),
    .A2(_10630_),
    .A3(_10632_),
    .ZN(_10633_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19539_ (.I(\sa20_sr[7] ),
    .Z(_10634_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19540_ (.I(\sa30_sr[7] ),
    .Z(_10635_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19541_ (.A1(\sa10_sr[6] ),
    .A2(\sa00_sr[6] ),
    .Z(_10636_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19542_ (.A1(net46),
    .A2(_10636_),
    .Z(_10637_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _19543_ (.A1(net47),
    .A2(net68),
    .A3(_10637_),
    .Z(_10638_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _19544_ (.I(_10483_),
    .Z(_10639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19545_ (.I0(_10638_),
    .I1(\text_in_r[127] ),
    .S(_10639_),
    .Z(_10640_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _19546_ (.A1(\u0.w[0][31] ),
    .A2(_10640_),
    .ZN(_10641_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19547_ (.I(_10641_),
    .Z(_10642_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _19548_ (.I(_10642_),
    .ZN(_10643_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19549_ (.A1(_10592_),
    .A2(_10633_),
    .A3(_10643_),
    .ZN(_10644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19550_ (.A1(net601),
    .A2(_10440_),
    .ZN(_10645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19551_ (.A1(_10435_),
    .A2(_10439_),
    .A3(_15676_),
    .ZN(_10646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19552_ (.A1(_10566_),
    .A2(_10646_),
    .ZN(_10647_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19553_ (.I(_10647_),
    .ZN(_10648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19554_ (.A1(_10440_),
    .A2(_10621_),
    .ZN(_10649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19555_ (.A1(_10649_),
    .A2(_10603_),
    .Z(_10650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _19556_ (.A1(_10645_),
    .A2(_10648_),
    .B(_10650_),
    .C(_10605_),
    .ZN(_10651_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19557_ (.I(_10499_),
    .ZN(_10652_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _19558_ (.I(_10597_),
    .ZN(_10653_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19559_ (.I(_10593_),
    .Z(_10654_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19560_ (.A1(_10652_),
    .A2(_10653_),
    .B(_10654_),
    .ZN(_10655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19561_ (.I(_10623_),
    .ZN(_10656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19562_ (.A1(_15698_),
    .A2(_15675_),
    .ZN(_10657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19563_ (.A1(_10656_),
    .A2(_10657_),
    .ZN(_10658_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19564_ (.I(_10572_),
    .Z(_10659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19565_ (.A1(_10655_),
    .A2(_10658_),
    .B(_10659_),
    .ZN(_10660_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19566_ (.I(_10555_),
    .Z(_10661_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19567_ (.A1(_10651_),
    .A2(_10660_),
    .B(_10661_),
    .ZN(_10662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19568_ (.A1(_10595_),
    .A2(_10593_),
    .Z(_10663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19569_ (.A1(_10383_),
    .A2(net630),
    .ZN(_10664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19570_ (.A1(net827),
    .A2(_10384_),
    .A3(_10382_),
    .ZN(_10665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19571_ (.A1(_10665_),
    .A2(_10664_),
    .ZN(_15674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19572_ (.A1(net1262),
    .A2(net33),
    .ZN(_10666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19573_ (.A1(_10663_),
    .A2(_10666_),
    .ZN(_10667_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19574_ (.I(_10573_),
    .Z(_10668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19575_ (.A1(net599),
    .A2(net598),
    .ZN(_10669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19576_ (.A1(_10669_),
    .A2(_10614_),
    .A3(_10497_),
    .ZN(_10670_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19577_ (.A1(_10667_),
    .A2(_10668_),
    .A3(_10670_),
    .ZN(_10671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19578_ (.A1(_15691_),
    .A2(_10596_),
    .ZN(_10672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19579_ (.A1(_10607_),
    .A2(_10672_),
    .ZN(_10673_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19580_ (.I(_10572_),
    .Z(_10674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19581_ (.A1(_10673_),
    .A2(_10540_),
    .B(_10674_),
    .ZN(_10675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19582_ (.A1(net591),
    .A2(_10566_),
    .Z(_10676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19583_ (.A1(net32),
    .A2(net80),
    .A3(_15698_),
    .ZN(_10677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19584_ (.A1(_10676_),
    .A2(_10677_),
    .ZN(_10678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19585_ (.A1(_10678_),
    .A2(_10675_),
    .ZN(_10679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19586_ (.A1(_10671_),
    .A2(_10679_),
    .A3(_10579_),
    .ZN(_10680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19587_ (.A1(_10662_),
    .A2(_10680_),
    .A3(_10591_),
    .ZN(_10681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19588_ (.A1(_10615_),
    .A2(_10492_),
    .ZN(_10682_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19589_ (.A1(_10682_),
    .A2(_10538_),
    .Z(_10683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19590_ (.A1(net32),
    .A2(_15698_),
    .A3(net33),
    .ZN(_10684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19591_ (.A1(_10604_),
    .A2(_10684_),
    .ZN(_10685_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19592_ (.I(_10555_),
    .Z(_10686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19593_ (.A1(_10683_),
    .A2(_10685_),
    .B(_10686_),
    .ZN(_10687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19594_ (.A1(_10445_),
    .A2(net597),
    .ZN(_10688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19595_ (.A1(_10688_),
    .A2(_10566_),
    .Z(_10689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19596_ (.A1(_10689_),
    .A2(_10684_),
    .ZN(_10690_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19597_ (.I(_15689_),
    .ZN(_10691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19598_ (.A1(_10691_),
    .A2(_10440_),
    .ZN(_10692_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19599_ (.A1(_10692_),
    .A2(_10504_),
    .Z(_10693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19600_ (.A1(_10693_),
    .A2(net592),
    .ZN(_10694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19601_ (.A1(_10690_),
    .A2(_10694_),
    .A3(_10659_),
    .ZN(_10695_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19602_ (.I(_10590_),
    .Z(_10696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19603_ (.A1(_10687_),
    .A2(_10695_),
    .B(_10696_),
    .ZN(_10697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19604_ (.A1(_10567_),
    .A2(_10538_),
    .ZN(_10698_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19605_ (.A1(net32),
    .A2(_15691_),
    .ZN(_10699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19606_ (.A1(_10699_),
    .A2(_10593_),
    .Z(_10700_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19607_ (.A1(_10698_),
    .A2(_10700_),
    .ZN(_10701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19608_ (.A1(_10701_),
    .A2(_10616_),
    .ZN(_10702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19609_ (.A1(net36),
    .A2(_15691_),
    .ZN(_10703_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19610_ (.I(_10703_),
    .Z(_10704_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19611_ (.A1(_10684_),
    .A2(_10654_),
    .A3(_10704_),
    .ZN(_10705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19612_ (.A1(_10691_),
    .A2(_15691_),
    .ZN(_10706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19613_ (.A1(_10615_),
    .A2(_10706_),
    .A3(_10505_),
    .ZN(_10707_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19614_ (.A1(_10705_),
    .A2(_10659_),
    .A3(_10707_),
    .ZN(_10708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19615_ (.A1(_10702_),
    .A2(_10708_),
    .A3(_10610_),
    .ZN(_10709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19616_ (.A1(_10697_),
    .A2(_10709_),
    .B(_10643_),
    .ZN(_10710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19617_ (.A1(_10681_),
    .A2(_10710_),
    .ZN(_10711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19618_ (.A1(_10711_),
    .A2(_10644_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19619_ (.I(_10682_),
    .ZN(_10712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19620_ (.A1(_10613_),
    .A2(_10712_),
    .ZN(_10713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19621_ (.A1(_10623_),
    .A2(_10533_),
    .Z(_10714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19622_ (.A1(_10713_),
    .A2(_10714_),
    .B(_10628_),
    .ZN(_10715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19623_ (.A1(_10706_),
    .A2(_10566_),
    .Z(_10716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19624_ (.I(_15677_),
    .ZN(_10717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19625_ (.A1(_15698_),
    .A2(_10717_),
    .ZN(_10718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19626_ (.A1(_10716_),
    .A2(_10718_),
    .B(_10605_),
    .ZN(_10719_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19627_ (.A1(_10677_),
    .A2(_10505_),
    .A3(_10646_),
    .ZN(_10720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19628_ (.A1(_10719_),
    .A2(_10720_),
    .ZN(_10721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19629_ (.A1(_10715_),
    .A2(_10721_),
    .B(_10696_),
    .ZN(_10722_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19630_ (.I(_10497_),
    .ZN(_10723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19631_ (.A1(_10723_),
    .A2(_10509_),
    .ZN(_10724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19632_ (.A1(_10724_),
    .A2(_10567_),
    .Z(_10725_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19633_ (.A1(_10652_),
    .A2(_10537_),
    .B(_10505_),
    .ZN(_10726_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19634_ (.A1(_10725_),
    .A2(_10668_),
    .A3(_10726_),
    .ZN(_10727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19635_ (.A1(_10663_),
    .A2(_10657_),
    .ZN(_10728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19636_ (.A1(net611),
    .A2(_10440_),
    .ZN(_10729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19637_ (.A1(_10604_),
    .A2(_10729_),
    .ZN(_10730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19638_ (.A1(_10728_),
    .A2(_10730_),
    .A3(_10564_),
    .ZN(_10731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19639_ (.A1(_10727_),
    .A2(_10731_),
    .A3(_10579_),
    .ZN(_10732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19640_ (.A1(_10722_),
    .A2(_10732_),
    .B(_10643_),
    .ZN(_10733_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19641_ (.A1(_10613_),
    .A2(_10540_),
    .A3(_10684_),
    .ZN(_10734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19642_ (.A1(_10689_),
    .A2(_10657_),
    .B(_10555_),
    .ZN(_10735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19643_ (.A1(_10734_),
    .A2(_10735_),
    .ZN(_10736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19644_ (.A1(_10663_),
    .A2(_10645_),
    .ZN(_10737_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19645_ (.A1(_10737_),
    .A2(_10730_),
    .A3(_10610_),
    .ZN(_10738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19646_ (.A1(_10736_),
    .A2(_10738_),
    .B(_10564_),
    .ZN(_10739_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19647_ (.A1(_10556_),
    .A2(_15699_),
    .A3(_10493_),
    .Z(_10740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19648_ (.A1(_10613_),
    .A2(_10576_),
    .ZN(_10741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19649_ (.A1(_10740_),
    .A2(_10564_),
    .A3(_10741_),
    .ZN(_10742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19650_ (.I(_10742_),
    .ZN(_10743_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19651_ (.A1(_10739_),
    .A2(_10743_),
    .B(_10591_),
    .ZN(_10744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19652_ (.A1(_10733_),
    .A2(_10744_),
    .ZN(_10745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19653_ (.A1(_10603_),
    .A2(_15698_),
    .Z(_10746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19654_ (.A1(_10746_),
    .A2(_10669_),
    .ZN(_10747_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19655_ (.A1(_10747_),
    .A2(_10533_),
    .Z(_10748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19656_ (.A1(_10446_),
    .A2(_10566_),
    .Z(_10749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19657_ (.A1(_10749_),
    .A2(_10666_),
    .ZN(_10750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19658_ (.A1(_10748_),
    .A2(_10750_),
    .ZN(_10751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19659_ (.A1(_10602_),
    .A2(_10593_),
    .ZN(_10752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19660_ (.A1(_10752_),
    .A2(_10723_),
    .Z(_10753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19661_ (.A1(_10656_),
    .A2(_10615_),
    .ZN(_10754_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19662_ (.I(_10573_),
    .Z(_10755_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19663_ (.A1(_10753_),
    .A2(_10754_),
    .A3(_10755_),
    .ZN(_10756_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19664_ (.A1(_10751_),
    .A2(_10756_),
    .A3(_10579_),
    .ZN(_10757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19665_ (.A1(_10650_),
    .A2(_10706_),
    .ZN(_10758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19666_ (.A1(_10758_),
    .A2(_10533_),
    .Z(_10759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19667_ (.A1(_10759_),
    .A2(_10496_),
    .ZN(_10760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19668_ (.A1(_10645_),
    .A2(_10603_),
    .ZN(_10761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19669_ (.A1(_10761_),
    .A2(_10704_),
    .Z(_10762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _19670_ (.A1(_10618_),
    .A2(_10493_),
    .B(_10538_),
    .ZN(_10763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19671_ (.A1(_10762_),
    .A2(_10763_),
    .B(_10628_),
    .ZN(_10764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19672_ (.A1(_10760_),
    .A2(_10764_),
    .ZN(_10765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19673_ (.A1(_10757_),
    .A2(_10765_),
    .A3(_10591_),
    .ZN(_10766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19674_ (.I(net591),
    .ZN(_10767_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19675_ (.A1(_10767_),
    .A2(_10618_),
    .B(_10505_),
    .ZN(_10768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19676_ (.A1(_10500_),
    .A2(_10654_),
    .ZN(_10769_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19677_ (.A1(_10768_),
    .A2(_10755_),
    .A3(_10769_),
    .ZN(_10770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19678_ (.A1(net32),
    .A2(net80),
    .ZN(_10771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19679_ (.A1(_10771_),
    .A2(_10688_),
    .ZN(_10772_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _19680_ (.I(_10504_),
    .Z(_10773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19681_ (.A1(_10772_),
    .A2(_10773_),
    .ZN(_10774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19682_ (.A1(_10536_),
    .A2(_10566_),
    .Z(_10775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19683_ (.A1(_10775_),
    .A2(_10688_),
    .ZN(_10776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19684_ (.A1(_10774_),
    .A2(_10776_),
    .A3(_10600_),
    .ZN(_10777_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19685_ (.A1(_10770_),
    .A2(_10777_),
    .A3(_10661_),
    .ZN(_10778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19686_ (.A1(_10693_),
    .A2(_10704_),
    .ZN(_10779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19687_ (.A1(_10771_),
    .A2(_15691_),
    .A3(_10493_),
    .ZN(_10780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19688_ (.A1(_10779_),
    .A2(_10780_),
    .A3(_10659_),
    .ZN(_10781_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19689_ (.A1(_15691_),
    .A2(_15680_),
    .Z(_10782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _19690_ (.I(_10572_),
    .Z(_10783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19691_ (.A1(_10782_),
    .A2(_10493_),
    .B(_10783_),
    .ZN(_10784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19692_ (.A1(_10720_),
    .A2(_10784_),
    .ZN(_10785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19693_ (.A1(_10781_),
    .A2(_10785_),
    .A3(_10557_),
    .ZN(_10786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19694_ (.A1(_10778_),
    .A2(_10786_),
    .A3(_10632_),
    .ZN(_10787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19695_ (.A1(_10766_),
    .A2(_10787_),
    .A3(_10643_),
    .ZN(_10788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19696_ (.A1(_10745_),
    .A2(_10788_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19697_ (.A1(_10688_),
    .A2(_10495_),
    .ZN(_10789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19698_ (.A1(_10789_),
    .A2(_10614_),
    .A3(_10704_),
    .ZN(_10790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19699_ (.A1(_10790_),
    .A2(_10605_),
    .A3(_10599_),
    .ZN(_10791_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19700_ (.A1(_10669_),
    .A2(_10446_),
    .A3(_10504_),
    .ZN(_10792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19701_ (.A1(_10692_),
    .A2(_10602_),
    .A3(_10593_),
    .ZN(_10793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19702_ (.A1(_10792_),
    .A2(_10793_),
    .ZN(_10794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19703_ (.A1(_10794_),
    .A2(_10659_),
    .ZN(_10795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19704_ (.A1(_10791_),
    .A2(_10795_),
    .A3(_10610_),
    .ZN(_10796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19705_ (.A1(_10684_),
    .A2(_10509_),
    .B(_10572_),
    .ZN(_10797_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19706_ (.A1(_10677_),
    .A2(_10614_),
    .A3(_10706_),
    .ZN(_10798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19707_ (.A1(_10797_),
    .A2(_10798_),
    .ZN(_10799_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19708_ (.A1(_10647_),
    .A2(_10699_),
    .ZN(_10800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19709_ (.A1(_10507_),
    .A2(_10603_),
    .ZN(_10801_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19710_ (.I(_10595_),
    .ZN(_10802_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19711_ (.A1(_10801_),
    .A2(_10802_),
    .ZN(_10803_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19712_ (.A1(_10800_),
    .A2(_10803_),
    .B(_10783_),
    .ZN(_10804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19713_ (.A1(_10799_),
    .A2(_10804_),
    .ZN(_10805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19714_ (.A1(_10805_),
    .A2(_10557_),
    .ZN(_10806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19715_ (.A1(_10796_),
    .A2(_10806_),
    .A3(_10591_),
    .ZN(_10807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19716_ (.A1(_10443_),
    .A2(net603),
    .A3(_15689_),
    .ZN(_10808_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19717_ (.A1(_10595_),
    .A2(_10566_),
    .A3(_10808_),
    .ZN(_10809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19718_ (.A1(_10809_),
    .A2(_10572_),
    .ZN(_10810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19719_ (.A1(_10625_),
    .A2(_10504_),
    .ZN(_10811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19720_ (.A1(_10811_),
    .A2(_10699_),
    .ZN(_10812_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19721_ (.A1(_10810_),
    .A2(_10812_),
    .ZN(_10813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19722_ (.A1(_10688_),
    .A2(_10593_),
    .A3(_10561_),
    .ZN(_10814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19723_ (.A1(net591),
    .A2(_10536_),
    .A3(_10504_),
    .ZN(_10815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19724_ (.A1(_10814_),
    .A2(_10815_),
    .B(_10573_),
    .ZN(_10816_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19725_ (.A1(_10813_),
    .A2(_10816_),
    .B(_10628_),
    .ZN(_10817_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19726_ (.A1(_10626_),
    .A2(_10509_),
    .B(_10572_),
    .ZN(_10818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19727_ (.A1(_10495_),
    .A2(_10603_),
    .Z(_10819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19728_ (.A1(_10819_),
    .A2(_10703_),
    .ZN(_10820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19729_ (.A1(_10818_),
    .A2(_10820_),
    .ZN(_10821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19730_ (.A1(_10625_),
    .A2(_10808_),
    .ZN(_10822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19731_ (.A1(_10822_),
    .A2(_10509_),
    .ZN(_10823_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19732_ (.A1(_10688_),
    .A2(_10495_),
    .A3(_10614_),
    .ZN(_10824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19733_ (.A1(_10823_),
    .A2(_10824_),
    .A3(_10573_),
    .ZN(_10825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19734_ (.A1(_10821_),
    .A2(_10825_),
    .A3(_10555_),
    .ZN(_10826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19735_ (.A1(_10817_),
    .A2(_10826_),
    .ZN(_10827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19736_ (.A1(_10827_),
    .A2(_10632_),
    .ZN(_10828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19737_ (.A1(_10807_),
    .A2(_10828_),
    .ZN(_10829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19738_ (.A1(_10829_),
    .A2(_10642_),
    .ZN(_10830_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19739_ (.A1(_10749_),
    .A2(_10607_),
    .Z(_10831_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19740_ (.A1(_10672_),
    .A2(_10614_),
    .A3(net609),
    .Z(_10832_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19741_ (.A1(_10831_),
    .A2(_10832_),
    .B(_10668_),
    .ZN(_10833_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19742_ (.A1(_10666_),
    .A2(_10446_),
    .A3(_10504_),
    .Z(_10834_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19743_ (.A1(_10834_),
    .A2(_10783_),
    .ZN(_10835_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19744_ (.A1(_10505_),
    .A2(_15699_),
    .Z(_10836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19745_ (.A1(_10835_),
    .A2(_10836_),
    .ZN(_10837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19746_ (.A1(_10833_),
    .A2(_10837_),
    .A3(_10661_),
    .ZN(_10838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19747_ (.A1(_10448_),
    .A2(_10650_),
    .ZN(_10839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19748_ (.A1(_15696_),
    .A2(_10654_),
    .B(_10783_),
    .ZN(_10840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19749_ (.A1(_10839_),
    .A2(_10840_),
    .B(_10686_),
    .ZN(_10841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19750_ (.A1(_10729_),
    .A2(_10603_),
    .Z(_10842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19751_ (.A1(_10842_),
    .A2(_10688_),
    .ZN(_10843_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19752_ (.A1(_10843_),
    .A2(_10755_),
    .A3(_10599_),
    .ZN(_10844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19753_ (.A1(_10841_),
    .A2(_10844_),
    .B(_10696_),
    .ZN(_10845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19754_ (.A1(_10838_),
    .A2(_10845_),
    .ZN(_10846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19755_ (.A1(_10746_),
    .A2(_10771_),
    .ZN(_10847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19756_ (.A1(_10847_),
    .A2(_10783_),
    .Z(_10848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19757_ (.A1(_10717_),
    .A2(_10494_),
    .Z(_10849_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19758_ (.A1(_10493_),
    .A2(_15698_),
    .A3(_10849_),
    .Z(_10850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19759_ (.A1(_10848_),
    .A2(_10741_),
    .A3(_10850_),
    .ZN(_10851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19760_ (.A1(_10652_),
    .A2(_10593_),
    .ZN(_10852_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19761_ (.A1(_10852_),
    .A2(_10538_),
    .Z(_10853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19762_ (.A1(_10656_),
    .A2(_10495_),
    .ZN(_10854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19763_ (.A1(_10854_),
    .A2(_10853_),
    .B(_10686_),
    .ZN(_10855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19764_ (.A1(_10851_),
    .A2(_10855_),
    .ZN(_10856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19765_ (.A1(_15703_),
    .A2(_10654_),
    .B(_10533_),
    .ZN(_10857_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19766_ (.A1(_10857_),
    .A2(_10792_),
    .B(_10628_),
    .ZN(_10858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19767_ (.A1(_10684_),
    .A2(_10654_),
    .ZN(_10859_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19768_ (.A1(_10509_),
    .A2(_15694_),
    .Z(_10860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19769_ (.A1(_10859_),
    .A2(_10600_),
    .A3(_10860_),
    .ZN(_10861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19770_ (.A1(_10858_),
    .A2(_10861_),
    .ZN(_10862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19771_ (.A1(_10856_),
    .A2(_10862_),
    .A3(_10591_),
    .ZN(_10863_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19772_ (.A1(_10846_),
    .A2(_10863_),
    .A3(_10643_),
    .ZN(_10864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19773_ (.A1(_10830_),
    .A2(_10864_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19774_ (.A1(_10669_),
    .A2(_10595_),
    .ZN(_10865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19775_ (.A1(_10865_),
    .A2(_10538_),
    .Z(_10866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19776_ (.A1(_10603_),
    .A2(_15691_),
    .Z(_10867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19777_ (.I(_10867_),
    .ZN(_10868_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19778_ (.A1(_10866_),
    .A2(_10868_),
    .B(_10590_),
    .ZN(_10869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19779_ (.A1(_10648_),
    .A2(_10561_),
    .ZN(_10870_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19780_ (.A1(_10779_),
    .A2(_10870_),
    .A3(_10755_),
    .ZN(_10871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19781_ (.A1(_10869_),
    .A2(_10871_),
    .B(_10557_),
    .ZN(_10872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19782_ (.A1(_10663_),
    .A2(_10669_),
    .ZN(_10873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19783_ (.A1(_10656_),
    .A2(_10729_),
    .ZN(_10874_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19784_ (.A1(_10873_),
    .A2(_10564_),
    .A3(_10874_),
    .ZN(_10875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19785_ (.A1(_10689_),
    .A2(_10729_),
    .ZN(_10876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19786_ (.I(_10650_),
    .ZN(_10877_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19787_ (.A1(_10876_),
    .A2(_10668_),
    .A3(_10877_),
    .ZN(_10878_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19788_ (.A1(_10696_),
    .A2(_10878_),
    .A3(_10875_),
    .ZN(_10879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19789_ (.A1(_10879_),
    .A2(_10872_),
    .B(_10642_),
    .ZN(_10880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19790_ (.A1(_10497_),
    .A2(_10672_),
    .Z(_10881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19791_ (.A1(_10842_),
    .A2(_10881_),
    .ZN(_10882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19792_ (.A1(_10882_),
    .A2(_10605_),
    .ZN(_10883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19793_ (.A1(_10775_),
    .A2(_10704_),
    .A3(_10688_),
    .Z(_10884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19794_ (.A1(_10883_),
    .A2(_10884_),
    .ZN(_10885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19795_ (.A1(_10676_),
    .A2(_10597_),
    .ZN(_10886_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19796_ (.A1(_10886_),
    .A2(_10674_),
    .A3(_10670_),
    .Z(_10887_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19797_ (.A1(_10885_),
    .A2(_10887_),
    .B(_10632_),
    .ZN(_10888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19798_ (.A1(_10706_),
    .A2(_10819_),
    .B(_10800_),
    .ZN(_10889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19799_ (.A1(_10889_),
    .A2(_10564_),
    .ZN(_10890_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19800_ (.A1(_10881_),
    .A2(_10614_),
    .Z(_10891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19801_ (.A1(_10867_),
    .A2(_10498_),
    .B(_10533_),
    .ZN(_10892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19802_ (.A1(_10746_),
    .A2(_10621_),
    .Z(_10893_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19803_ (.I(_10893_),
    .ZN(_10894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19804_ (.A1(_10891_),
    .A2(_10892_),
    .A3(_10894_),
    .ZN(_10895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19805_ (.A1(_10890_),
    .A2(_10895_),
    .A3(_10591_),
    .ZN(_10896_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19806_ (.A1(_10888_),
    .A2(_10896_),
    .A3(_10579_),
    .ZN(_10897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19807_ (.A1(_10880_),
    .A2(_10897_),
    .ZN(_10898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19808_ (.A1(_10576_),
    .A2(_10446_),
    .Z(_10899_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19809_ (.A1(_10899_),
    .A2(_10893_),
    .B(_10555_),
    .ZN(_10900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19810_ (.A1(_10767_),
    .A2(_10593_),
    .Z(_10901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _19811_ (.A1(_10901_),
    .A2(_10628_),
    .B1(_10773_),
    .B2(_10565_),
    .ZN(_10902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19812_ (.A1(_10900_),
    .A2(_10902_),
    .ZN(_10903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19813_ (.A1(_10903_),
    .A2(_10668_),
    .ZN(_10904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19814_ (.I(_10625_),
    .ZN(_10905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19815_ (.A1(_10905_),
    .A2(_10504_),
    .ZN(_10906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19816_ (.A1(_10906_),
    .A2(_10556_),
    .Z(_10907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19817_ (.A1(_10907_),
    .A2(_10814_),
    .B(_10659_),
    .ZN(_10908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19818_ (.A1(_10712_),
    .A2(net591),
    .ZN(_10909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19819_ (.A1(_15691_),
    .A2(_10849_),
    .ZN(_10910_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19820_ (.A1(_10692_),
    .A2(_10910_),
    .A3(_10505_),
    .ZN(_10911_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19821_ (.A1(_10909_),
    .A2(_10911_),
    .A3(_10610_),
    .ZN(_10912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19822_ (.A1(_10908_),
    .A2(_10912_),
    .B(_10631_),
    .ZN(_10913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19823_ (.A1(_10904_),
    .A2(_10913_),
    .ZN(_10914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19824_ (.A1(_10562_),
    .A2(_10910_),
    .ZN(_10915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19825_ (.A1(_10741_),
    .A2(_10915_),
    .A3(_10600_),
    .ZN(_10916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19826_ (.I(_10809_),
    .ZN(_10917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19827_ (.A1(_10917_),
    .A2(_10659_),
    .B(_10628_),
    .ZN(_10918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19828_ (.A1(_10916_),
    .A2(_10918_),
    .B(_10696_),
    .ZN(_10919_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19829_ (.A1(_10906_),
    .A2(_10573_),
    .Z(_10920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19830_ (.A1(_10676_),
    .A2(_10692_),
    .ZN(_10921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19831_ (.A1(_10746_),
    .A2(net33),
    .ZN(_10922_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19832_ (.A1(_10920_),
    .A2(_10921_),
    .A3(_10922_),
    .ZN(_10923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19833_ (.A1(_10750_),
    .A2(_10600_),
    .A3(_10506_),
    .ZN(_10924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19834_ (.A1(_10923_),
    .A2(_10924_),
    .A3(_10579_),
    .ZN(_10925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19835_ (.A1(_10919_),
    .A2(_10925_),
    .ZN(_10926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19836_ (.A1(_10914_),
    .A2(_10926_),
    .A3(_10642_),
    .ZN(_10927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19837_ (.A1(_10898_),
    .A2(_10927_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19838_ (.A1(_10699_),
    .A2(_10594_),
    .ZN(_10928_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _19839_ (.A1(_10668_),
    .A2(_10730_),
    .A3(_10852_),
    .A4(_10928_),
    .ZN(_10929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19840_ (.A1(_10663_),
    .A2(_10692_),
    .ZN(_10930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19841_ (.A1(_10746_),
    .A2(_10674_),
    .ZN(_10931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19842_ (.A1(_10930_),
    .A2(_10931_),
    .B(_10557_),
    .ZN(_10932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19843_ (.A1(_10929_),
    .A2(_10932_),
    .ZN(_10933_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19844_ (.A1(_10537_),
    .A2(_10752_),
    .Z(_10934_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19845_ (.A1(_10616_),
    .A2(_10934_),
    .A3(_10564_),
    .ZN(_10935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19846_ (.A1(_10718_),
    .A2(_10509_),
    .ZN(_10936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19847_ (.A1(_10936_),
    .A2(_10783_),
    .Z(_10937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19848_ (.A1(_10677_),
    .A2(_10540_),
    .ZN(_10938_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19849_ (.A1(_10937_),
    .A2(_10938_),
    .B(_10610_),
    .ZN(_10939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19850_ (.A1(_10939_),
    .A2(_10935_),
    .ZN(_10940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19851_ (.A1(_10940_),
    .A2(_10933_),
    .A3(_10632_),
    .ZN(_10941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19852_ (.A1(_10802_),
    .A2(_10593_),
    .ZN(_10942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19853_ (.A1(_10942_),
    .A2(_10783_),
    .Z(_10943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19854_ (.A1(_10562_),
    .A2(_10703_),
    .ZN(_10944_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19855_ (.A1(_10704_),
    .A2(_10614_),
    .Z(_10945_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19856_ (.A1(_10943_),
    .A2(_10944_),
    .A3(_10945_),
    .ZN(_10946_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19857_ (.I(_15687_),
    .ZN(_10947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19858_ (.A1(_10947_),
    .A2(_10654_),
    .B(_10783_),
    .ZN(_10948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19859_ (.A1(_10536_),
    .A2(_10773_),
    .ZN(_10949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19860_ (.A1(_10949_),
    .A2(_10948_),
    .B(_10686_),
    .ZN(_10950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19861_ (.A1(_10946_),
    .A2(_10950_),
    .B(_10631_),
    .ZN(_10951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19862_ (.A1(_10729_),
    .A2(_10566_),
    .ZN(_10952_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19863_ (.I(_10669_),
    .ZN(_10953_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19864_ (.A1(_10952_),
    .A2(_10953_),
    .ZN(_10954_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19865_ (.I(_10954_),
    .ZN(_10955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19866_ (.A1(_10562_),
    .A2(_10595_),
    .ZN(_10956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19867_ (.A1(_10955_),
    .A2(_10956_),
    .A3(_10755_),
    .ZN(_10957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19868_ (.A1(_10609_),
    .A2(_10600_),
    .A3(_10670_),
    .ZN(_10958_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19869_ (.A1(_10957_),
    .A2(_10958_),
    .A3(_10661_),
    .ZN(_10959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19870_ (.A1(_10959_),
    .A2(_10951_),
    .ZN(_10960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19871_ (.A1(_10960_),
    .A2(_10642_),
    .A3(_10941_),
    .ZN(_10961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19872_ (.A1(_10716_),
    .A2(_10649_),
    .ZN(_10962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19873_ (.A1(_10563_),
    .A2(_10564_),
    .A3(_10962_),
    .ZN(_10963_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19874_ (.A1(_10509_),
    .A2(_10536_),
    .ZN(_10964_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19875_ (.A1(_10964_),
    .A2(_10905_),
    .ZN(_10965_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19876_ (.A1(_10763_),
    .A2(_10965_),
    .B(_10686_),
    .ZN(_10966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19877_ (.A1(_10963_),
    .A2(_10966_),
    .B(_10631_),
    .ZN(_10967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19878_ (.A1(_10842_),
    .A2(_10448_),
    .ZN(_10968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19879_ (.A1(_10968_),
    .A2(_10755_),
    .A3(_10793_),
    .ZN(_10969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19880_ (.A1(_10645_),
    .A2(_10499_),
    .ZN(_10970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19881_ (.A1(_10970_),
    .A2(_10773_),
    .B(_10674_),
    .ZN(_10971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19882_ (.A1(_10496_),
    .A2(_10971_),
    .ZN(_10972_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19883_ (.A1(_10969_),
    .A2(_10972_),
    .A3(_10661_),
    .ZN(_10973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19884_ (.A1(_10967_),
    .A2(_10973_),
    .B(_10642_),
    .ZN(_10974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19885_ (.A1(_10835_),
    .A2(_10737_),
    .ZN(_10975_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19886_ (.A1(_10446_),
    .A2(_10614_),
    .A3(_10607_),
    .Z(_10976_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19887_ (.A1(_10976_),
    .A2(_10954_),
    .B(_10755_),
    .ZN(_10977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19888_ (.A1(_10975_),
    .A2(_10977_),
    .A3(_10661_),
    .ZN(_10978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19889_ (.I(_10761_),
    .ZN(_10979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19890_ (.A1(_10979_),
    .A2(_10688_),
    .ZN(_10980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19891_ (.A1(_10689_),
    .A2(_10657_),
    .ZN(_10981_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19892_ (.A1(_10980_),
    .A2(_10600_),
    .A3(_10981_),
    .ZN(_10982_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19893_ (.A1(_10562_),
    .A2(_10533_),
    .A3(_10565_),
    .Z(_10983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19894_ (.A1(_10982_),
    .A2(_10557_),
    .A3(_10983_),
    .ZN(_10984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19895_ (.A1(_10978_),
    .A2(_10632_),
    .A3(_10984_),
    .ZN(_10985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19896_ (.A1(_10974_),
    .A2(_10985_),
    .ZN(_10986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19897_ (.A1(_10986_),
    .A2(_10961_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19898_ (.A1(net826),
    .A2(_10575_),
    .ZN(_10987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19899_ (.A1(_10712_),
    .A2(_10771_),
    .ZN(_10988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19900_ (.A1(_10988_),
    .A2(_10674_),
    .ZN(_10989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19901_ (.A1(_10987_),
    .A2(_10540_),
    .B(_10989_),
    .ZN(_10990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19902_ (.A1(_10505_),
    .A2(net1262),
    .ZN(_10991_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19903_ (.A1(_10955_),
    .A2(_10605_),
    .A3(_10991_),
    .Z(_10992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19904_ (.A1(_10990_),
    .A2(_10992_),
    .B(_10579_),
    .ZN(_10993_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19905_ (.A1(_10936_),
    .A2(_10447_),
    .ZN(_10994_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19906_ (.A1(_10994_),
    .A2(_10964_),
    .B(_10674_),
    .ZN(_10995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19907_ (.A1(_10808_),
    .A2(_10493_),
    .ZN(_10996_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19908_ (.A1(_10623_),
    .A2(_10608_),
    .B(_10605_),
    .C(_10996_),
    .ZN(_10997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19909_ (.A1(_10995_),
    .A2(_10997_),
    .ZN(_10998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19910_ (.A1(_10998_),
    .A2(_10661_),
    .B(_10632_),
    .ZN(_10999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19911_ (.A1(_10993_),
    .A2(_10999_),
    .ZN(_11000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _19912_ (.A1(_10746_),
    .A2(net33),
    .B(_10573_),
    .ZN(_11001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19913_ (.I(_10676_),
    .ZN(_11002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19914_ (.A1(_11001_),
    .A2(_11002_),
    .A3(_10906_),
    .ZN(_11003_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19915_ (.A1(_10752_),
    .A2(_10573_),
    .Z(_11004_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19916_ (.A1(_11004_),
    .A2(_10747_),
    .B(_10628_),
    .ZN(_11005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19917_ (.A1(_11003_),
    .A2(_11005_),
    .B(_10696_),
    .ZN(_11006_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19918_ (.A1(_10561_),
    .A2(_10492_),
    .Z(_11007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19919_ (.A1(_10448_),
    .A2(_11007_),
    .ZN(_11008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19920_ (.A1(_10540_),
    .A2(_15680_),
    .ZN(_11009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19921_ (.A1(_10574_),
    .A2(_11008_),
    .A3(_11009_),
    .ZN(_11010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19922_ (.A1(_10693_),
    .A2(_10602_),
    .ZN(_11011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19923_ (.A1(_10701_),
    .A2(_11011_),
    .ZN(_11012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19924_ (.A1(_11010_),
    .A2(_11012_),
    .A3(_10579_),
    .ZN(_11013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19925_ (.A1(_11006_),
    .A2(_11013_),
    .B(_10642_),
    .ZN(_11014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19926_ (.A1(_11000_),
    .A2(_11014_),
    .ZN(_11015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19927_ (.I(net826),
    .ZN(_11016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19928_ (.A1(_10910_),
    .A2(_10773_),
    .ZN(_11017_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19929_ (.A1(_11016_),
    .A2(_10859_),
    .B(_10600_),
    .C(_11017_),
    .ZN(_11018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19930_ (.I(_10693_),
    .ZN(_11019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19931_ (.A1(_10763_),
    .A2(_11019_),
    .B(_10686_),
    .ZN(_11020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19932_ (.A1(_11018_),
    .A2(_11020_),
    .ZN(_11021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19933_ (.A1(_10656_),
    .A2(_10575_),
    .ZN(_11022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19934_ (.A1(_10648_),
    .A2(_10692_),
    .ZN(_11023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19935_ (.A1(_11022_),
    .A2(_11023_),
    .A3(_10755_),
    .ZN(_11024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19936_ (.A1(net826),
    .A2(_10594_),
    .ZN(_11025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19937_ (.A1(_10596_),
    .A2(_10773_),
    .B(_10783_),
    .ZN(_11026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19938_ (.A1(_11025_),
    .A2(_11026_),
    .ZN(_11027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19939_ (.A1(_11024_),
    .A2(_11027_),
    .A3(_10610_),
    .ZN(_11028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19940_ (.A1(_11021_),
    .A2(_11028_),
    .A3(_10591_),
    .ZN(_11029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19941_ (.A1(net80),
    .A2(_10505_),
    .B(_10783_),
    .ZN(_11030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19942_ (.A1(_11030_),
    .A2(_10667_),
    .B(_10686_),
    .ZN(_11031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19943_ (.A1(_10656_),
    .A2(_10684_),
    .ZN(_11032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19944_ (.A1(_11007_),
    .A2(_10704_),
    .ZN(_11033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19945_ (.A1(_11032_),
    .A2(_11033_),
    .A3(_10659_),
    .ZN(_11034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19946_ (.A1(_11031_),
    .A2(_11034_),
    .B(_10696_),
    .ZN(_11035_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19947_ (.A1(_10613_),
    .A2(_10594_),
    .A3(_10692_),
    .ZN(_11036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19948_ (.A1(_10653_),
    .A2(_10773_),
    .B(_10533_),
    .ZN(_11037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19949_ (.A1(_11036_),
    .A2(_11037_),
    .B(_10628_),
    .ZN(_11038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19950_ (.A1(_10616_),
    .A2(_10619_),
    .A3(_10942_),
    .ZN(_11039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19951_ (.A1(_11038_),
    .A2(_11039_),
    .ZN(_11040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19952_ (.A1(_11035_),
    .A2(_11040_),
    .ZN(_11041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19953_ (.A1(_11029_),
    .A2(_11041_),
    .A3(_10642_),
    .ZN(_11042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19954_ (.A1(_11015_),
    .A2(_11042_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19955_ (.A1(_11007_),
    .A2(_10706_),
    .ZN(_11043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19956_ (.A1(_11043_),
    .A2(_10847_),
    .A3(_10569_),
    .ZN(_11044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19957_ (.A1(_11044_),
    .A2(_10605_),
    .Z(_11045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19958_ (.A1(_10626_),
    .A2(_10801_),
    .Z(_11046_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19959_ (.A1(_11046_),
    .A2(_10539_),
    .A3(_10942_),
    .Z(_11047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19960_ (.A1(_11045_),
    .A2(_11047_),
    .B(_10661_),
    .ZN(_11048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19961_ (.A1(_10508_),
    .A2(_10614_),
    .ZN(_11049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19962_ (.A1(_10852_),
    .A2(_11049_),
    .Z(_11050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19963_ (.A1(_11050_),
    .A2(_10920_),
    .B(_10686_),
    .ZN(_11051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19964_ (.A1(_10842_),
    .A2(_10669_),
    .ZN(_11052_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19965_ (.A1(_15692_),
    .A2(_15701_),
    .B(_10654_),
    .ZN(_11053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19966_ (.A1(_11052_),
    .A2(_10564_),
    .A3(_11053_),
    .ZN(_11054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19967_ (.A1(_11051_),
    .A2(_11054_),
    .B(_10696_),
    .ZN(_11055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19968_ (.A1(_11048_),
    .A2(_11055_),
    .ZN(_11056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19969_ (.A1(_10979_),
    .A2(_10669_),
    .ZN(_11057_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19970_ (.A1(_10653_),
    .A2(_10654_),
    .B(_10533_),
    .ZN(_11058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19971_ (.A1(_11057_),
    .A2(_11058_),
    .B(_10628_),
    .ZN(_11059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19972_ (.A1(_10775_),
    .A2(_10910_),
    .ZN(_11060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19973_ (.A1(_11001_),
    .A2(_10670_),
    .A3(_11060_),
    .ZN(_11061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19974_ (.A1(_11059_),
    .A2(_11061_),
    .B(_10632_),
    .ZN(_11062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19975_ (.A1(_10684_),
    .A2(_10594_),
    .A3(_10622_),
    .ZN(_11063_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19976_ (.A1(_11063_),
    .A2(_10668_),
    .A3(_10860_),
    .ZN(_11064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19977_ (.A1(_10684_),
    .A2(_10773_),
    .A3(_10704_),
    .ZN(_11065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19978_ (.A1(_10718_),
    .A2(_10646_),
    .A3(_10654_),
    .ZN(_11066_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19979_ (.A1(_11065_),
    .A2(_11066_),
    .A3(_10564_),
    .ZN(_11067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19980_ (.A1(_11064_),
    .A2(_11067_),
    .A3(_10579_),
    .ZN(_11068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19981_ (.A1(_11062_),
    .A2(_11068_),
    .ZN(_11069_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19982_ (.A1(_11056_),
    .A2(_11069_),
    .A3(_10643_),
    .ZN(_11070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19983_ (.I(_10576_),
    .ZN(_11071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19984_ (.A1(_10944_),
    .A2(_11071_),
    .ZN(_11072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19985_ (.A1(_11072_),
    .A2(_10674_),
    .ZN(_11073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19986_ (.A1(_10790_),
    .A2(_10605_),
    .ZN(_11074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19987_ (.A1(_11073_),
    .A2(_11074_),
    .ZN(_11075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19988_ (.A1(_11075_),
    .A2(_10661_),
    .ZN(_11076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19989_ (.A1(_10693_),
    .A2(_10646_),
    .ZN(_11077_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19990_ (.A1(_11077_),
    .A2(_10755_),
    .A3(_10724_),
    .ZN(_11078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19991_ (.I(_15693_),
    .ZN(_11079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19992_ (.A1(_11079_),
    .A2(_10773_),
    .B(_10674_),
    .ZN(_11080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19993_ (.A1(_11080_),
    .A2(_11033_),
    .ZN(_11081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19994_ (.A1(_11078_),
    .A2(_11081_),
    .A3(_10557_),
    .ZN(_11082_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19995_ (.A1(_11076_),
    .A2(_11082_),
    .A3(_10591_),
    .ZN(_11083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19996_ (.A1(_10690_),
    .A2(_10755_),
    .A3(_10761_),
    .ZN(_11084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19997_ (.A1(_10811_),
    .A2(_10647_),
    .ZN(_11085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19998_ (.A1(_11001_),
    .A2(_11085_),
    .ZN(_11086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19999_ (.A1(_11084_),
    .A2(_11086_),
    .A3(_10610_),
    .ZN(_11087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20000_ (.A1(_10566_),
    .A2(net1262),
    .ZN(_11088_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20001_ (.A1(_10866_),
    .A2(_11088_),
    .B(_10686_),
    .ZN(_11089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20002_ (.A1(_10716_),
    .A2(_10497_),
    .ZN(_11090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20003_ (.A1(_10865_),
    .A2(_10773_),
    .ZN(_11091_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20004_ (.A1(_11090_),
    .A2(_11091_),
    .A3(_10659_),
    .ZN(_11092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20005_ (.A1(_11089_),
    .A2(_11092_),
    .ZN(_11093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20006_ (.A1(_11087_),
    .A2(_11093_),
    .A3(_10632_),
    .ZN(_11094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20007_ (.A1(_11083_),
    .A2(_11094_),
    .A3(_10642_),
    .ZN(_11095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20008_ (.A1(_11070_),
    .A2(_11095_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20009_ (.A1(_10538_),
    .A2(_10499_),
    .Z(_11096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20010_ (.A1(_11096_),
    .A2(_10510_),
    .Z(_11097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20011_ (.A1(_10699_),
    .A2(_10540_),
    .ZN(_11098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20012_ (.A1(_11097_),
    .A2(_11098_),
    .B(_10557_),
    .ZN(_11099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20013_ (.A1(_10594_),
    .A2(_15680_),
    .ZN(_11100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20014_ (.A1(_11052_),
    .A2(_10668_),
    .A3(_11100_),
    .ZN(_11101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20015_ (.A1(_11099_),
    .A2(_11101_),
    .B(_10696_),
    .ZN(_11102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20016_ (.I(_10615_),
    .ZN(_11103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20017_ (.A1(net593),
    .A2(_10597_),
    .ZN(_11104_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20018_ (.A1(_11103_),
    .A2(_10952_),
    .B1(_11104_),
    .B2(_10594_),
    .ZN(_11105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20019_ (.A1(_11105_),
    .A2(_10853_),
    .ZN(_11106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20020_ (.A1(_11088_),
    .A2(_10572_),
    .Z(_11107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20021_ (.A1(_11103_),
    .A2(_10509_),
    .ZN(_11108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20022_ (.A1(_11107_),
    .A2(_11108_),
    .Z(_11109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20023_ (.A1(_11109_),
    .A2(_10915_),
    .B(_10610_),
    .ZN(_11110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20024_ (.A1(_11106_),
    .A2(_11110_),
    .ZN(_11111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20025_ (.A1(_11102_),
    .A2(_11111_),
    .ZN(_11112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20026_ (.A1(_10712_),
    .A2(_10704_),
    .ZN(_11113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20027_ (.A1(_10650_),
    .A2(_10646_),
    .ZN(_11114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20028_ (.A1(_11113_),
    .A2(_11114_),
    .A3(_10668_),
    .ZN(_11115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20029_ (.A1(_10649_),
    .A2(_10625_),
    .Z(_11116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20030_ (.A1(_10505_),
    .A2(_15701_),
    .ZN(_11117_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20031_ (.A1(_11116_),
    .A2(_10540_),
    .B(_10600_),
    .C(_11117_),
    .ZN(_11118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20032_ (.A1(_11115_),
    .A2(_11118_),
    .A3(_10661_),
    .ZN(_11119_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20033_ (.A1(_15687_),
    .A2(_10594_),
    .B(_10510_),
    .C(_10605_),
    .ZN(_11120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20034_ (.A1(_10730_),
    .A2(_10942_),
    .A3(_11107_),
    .ZN(_11121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20035_ (.A1(_11120_),
    .A2(_11121_),
    .A3(_10557_),
    .ZN(_11122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20036_ (.A1(_11119_),
    .A2(_11122_),
    .A3(_10591_),
    .ZN(_11123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20037_ (.A1(_11112_),
    .A2(_11123_),
    .A3(_10643_),
    .ZN(_11124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20038_ (.A1(_10448_),
    .A2(_10540_),
    .B(_10533_),
    .ZN(_11125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20039_ (.A1(_10648_),
    .A2(_10677_),
    .ZN(_11126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20040_ (.A1(_11125_),
    .A2(_11126_),
    .B(_10557_),
    .ZN(_11127_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20041_ (.A1(_10867_),
    .A2(_10771_),
    .Z(_11128_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20042_ (.A1(_10901_),
    .A2(_10674_),
    .A3(_11128_),
    .Z(_11129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20043_ (.A1(_11129_),
    .A2(_11127_),
    .B(_10632_),
    .ZN(_11130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20044_ (.A1(net80),
    .A2(_10540_),
    .B(_10980_),
    .ZN(_11131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20045_ (.A1(_11131_),
    .A2(_10668_),
    .ZN(_11132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20046_ (.A1(_10677_),
    .A2(_10594_),
    .A3(_10704_),
    .ZN(_11133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20047_ (.A1(_10835_),
    .A2(_11133_),
    .ZN(_11134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20048_ (.A1(_11132_),
    .A2(_11134_),
    .A3(_10579_),
    .ZN(_11135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20049_ (.A1(_11135_),
    .A2(_11130_),
    .ZN(_11136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20050_ (.A1(_10448_),
    .A2(_10712_),
    .ZN(_11137_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20051_ (.A1(_10892_),
    .A2(_11137_),
    .A3(_10847_),
    .ZN(_11138_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20052_ (.A1(_10716_),
    .A2(_10674_),
    .ZN(_11139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20053_ (.A1(_11139_),
    .A2(_10944_),
    .B(_10686_),
    .ZN(_11140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20054_ (.A1(_11138_),
    .A2(_11140_),
    .B(_10696_),
    .ZN(_11141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20055_ (.A1(_10843_),
    .A2(_10600_),
    .A3(_11043_),
    .ZN(_11142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20056_ (.A1(_10909_),
    .A2(_10758_),
    .A3(_10659_),
    .ZN(_11143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20057_ (.A1(_11142_),
    .A2(_11143_),
    .A3(_10610_),
    .ZN(_11144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20058_ (.A1(_11141_),
    .A2(_11144_),
    .B(_10643_),
    .ZN(_11145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20059_ (.A1(_11145_),
    .A2(_11136_),
    .ZN(_11146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20060_ (.A1(_11146_),
    .A2(_11124_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20061_ (.A1(\sa21_sr[1] ),
    .A2(\sa30_sub[1] ),
    .Z(_11147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20062_ (.I(\sa01_sr[7] ),
    .ZN(_11148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20063_ (.I(\sa01_sr[0] ),
    .ZN(_11149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20064_ (.A1(_11149_),
    .A2(_11148_),
    .ZN(_11150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20065_ (.A1(net1022),
    .A2(net799),
    .ZN(_11151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20066_ (.A1(_11151_),
    .A2(_11150_),
    .ZN(_11152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20067_ (.A1(_11152_),
    .A2(_11147_),
    .ZN(_11153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20068_ (.A1(_11149_),
    .A2(net1022),
    .ZN(_11154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20069_ (.A1(_11148_),
    .A2(\sa01_sr[0] ),
    .ZN(_11155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20070_ (.A1(_11155_),
    .A2(_11154_),
    .ZN(_11156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20071_ (.I(\sa21_sr[1] ),
    .ZN(_11157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20072_ (.I(\sa30_sub[1] ),
    .ZN(_11158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20073_ (.A1(_11157_),
    .A2(_11158_),
    .ZN(_11159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20074_ (.A1(net947),
    .A2(\sa30_sub[1] ),
    .ZN(_11160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20075_ (.A1(_11159_),
    .A2(_11160_),
    .ZN(_11161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20076_ (.A1(_11156_),
    .A2(_11161_),
    .ZN(_11162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20077_ (.A1(_11153_),
    .A2(_11162_),
    .ZN(_11163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20078_ (.I(_11163_),
    .ZN(_11164_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20079_ (.I(\sa11_sr[7] ),
    .ZN(_11165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20080_ (.I(\sa11_sr[0] ),
    .ZN(_11166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20081_ (.A1(_11166_),
    .A2(_11165_),
    .ZN(_11167_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20082_ (.I(\sa11_sr[7] ),
    .Z(_11168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20083_ (.A1(_11168_),
    .A2(\sa11_sr[0] ),
    .ZN(_11169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20084_ (.A1(_11169_),
    .A2(_11167_),
    .ZN(_11170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20085_ (.A1(_11170_),
    .A2(net805),
    .ZN(_11171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20086_ (.A1(_11166_),
    .A2(_11168_),
    .ZN(_11172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20087_ (.A1(_11165_),
    .A2(\sa11_sr[0] ),
    .ZN(_11173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20088_ (.A1(_11172_),
    .A2(_11173_),
    .ZN(_11174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20089_ (.I(\sa11_sr[1] ),
    .ZN(_11175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20090_ (.A1(_11174_),
    .A2(_11175_),
    .ZN(_11176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20091_ (.A1(_11171_),
    .A2(_11176_),
    .ZN(_11177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20092_ (.I(_11177_),
    .ZN(_11178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20093_ (.A1(_11164_),
    .A2(_11178_),
    .ZN(_11179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20094_ (.A1(_11163_),
    .A2(_11177_),
    .ZN(_11180_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20095_ (.A1(_11180_),
    .A2(_10522_),
    .A3(_11179_),
    .ZN(_11181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20096_ (.A1(_10525_),
    .A2(\text_in_r[89] ),
    .ZN(_11182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20097_ (.A1(_11182_),
    .A2(_11181_),
    .ZN(_11183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20098_ (.A1(_11183_),
    .A2(_07913_),
    .ZN(_11184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20099_ (.A1(_11181_),
    .A2(net654),
    .A3(_11182_),
    .ZN(_11185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20100_ (.A1(_11185_),
    .A2(_11184_),
    .ZN(_11186_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20101_ (.I(_11186_),
    .Z(_15711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20102_ (.A1(_11148_),
    .A2(_11165_),
    .ZN(_11187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20103_ (.A1(\sa01_sr[7] ),
    .A2(_11168_),
    .ZN(_11188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20104_ (.A1(_11187_),
    .A2(_11188_),
    .ZN(_11189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20105_ (.I(\sa30_sub[0] ),
    .ZN(_11190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20106_ (.A1(_11189_),
    .A2(_11190_),
    .ZN(_11191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20107_ (.A1(_11187_),
    .A2(net517),
    .A3(_11188_),
    .ZN(_11192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20108_ (.A1(_11166_),
    .A2(net814),
    .ZN(_11193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20109_ (.I(\sa21_sr[0] ),
    .ZN(_11194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20110_ (.A1(_11194_),
    .A2(net796),
    .ZN(_11195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20111_ (.A1(_11193_),
    .A2(_11195_),
    .ZN(_11196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20112_ (.A1(_11191_),
    .A2(_11192_),
    .A3(_11196_),
    .ZN(_11197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20113_ (.A1(_11189_),
    .A2(net517),
    .ZN(_11198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20114_ (.A1(_11187_),
    .A2(_11190_),
    .A3(_11188_),
    .ZN(_11199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20115_ (.I(_11196_),
    .ZN(_11200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20116_ (.A1(_11198_),
    .A2(_11199_),
    .A3(_11200_),
    .ZN(_11201_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _20117_ (.I(net475),
    .Z(_11202_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _20118_ (.I(_11202_),
    .Z(_11203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20119_ (.A1(_11197_),
    .A2(_11201_),
    .B(_11203_),
    .ZN(_11204_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20120_ (.I(\text_in_r[88] ),
    .ZN(_11205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20121_ (.A1(_11205_),
    .A2(_10431_),
    .Z(_11206_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20122_ (.A1(_11204_),
    .A2(_11206_),
    .B(net699),
    .ZN(_11207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20123_ (.A1(_11197_),
    .A2(_11201_),
    .ZN(_11208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20124_ (.A1(_11208_),
    .A2(_10489_),
    .ZN(_11209_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20125_ (.I(_11206_),
    .ZN(_11210_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20126_ (.A1(_11209_),
    .A2(_07908_),
    .A3(_11210_),
    .ZN(_11211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20127_ (.A1(_11207_),
    .A2(_11211_),
    .ZN(_15714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20128_ (.I(\sa01_sr[1] ),
    .ZN(_11212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20129_ (.A1(_11175_),
    .A2(_11212_),
    .ZN(_11213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20130_ (.A1(net807),
    .A2(\sa01_sr[1] ),
    .ZN(_11214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20131_ (.A1(_11213_),
    .A2(_11214_),
    .ZN(_11215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20132_ (.I(\sa21_sr[2] ),
    .ZN(_11216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20133_ (.A1(net1239),
    .A2(_11216_),
    .ZN(_11217_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20134_ (.I(\sa21_sr[2] ),
    .Z(_11218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20135_ (.A1(_11213_),
    .A2(_11218_),
    .A3(_11214_),
    .ZN(_11219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20136_ (.A1(_11217_),
    .A2(_11219_),
    .ZN(_11220_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20137_ (.I(\sa30_sub[2] ),
    .ZN(_11221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20138_ (.A1(_11221_),
    .A2(\sa11_sr[2] ),
    .ZN(_11222_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20139_ (.I(\sa11_sr[2] ),
    .ZN(_11223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20140_ (.A1(_11223_),
    .A2(\sa30_sub[2] ),
    .ZN(_11224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20141_ (.A1(_11222_),
    .A2(_11224_),
    .ZN(_11225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20142_ (.I(_11225_),
    .ZN(_11226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20143_ (.A1(_11220_),
    .A2(_11226_),
    .ZN(_11227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20144_ (.A1(_11217_),
    .A2(_11219_),
    .A3(_11225_),
    .ZN(_11228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20145_ (.A1(_11227_),
    .A2(_11228_),
    .B(_10482_),
    .ZN(_11229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20146_ (.I(\text_in_r[90] ),
    .ZN(_11230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20147_ (.A1(_11230_),
    .A2(_11202_),
    .Z(_11231_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20148_ (.A1(_11229_),
    .A2(_11231_),
    .B(_07917_),
    .ZN(_11232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20149_ (.A1(_11227_),
    .A2(_11228_),
    .ZN(_11233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20150_ (.A1(_11233_),
    .A2(_10402_),
    .ZN(_11234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20151_ (.I(_11231_),
    .ZN(_11235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20152_ (.A1(_11234_),
    .A2(net767),
    .A3(_11235_),
    .ZN(_11236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20153_ (.A1(_11232_),
    .A2(_11236_),
    .ZN(_11237_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20154_ (.I(_11237_),
    .Z(_11238_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20155_ (.I(_11238_),
    .Z(_15730_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20156_ (.A1(_11204_),
    .A2(_11206_),
    .B(_07908_),
    .ZN(_11239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20157_ (.A1(_11209_),
    .A2(net698),
    .A3(_11210_),
    .ZN(_11240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20158_ (.A1(_11240_),
    .A2(_11239_),
    .ZN(_15705_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20159_ (.A1(_11229_),
    .A2(_11231_),
    .B(net767),
    .ZN(_11241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20160_ (.A1(_11234_),
    .A2(_07917_),
    .A3(_11235_),
    .ZN(_11242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20161_ (.A1(_11241_),
    .A2(_11242_),
    .ZN(_11243_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20162_ (.I(_11243_),
    .Z(_15723_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20163_ (.I(_15715_),
    .ZN(_11244_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20164_ (.A1(_11238_),
    .A2(_11244_),
    .Z(_11245_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20165_ (.I(_15707_),
    .ZN(_11246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20166_ (.A1(_11232_),
    .A2(_11236_),
    .A3(_11246_),
    .ZN(_11247_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20167_ (.I(_11247_),
    .ZN(_11248_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20168_ (.A1(\sa21_sr[3] ),
    .A2(\sa30_sub[3] ),
    .Z(_11249_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20169_ (.I(\sa01_sr[2] ),
    .ZN(_11250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20170_ (.A1(_11148_),
    .A2(_11250_),
    .ZN(_11251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20171_ (.A1(net1022),
    .A2(\sa01_sr[2] ),
    .ZN(_11252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20172_ (.A1(_11251_),
    .A2(_11252_),
    .ZN(_11253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20173_ (.A1(_11249_),
    .A2(_11253_),
    .ZN(_11254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20174_ (.A1(_11250_),
    .A2(net35),
    .ZN(_11255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20175_ (.A1(_11148_),
    .A2(\sa01_sr[2] ),
    .ZN(_11256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20176_ (.A1(_11255_),
    .A2(_11256_),
    .ZN(_11257_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20177_ (.I(\sa21_sr[3] ),
    .ZN(_11258_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20178_ (.I(\sa30_sub[3] ),
    .ZN(_11259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20179_ (.A1(_11258_),
    .A2(_11259_),
    .ZN(_11260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20180_ (.A1(\sa21_sr[3] ),
    .A2(\sa30_sub[3] ),
    .ZN(_11261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20181_ (.A1(_11260_),
    .A2(_11261_),
    .ZN(_11262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20182_ (.A1(_11257_),
    .A2(_11262_),
    .ZN(_11263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20183_ (.A1(_11254_),
    .A2(_11263_),
    .ZN(_11264_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20184_ (.I(_11264_),
    .ZN(_11265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20185_ (.I(\sa11_sr[3] ),
    .ZN(_11266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20186_ (.A1(_11266_),
    .A2(net523),
    .ZN(_11267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20187_ (.A1(_11165_),
    .A2(\sa11_sr[3] ),
    .ZN(_11268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20188_ (.A1(_11267_),
    .A2(_11268_),
    .ZN(_11269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20189_ (.A1(_11269_),
    .A2(\sa11_sr[2] ),
    .ZN(_11270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20190_ (.A1(_11165_),
    .A2(_11266_),
    .ZN(_11271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20191_ (.A1(\sa11_sr[7] ),
    .A2(\sa11_sr[3] ),
    .ZN(_11272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20192_ (.A1(_11271_),
    .A2(_11272_),
    .ZN(_11273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20193_ (.A1(_11273_),
    .A2(_11223_),
    .ZN(_11274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20194_ (.A1(_11270_),
    .A2(_11274_),
    .ZN(_11275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20195_ (.A1(_11265_),
    .A2(_11275_),
    .ZN(_11276_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20196_ (.I(_11275_),
    .ZN(_11277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20197_ (.A1(_11277_),
    .A2(_11264_),
    .ZN(_11278_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20198_ (.I(_10402_),
    .Z(_11279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20199_ (.A1(_11276_),
    .A2(_11278_),
    .A3(_11279_),
    .ZN(_11280_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20200_ (.A1(_10411_),
    .A2(\text_in_r[91] ),
    .ZN(_11281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20201_ (.A1(_11280_),
    .A2(_07921_),
    .A3(_11281_),
    .ZN(_11282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20202_ (.A1(_11265_),
    .A2(_11277_),
    .ZN(_11283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20203_ (.A1(_11264_),
    .A2(_11275_),
    .ZN(_11284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20204_ (.A1(_11283_),
    .A2(_11279_),
    .A3(_11284_),
    .ZN(_11285_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20205_ (.A1(_10489_),
    .A2(\text_in_r[91] ),
    .Z(_11286_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20206_ (.A1(_11285_),
    .A2(\u0.w[1][27] ),
    .A3(_11286_),
    .ZN(_11287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20207_ (.A1(_11282_),
    .A2(_11287_),
    .ZN(_11288_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20208_ (.I(_11288_),
    .Z(_11289_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20209_ (.I(_11289_),
    .Z(_11290_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20210_ (.A1(_11245_),
    .A2(_11248_),
    .B(_11290_),
    .ZN(_11291_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20211_ (.I(_15708_),
    .ZN(_11292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20212_ (.A1(_11232_),
    .A2(_11236_),
    .A3(_11292_),
    .ZN(_11293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20213_ (.A1(_11280_),
    .A2(\u0.w[1][27] ),
    .A3(_11281_),
    .ZN(_11294_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20214_ (.A1(_11285_),
    .A2(_07921_),
    .A3(_11286_),
    .ZN(_11295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20215_ (.A1(_11294_),
    .A2(_11295_),
    .ZN(_11296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20216_ (.A1(_11293_),
    .A2(_11296_),
    .ZN(_11297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20217_ (.I(_11297_),
    .ZN(_11298_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20218_ (.A1(_11241_),
    .A2(_11242_),
    .A3(_15707_),
    .ZN(_11299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20219_ (.A1(_11298_),
    .A2(_11299_),
    .ZN(_11300_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20220_ (.A1(net35),
    .A2(\sa01_sr[3] ),
    .Z(_11301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20221_ (.A1(\sa21_sr[4] ),
    .A2(\sa30_sub[4] ),
    .Z(_11302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20222_ (.A1(\sa21_sr[4] ),
    .A2(\sa30_sub[4] ),
    .ZN(_11303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20223_ (.A1(_11302_),
    .A2(_11303_),
    .ZN(_11304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20224_ (.I(_11304_),
    .ZN(_11305_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20225_ (.A1(_11301_),
    .A2(_11305_),
    .Z(_11306_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20226_ (.A1(\sa11_sr[4] ),
    .A2(_11273_),
    .Z(_11307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20227_ (.I(_11307_),
    .ZN(_11308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20228_ (.A1(_11306_),
    .A2(_11308_),
    .ZN(_11309_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20229_ (.A1(_11304_),
    .A2(_11301_),
    .Z(_11310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20230_ (.A1(_11310_),
    .A2(_11307_),
    .ZN(_11311_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20231_ (.A1(_11309_),
    .A2(_11311_),
    .A3(_10523_),
    .ZN(_11312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20232_ (.A1(_10526_),
    .A2(\text_in_r[92] ),
    .ZN(_11313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20233_ (.A1(_11312_),
    .A2(_11313_),
    .ZN(_11314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20234_ (.A1(_11314_),
    .A2(\u0.w[1][28] ),
    .ZN(_11315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20235_ (.A1(_11312_),
    .A2(_07925_),
    .A3(_11313_),
    .ZN(_11316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20236_ (.A1(_11315_),
    .A2(_11316_),
    .ZN(_11317_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20237_ (.I(_11317_),
    .Z(_11318_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20238_ (.I(_11318_),
    .Z(_11319_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20239_ (.A1(_11291_),
    .A2(_11300_),
    .A3(_11319_),
    .ZN(_11320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20240_ (.A1(net654),
    .A2(_11183_),
    .ZN(_11321_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20241_ (.A1(_11181_),
    .A2(_07913_),
    .A3(_11182_),
    .ZN(_11322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20242_ (.A1(_11322_),
    .A2(_11321_),
    .ZN(_15706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20243_ (.A1(net1),
    .A2(_11289_),
    .A3(_15730_),
    .ZN(_11323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20244_ (.I(_11293_),
    .ZN(_11324_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20245_ (.I(_11288_),
    .Z(_11325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20246_ (.A1(_11325_),
    .A2(_11324_),
    .ZN(_11326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20247_ (.A1(_11238_),
    .A2(_11292_),
    .ZN(_11327_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20248_ (.I(_11296_),
    .Z(_11328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20249_ (.A1(_11327_),
    .A2(_11328_),
    .ZN(_11329_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20250_ (.A1(_11323_),
    .A2(_11326_),
    .A3(_11329_),
    .ZN(_11330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20251_ (.A1(_11314_),
    .A2(_07925_),
    .ZN(_11331_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20252_ (.A1(_11312_),
    .A2(\u0.w[1][28] ),
    .A3(_11313_),
    .ZN(_11332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20253_ (.A1(_11331_),
    .A2(_11332_),
    .ZN(_11333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20254_ (.I(_11333_),
    .Z(_11334_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20255_ (.I(_11334_),
    .Z(_11335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20256_ (.A1(_11330_),
    .A2(_11335_),
    .ZN(_11336_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20257_ (.A1(\sa21_sr[5] ),
    .A2(\sa30_sub[5] ),
    .Z(_11337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20258_ (.A1(\sa21_sr[5] ),
    .A2(\sa30_sub[5] ),
    .ZN(_11338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20259_ (.A1(_11337_),
    .A2(_11338_),
    .ZN(_11339_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20260_ (.A1(\sa11_sr[5] ),
    .A2(_11339_),
    .Z(_11340_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20261_ (.A1(\sa11_sr[4] ),
    .A2(\sa01_sr[4] ),
    .Z(_11341_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20262_ (.I(_11341_),
    .ZN(_11342_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20263_ (.A1(_11340_),
    .A2(_11342_),
    .Z(_11343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20264_ (.A1(_11340_),
    .A2(_11342_),
    .ZN(_11344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20265_ (.A1(_11343_),
    .A2(_11344_),
    .ZN(_11345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20266_ (.A1(_10587_),
    .A2(\text_in_r[93] ),
    .ZN(_11346_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20267_ (.A1(_11345_),
    .A2(_10639_),
    .B(_07929_),
    .C(_11346_),
    .ZN(_11347_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _20268_ (.I(_10489_),
    .Z(_11348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20269_ (.A1(_11343_),
    .A2(_11348_),
    .A3(_11344_),
    .ZN(_11349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20270_ (.A1(_11349_),
    .A2(_11346_),
    .ZN(_11350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20271_ (.A1(_11350_),
    .A2(\u0.w[1][29] ),
    .ZN(_11351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20272_ (.A1(_11347_),
    .A2(_11351_),
    .ZN(_11352_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20273_ (.I(_11352_),
    .Z(_11353_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20274_ (.I(_11353_),
    .Z(_11354_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20275_ (.A1(_11320_),
    .A2(_11336_),
    .A3(_11354_),
    .ZN(_11355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20276_ (.A1(_11243_),
    .A2(_15714_),
    .ZN(_11356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20277_ (.A1(_11356_),
    .A2(_11288_),
    .ZN(_11357_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20278_ (.I(_11357_),
    .ZN(_11358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20279_ (.A1(net1),
    .A2(net843),
    .ZN(_11359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20280_ (.A1(_11358_),
    .A2(_11359_),
    .ZN(_11360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20281_ (.A1(_15711_),
    .A2(net844),
    .ZN(_11361_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20282_ (.I(_11296_),
    .Z(_11362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20283_ (.A1(_11238_),
    .A2(_15714_),
    .ZN(_11363_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20284_ (.A1(_11361_),
    .A2(_11362_),
    .A3(_11363_),
    .ZN(_11364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20285_ (.A1(_11360_),
    .A2(_11364_),
    .A3(_11335_),
    .ZN(_11365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20286_ (.A1(_15711_),
    .A2(_15714_),
    .A3(_11238_),
    .ZN(_11366_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20287_ (.A1(_11293_),
    .A2(_11325_),
    .Z(_11367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20288_ (.A1(_11366_),
    .A2(_11367_),
    .ZN(_11368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20289_ (.A1(_15730_),
    .A2(_11246_),
    .ZN(_11369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20290_ (.A1(_15723_),
    .A2(_11244_),
    .ZN(_11370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20291_ (.A1(_11369_),
    .A2(_11370_),
    .ZN(_11371_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20292_ (.I(_11328_),
    .Z(_11372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20293_ (.A1(_11371_),
    .A2(_11372_),
    .ZN(_11373_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20294_ (.I(_11318_),
    .Z(_11374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20295_ (.A1(_11368_),
    .A2(_11373_),
    .A3(_11374_),
    .ZN(_11375_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20296_ (.I(_11352_),
    .ZN(_11376_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20297_ (.I(_11376_),
    .Z(_11377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20298_ (.A1(_11365_),
    .A2(_11375_),
    .A3(_11377_),
    .ZN(_11378_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20299_ (.A1(\sa11_sr[5] ),
    .A2(\sa01_sr[5] ),
    .ZN(_11379_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20300_ (.A1(\sa21_sr[6] ),
    .A2(\sa30_sub[6] ),
    .Z(_11380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20301_ (.A1(\sa21_sr[6] ),
    .A2(\sa30_sub[6] ),
    .ZN(_11381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20302_ (.A1(_11380_),
    .A2(_11381_),
    .ZN(_11382_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20303_ (.A1(\sa11_sr[6] ),
    .A2(_11382_),
    .Z(_11383_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20304_ (.A1(_11379_),
    .A2(_11383_),
    .Z(_11384_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20305_ (.I(_10525_),
    .Z(_11385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20306_ (.A1(_11385_),
    .A2(\text_in_r[94] ),
    .Z(_11386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20307_ (.A1(_11384_),
    .A2(_10585_),
    .B(_11386_),
    .ZN(_11387_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _20308_ (.A1(_07729_),
    .A2(_11387_),
    .Z(_11388_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20309_ (.I(_11388_),
    .ZN(_11389_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20310_ (.I(_11389_),
    .Z(_11390_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20311_ (.A1(_11355_),
    .A2(_11378_),
    .A3(_11390_),
    .ZN(_11391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20312_ (.A1(_11237_),
    .A2(_15705_),
    .ZN(_11392_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20313_ (.I(_11392_),
    .ZN(_11393_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20314_ (.I(_15721_),
    .ZN(_11394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20315_ (.A1(_15723_),
    .A2(_11394_),
    .ZN(_11395_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20316_ (.I(_11395_),
    .ZN(_11396_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20317_ (.I(_11288_),
    .Z(_11397_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20318_ (.A1(_11393_),
    .A2(_11396_),
    .A3(_11397_),
    .Z(_11398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20319_ (.A1(net42),
    .A2(_11393_),
    .ZN(_11399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20320_ (.A1(net1023),
    .A2(_11243_),
    .ZN(_11400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20321_ (.A1(_11399_),
    .A2(_11290_),
    .A3(_11400_),
    .ZN(_11401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20322_ (.A1(_11398_),
    .A2(_11401_),
    .A3(_11335_),
    .ZN(_11402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20323_ (.A1(_11232_),
    .A2(_11236_),
    .A3(_15709_),
    .ZN(_11403_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20324_ (.I(_11296_),
    .Z(_11404_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20325_ (.A1(_11403_),
    .A2(_11404_),
    .ZN(_11405_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20326_ (.I(_11405_),
    .ZN(_11406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20327_ (.A1(_11406_),
    .A2(_11323_),
    .Z(_11407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20328_ (.A1(_11404_),
    .A2(_15723_),
    .ZN(_11408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20329_ (.A1(_11404_),
    .A2(_15714_),
    .ZN(_11409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20330_ (.A1(_11408_),
    .A2(_11409_),
    .ZN(_11410_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20331_ (.I(_11356_),
    .ZN(_11411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20332_ (.A1(_11411_),
    .A2(net42),
    .ZN(_11412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20333_ (.A1(_11410_),
    .A2(_11412_),
    .ZN(_11413_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20334_ (.A1(_11407_),
    .A2(_11413_),
    .A3(_11319_),
    .ZN(_11414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20335_ (.A1(_11402_),
    .A2(_11354_),
    .A3(_11414_),
    .ZN(_11415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20336_ (.A1(_11392_),
    .A2(_11288_),
    .ZN(_11416_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20337_ (.I(_11317_),
    .Z(_11417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20338_ (.A1(_11416_),
    .A2(_11417_),
    .Z(_11418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20339_ (.A1(_11241_),
    .A2(_11242_),
    .B(_15712_),
    .ZN(_11419_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20340_ (.A1(_11419_),
    .A2(_11325_),
    .ZN(_11420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20341_ (.A1(_11399_),
    .A2(_11420_),
    .ZN(_11421_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20342_ (.I(_11352_),
    .Z(_11422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20343_ (.A1(_11418_),
    .A2(_11421_),
    .B(_11422_),
    .ZN(_11423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20344_ (.A1(_11243_),
    .A2(net841),
    .ZN(_11424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20345_ (.A1(_15730_),
    .A2(_15721_),
    .ZN(_11425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20346_ (.A1(_11424_),
    .A2(_11425_),
    .ZN(_11426_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20347_ (.I(_11318_),
    .Z(_11427_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20348_ (.A1(_11426_),
    .A2(_11372_),
    .B(_11427_),
    .ZN(_11428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20349_ (.A1(_11243_),
    .A2(net843),
    .ZN(_11429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20350_ (.A1(_11429_),
    .A2(_11325_),
    .Z(_11430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20351_ (.A1(_11430_),
    .A2(_11361_),
    .ZN(_11431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20352_ (.A1(_11428_),
    .A2(_11431_),
    .ZN(_11432_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20353_ (.I(_11389_),
    .Z(_11433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20354_ (.A1(_11423_),
    .A2(_11432_),
    .B(_11433_),
    .ZN(_11434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20355_ (.A1(_11415_),
    .A2(_11434_),
    .ZN(_11435_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _20356_ (.I(\sa21_sr[7] ),
    .Z(_11436_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20357_ (.A1(\sa11_sr[6] ),
    .A2(\sa01_sr[6] ),
    .Z(_11437_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20358_ (.A1(net524),
    .A2(_11437_),
    .Z(_11438_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _20359_ (.A1(net26),
    .A2(net819),
    .A3(_11438_),
    .Z(_11439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20360_ (.I0(_11439_),
    .I1(\text_in_r[95] ),
    .S(_10639_),
    .Z(_11440_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20361_ (.A1(_07936_),
    .A2(_11440_),
    .Z(_11441_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20362_ (.I(_11441_),
    .Z(_11442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20363_ (.A1(_11391_),
    .A2(_11435_),
    .A3(_11442_),
    .ZN(_11443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20364_ (.A1(_11241_),
    .A2(_11242_),
    .A3(_15708_),
    .ZN(_11444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20365_ (.A1(_11328_),
    .A2(_11444_),
    .B(_11333_),
    .ZN(_11445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20366_ (.A1(_11404_),
    .A2(_15728_),
    .Z(_11446_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20367_ (.A1(_11445_),
    .A2(_11446_),
    .Z(_11447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20368_ (.A1(_11447_),
    .A2(_11353_),
    .Z(_11448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20369_ (.A1(_11363_),
    .A2(_11247_),
    .ZN(_11449_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20370_ (.I(_11404_),
    .Z(_11450_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20371_ (.I(_11333_),
    .Z(_11451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20372_ (.A1(_11449_),
    .A2(_11450_),
    .B(_11451_),
    .ZN(_11452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20373_ (.A1(_11243_),
    .A2(net980),
    .ZN(_11453_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20374_ (.I(_15712_),
    .ZN(_11454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20375_ (.A1(_15730_),
    .A2(_11454_),
    .ZN(_11455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20376_ (.A1(_11453_),
    .A2(_11289_),
    .A3(_11455_),
    .ZN(_11456_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20377_ (.I(_15709_),
    .ZN(_11457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20378_ (.A1(_15730_),
    .A2(_11457_),
    .ZN(_11458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20379_ (.A1(_11430_),
    .A2(_11458_),
    .ZN(_11459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20380_ (.A1(_11452_),
    .A2(_11456_),
    .A3(_11459_),
    .ZN(_11460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20381_ (.A1(_11448_),
    .A2(_11460_),
    .ZN(_11461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20382_ (.I(_11403_),
    .ZN(_11462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20383_ (.A1(_11462_),
    .A2(_11328_),
    .ZN(_11463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20384_ (.A1(_11463_),
    .A2(_11334_),
    .Z(_11464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20385_ (.I(_11429_),
    .ZN(_11465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20386_ (.A1(_11465_),
    .A2(net42),
    .ZN(_11466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20387_ (.A1(_11238_),
    .A2(_15715_),
    .ZN(_11467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20388_ (.A1(_11467_),
    .A2(_11288_),
    .ZN(_11468_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20389_ (.I(_11468_),
    .ZN(_11469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20390_ (.A1(_11466_),
    .A2(_11469_),
    .ZN(_11470_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20391_ (.A1(_11464_),
    .A2(_11470_),
    .B(_11422_),
    .ZN(_11471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20392_ (.I(_15717_),
    .ZN(_11472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20393_ (.A1(_11238_),
    .A2(_11472_),
    .ZN(_11473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20394_ (.A1(_11473_),
    .A2(_11296_),
    .ZN(_11474_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20395_ (.I(_11474_),
    .ZN(_11475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20396_ (.A1(_11466_),
    .A2(_11475_),
    .ZN(_11476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20397_ (.A1(_11476_),
    .A2(_11319_),
    .A3(_11406_),
    .ZN(_11477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20398_ (.A1(_11471_),
    .A2(_11477_),
    .ZN(_11478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20399_ (.A1(_11461_),
    .A2(_11478_),
    .A3(_11390_),
    .ZN(_11479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20400_ (.A1(_11453_),
    .A2(_11288_),
    .Z(_11480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20401_ (.A1(_11480_),
    .A2(_11444_),
    .ZN(_11481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20402_ (.A1(_11467_),
    .A2(_11328_),
    .Z(_11482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20403_ (.A1(_11482_),
    .A2(_11429_),
    .ZN(_11483_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20404_ (.A1(_11481_),
    .A2(_11319_),
    .A3(_11483_),
    .ZN(_11484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20405_ (.I(_11369_),
    .ZN(_11485_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20406_ (.A1(_11485_),
    .A2(_11462_),
    .B(_11397_),
    .ZN(_11486_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20407_ (.A1(_11420_),
    .A2(_11427_),
    .ZN(_11487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20408_ (.A1(_11486_),
    .A2(_11487_),
    .B(_11353_),
    .ZN(_11488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20409_ (.A1(_11484_),
    .A2(_11488_),
    .B(_11433_),
    .ZN(_11489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20410_ (.A1(_11238_),
    .A2(_15712_),
    .ZN(_11490_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20411_ (.A1(_11490_),
    .A2(_11404_),
    .Z(_11491_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20412_ (.A1(_11491_),
    .A2(_11334_),
    .Z(_11492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20413_ (.A1(_11243_),
    .A2(_15717_),
    .ZN(_11493_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20414_ (.A1(_11493_),
    .A2(_11404_),
    .ZN(_11494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20415_ (.I(_11494_),
    .ZN(_11495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20416_ (.A1(_11492_),
    .A2(_11297_),
    .A3(_11495_),
    .ZN(_11496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20417_ (.A1(_11413_),
    .A2(_11491_),
    .A3(_11374_),
    .ZN(_11497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20418_ (.A1(_11496_),
    .A2(_11354_),
    .A3(_11497_),
    .ZN(_11498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20419_ (.A1(_11489_),
    .A2(_11498_),
    .ZN(_11499_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _20420_ (.I(_11442_),
    .ZN(_11500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20421_ (.A1(_11479_),
    .A2(_11499_),
    .A3(_11500_),
    .ZN(_11501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20422_ (.A1(_11443_),
    .A2(_11501_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20423_ (.A1(_11241_),
    .A2(_11394_),
    .A3(_11242_),
    .ZN(_11502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20424_ (.A1(_11502_),
    .A2(_11296_),
    .Z(_11503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20425_ (.A1(_11503_),
    .A2(_11400_),
    .B(_11318_),
    .ZN(_11504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20426_ (.A1(_11400_),
    .A2(_11429_),
    .ZN(_11505_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20427_ (.I(_11288_),
    .Z(_11506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20428_ (.A1(_11505_),
    .A2(_11506_),
    .ZN(_11507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20429_ (.A1(_11504_),
    .A2(_11507_),
    .ZN(_11508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20430_ (.A1(_11366_),
    .A2(_11362_),
    .A3(_11424_),
    .ZN(_11509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20431_ (.A1(_15723_),
    .A2(net979),
    .Z(_11510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20432_ (.A1(_11510_),
    .A2(_11506_),
    .B(_11334_),
    .ZN(_11511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20433_ (.A1(_11509_),
    .A2(_11511_),
    .ZN(_11512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20434_ (.A1(_11508_),
    .A2(_11512_),
    .ZN(_11513_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20435_ (.I(_11376_),
    .Z(_11514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20436_ (.A1(_11513_),
    .A2(_11514_),
    .ZN(_11515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20437_ (.A1(_11444_),
    .A2(_11325_),
    .ZN(_11516_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20438_ (.A1(_11516_),
    .A2(_11465_),
    .B(_11417_),
    .ZN(_11517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20439_ (.A1(_15711_),
    .A2(_15714_),
    .ZN(_11518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20440_ (.A1(_11518_),
    .A2(_11429_),
    .B(_11397_),
    .ZN(_11519_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20441_ (.A1(_11517_),
    .A2(_11519_),
    .ZN(_11520_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20442_ (.A1(_11363_),
    .A2(_11247_),
    .A3(_11397_),
    .ZN(_11521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20443_ (.A1(_11490_),
    .A2(_11293_),
    .A3(_11450_),
    .ZN(_11522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20444_ (.A1(_11521_),
    .A2(_11522_),
    .B(_11427_),
    .ZN(_11523_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20445_ (.I(_11352_),
    .Z(_11524_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20446_ (.A1(_11520_),
    .A2(_11523_),
    .B(_11524_),
    .ZN(_11525_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20447_ (.I(_11388_),
    .Z(_11526_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20448_ (.A1(_11515_),
    .A2(_11525_),
    .A3(_11526_),
    .ZN(_11527_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20449_ (.A1(_11296_),
    .A2(_15730_),
    .Z(_11528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20450_ (.A1(_11528_),
    .A2(_11361_),
    .B(_11334_),
    .ZN(_11529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20451_ (.A1(_11453_),
    .A2(_11359_),
    .A3(_11506_),
    .ZN(_11530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20452_ (.A1(_11529_),
    .A2(_11530_),
    .ZN(_11531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20453_ (.A1(_11243_),
    .A2(_11454_),
    .ZN(_11532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20454_ (.A1(_11363_),
    .A2(_11532_),
    .A3(_11506_),
    .ZN(_11533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20455_ (.A1(_11392_),
    .A2(_11293_),
    .A3(_11362_),
    .ZN(_11534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20456_ (.A1(_11533_),
    .A2(_11534_),
    .A3(_11451_),
    .ZN(_11535_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20457_ (.A1(_11531_),
    .A2(_11535_),
    .A3(_11376_),
    .ZN(_11536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20458_ (.A1(net42),
    .A2(_15730_),
    .ZN(_11537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20459_ (.A1(_11537_),
    .A2(_11362_),
    .B(_11318_),
    .ZN(_11538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20460_ (.A1(_11538_),
    .A2(_11456_),
    .B(_11376_),
    .ZN(_11539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20461_ (.A1(_11356_),
    .A2(_11490_),
    .ZN(_11540_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20462_ (.I(_11400_),
    .ZN(_11541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20463_ (.A1(_11540_),
    .A2(_11541_),
    .B(_11506_),
    .ZN(_11542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20464_ (.A1(_11243_),
    .A2(_15721_),
    .ZN(_11543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20465_ (.A1(_11543_),
    .A2(_11444_),
    .ZN(_11544_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20466_ (.A1(_11544_),
    .A2(_11362_),
    .B(_11333_),
    .ZN(_11545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20467_ (.A1(_11542_),
    .A2(_11545_),
    .ZN(_11546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20468_ (.A1(_11539_),
    .A2(_11546_),
    .ZN(_11547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20469_ (.A1(_11536_),
    .A2(_11547_),
    .ZN(_11548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20470_ (.A1(_11548_),
    .A2(_11390_),
    .ZN(_11549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20471_ (.A1(_11527_),
    .A2(_11549_),
    .ZN(_11550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20472_ (.A1(_11550_),
    .A2(_11500_),
    .ZN(_11551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20473_ (.I(_11363_),
    .ZN(_11552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20474_ (.A1(_11552_),
    .A2(_11397_),
    .B(_11417_),
    .ZN(_11553_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20475_ (.A1(_11247_),
    .A2(_11325_),
    .ZN(_11554_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20476_ (.A1(_11405_),
    .A2(_11554_),
    .ZN(_11555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20477_ (.I(_11444_),
    .ZN(_11556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20478_ (.A1(_11556_),
    .A2(_11328_),
    .ZN(_11557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20479_ (.A1(_11553_),
    .A2(_11555_),
    .A3(_11557_),
    .ZN(_11558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20480_ (.A1(net1),
    .A2(_11238_),
    .ZN(_11559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20481_ (.A1(_11420_),
    .A2(_11559_),
    .ZN(_11560_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20482_ (.A1(_11356_),
    .A2(_11299_),
    .A3(_11397_),
    .ZN(_11561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20483_ (.A1(_11560_),
    .A2(_11374_),
    .A3(_11561_),
    .ZN(_11562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20484_ (.A1(_11558_),
    .A2(_11562_),
    .A3(_11514_),
    .ZN(_11563_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20485_ (.I(_11416_),
    .ZN(_11564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20486_ (.A1(_11564_),
    .A2(_11412_),
    .ZN(_11565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20487_ (.A1(_11318_),
    .A2(_11297_),
    .Z(_11566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20488_ (.A1(_11565_),
    .A2(_11566_),
    .B(_11376_),
    .ZN(_11567_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20489_ (.A1(_11395_),
    .A2(_11289_),
    .Z(_11568_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20490_ (.A1(_11568_),
    .A2(_11458_),
    .B(_11427_),
    .ZN(_11569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20491_ (.A1(_11569_),
    .A2(_11509_),
    .ZN(_11570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20492_ (.A1(_11567_),
    .A2(_11570_),
    .ZN(_11571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20493_ (.A1(_11571_),
    .A2(_11563_),
    .B(_11390_),
    .ZN(_11572_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20494_ (.A1(_11429_),
    .A2(_11363_),
    .A3(net42),
    .ZN(_11573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20495_ (.A1(_11573_),
    .A2(_11372_),
    .ZN(_11574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20496_ (.A1(_11430_),
    .A2(_11299_),
    .ZN(_11575_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20497_ (.A1(_11574_),
    .A2(_11514_),
    .A3(_11575_),
    .ZN(_11576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20498_ (.A1(_11358_),
    .A2(_11537_),
    .ZN(_11577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20499_ (.A1(_11577_),
    .A2(_11422_),
    .A3(_11560_),
    .ZN(_11578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20500_ (.A1(_11576_),
    .A2(_11578_),
    .ZN(_11579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20501_ (.I(_15731_),
    .ZN(_11580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20502_ (.A1(_11362_),
    .A2(_11580_),
    .Z(_11581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20503_ (.A1(_11581_),
    .A2(_11353_),
    .B(_11451_),
    .ZN(_11582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20504_ (.A1(_11469_),
    .A2(_11412_),
    .ZN(_11583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20505_ (.A1(_11582_),
    .A2(_11583_),
    .ZN(_11584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20506_ (.A1(_11584_),
    .A2(_11433_),
    .ZN(_11585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20507_ (.A1(_11579_),
    .A2(_11335_),
    .B(_11585_),
    .ZN(_11586_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20508_ (.A1(_11572_),
    .A2(_11586_),
    .B(_11442_),
    .ZN(_11587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20509_ (.A1(_11551_),
    .A2(_11587_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20510_ (.A1(_11559_),
    .A2(_11404_),
    .Z(_11588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20511_ (.A1(_11588_),
    .A2(_11429_),
    .ZN(_11589_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20512_ (.A1(_11481_),
    .A2(_11589_),
    .B(_11524_),
    .ZN(_11590_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20513_ (.A1(_11444_),
    .A2(_11328_),
    .Z(_11591_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20514_ (.A1(_11591_),
    .A2(_11370_),
    .B(_11376_),
    .ZN(_11592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20515_ (.A1(_11480_),
    .A2(_11369_),
    .ZN(_11593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20516_ (.A1(_11592_),
    .A2(_11593_),
    .Z(_11594_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20517_ (.A1(_11590_),
    .A2(_11594_),
    .B(_11335_),
    .ZN(_11595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20518_ (.I(_11329_),
    .ZN(_11596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20519_ (.A1(_11466_),
    .A2(_11596_),
    .ZN(_11597_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20520_ (.I(_11289_),
    .Z(_11598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20521_ (.A1(_15728_),
    .A2(_11598_),
    .B(_11353_),
    .ZN(_11599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20522_ (.I(_11333_),
    .Z(_11600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20523_ (.A1(_11597_),
    .A2(_11599_),
    .B(_11600_),
    .ZN(_11601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20524_ (.A1(_11453_),
    .A2(_11359_),
    .A3(_11450_),
    .ZN(_11602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20525_ (.A1(_11290_),
    .A2(_11580_),
    .ZN(_11603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20526_ (.A1(_11602_),
    .A2(_11524_),
    .A3(_11603_),
    .ZN(_11604_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20527_ (.A1(_11601_),
    .A2(_11604_),
    .B(_11433_),
    .ZN(_11605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20528_ (.A1(_11595_),
    .A2(_11605_),
    .ZN(_11606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20529_ (.A1(_11457_),
    .A2(_11454_),
    .Z(_11607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20530_ (.I(_11607_),
    .ZN(_11608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20531_ (.A1(_15723_),
    .A2(_11608_),
    .ZN(_11609_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20532_ (.A1(_11559_),
    .A2(_11392_),
    .A3(_11609_),
    .ZN(_11610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20533_ (.A1(_11610_),
    .A2(_11372_),
    .ZN(_11611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20534_ (.A1(_11611_),
    .A2(_11335_),
    .A3(_11583_),
    .ZN(_11612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20535_ (.A1(_11248_),
    .A2(_11289_),
    .ZN(_11613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20536_ (.A1(_11613_),
    .A2(_11417_),
    .Z(_11614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20537_ (.A1(_11298_),
    .A2(_11455_),
    .ZN(_11615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20538_ (.A1(_11614_),
    .A2(_11615_),
    .B(_11422_),
    .ZN(_11616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20539_ (.A1(_11612_),
    .A2(_11616_),
    .ZN(_11617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20540_ (.A1(_11453_),
    .A2(_11361_),
    .A3(_11362_),
    .ZN(_11618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20541_ (.A1(_15735_),
    .A2(_11598_),
    .B(_11427_),
    .ZN(_11619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20542_ (.A1(_11618_),
    .A2(_11619_),
    .B(_11514_),
    .ZN(_11620_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20543_ (.A1(_11325_),
    .A2(_15726_),
    .Z(_11621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20544_ (.A1(net1),
    .A2(_11325_),
    .ZN(_11622_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20545_ (.A1(_11416_),
    .A2(_11621_),
    .A3(_11622_),
    .ZN(_11623_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20546_ (.A1(_11623_),
    .A2(_11600_),
    .Z(_11624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20547_ (.A1(_11620_),
    .A2(_11624_),
    .ZN(_11625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20548_ (.A1(_11617_),
    .A2(_11625_),
    .A3(_11390_),
    .ZN(_11626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20549_ (.A1(_11606_),
    .A2(_11626_),
    .A3(_11500_),
    .ZN(_11627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20550_ (.A1(_11366_),
    .A2(_11450_),
    .ZN(_11628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20551_ (.A1(_11399_),
    .A2(_11598_),
    .ZN(_11629_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20552_ (.A1(_11396_),
    .A2(_11628_),
    .B(_11629_),
    .C(_11374_),
    .ZN(_11630_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20553_ (.A1(_11424_),
    .A2(_11288_),
    .Z(_11631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20554_ (.A1(_11631_),
    .A2(_11559_),
    .ZN(_11632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20555_ (.A1(_11238_),
    .A2(_15709_),
    .ZN(_11633_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20556_ (.A1(_11356_),
    .A2(_11633_),
    .A3(_11450_),
    .ZN(_11634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20557_ (.A1(_11632_),
    .A2(_11634_),
    .ZN(_11635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20558_ (.A1(_11635_),
    .A2(_11335_),
    .B(_11422_),
    .ZN(_11636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20559_ (.A1(_11630_),
    .A2(_11636_),
    .B(_11526_),
    .ZN(_11637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20560_ (.A1(_11356_),
    .A2(_11490_),
    .A3(_11404_),
    .ZN(_11638_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20561_ (.A1(_11638_),
    .A2(_11541_),
    .B(_11318_),
    .ZN(_11639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20562_ (.I(_11481_),
    .ZN(_11640_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20563_ (.A1(_11639_),
    .A2(_11640_),
    .Z(_11641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20564_ (.I(_11618_),
    .ZN(_11642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20565_ (.A1(_11532_),
    .A2(_11325_),
    .ZN(_11643_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20566_ (.I(_11502_),
    .ZN(_11644_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20567_ (.A1(_11644_),
    .A2(_11643_),
    .ZN(_11645_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _20568_ (.I(_11333_),
    .Z(_11646_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20569_ (.A1(_11642_),
    .A2(_11645_),
    .B(_11646_),
    .ZN(_11647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20570_ (.A1(_11641_),
    .A2(_11647_),
    .ZN(_11648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20571_ (.A1(_11648_),
    .A2(_11354_),
    .ZN(_11649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20572_ (.A1(_11637_),
    .A2(_11649_),
    .ZN(_11650_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20573_ (.A1(_11473_),
    .A2(_11325_),
    .Z(_11651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20574_ (.A1(_11651_),
    .A2(_11429_),
    .ZN(_11652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20575_ (.A1(_11591_),
    .A2(_11293_),
    .ZN(_11653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20576_ (.A1(_11652_),
    .A2(_11653_),
    .B(_11600_),
    .ZN(_11654_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20577_ (.I(_11425_),
    .ZN(_11655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20578_ (.A1(_11357_),
    .A2(_11655_),
    .B(_11451_),
    .ZN(_11656_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20579_ (.A1(_11559_),
    .A2(_11450_),
    .A3(_11493_),
    .Z(_11657_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20580_ (.A1(_11656_),
    .A2(_11657_),
    .ZN(_11658_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20581_ (.A1(_11654_),
    .A2(_11658_),
    .B(_11377_),
    .ZN(_11659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20582_ (.A1(_11318_),
    .A2(_11490_),
    .ZN(_11660_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20583_ (.A1(_11494_),
    .A2(_11660_),
    .ZN(_11661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20584_ (.A1(net42),
    .A2(_11328_),
    .Z(_11662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20585_ (.A1(_11662_),
    .A2(_15723_),
    .ZN(_11663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20586_ (.A1(_11661_),
    .A2(_11663_),
    .B(_11376_),
    .ZN(_11664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20587_ (.A1(_11495_),
    .A2(_11451_),
    .Z(_11665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20588_ (.A1(_11425_),
    .A2(_11506_),
    .ZN(_11666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20589_ (.A1(_11638_),
    .A2(_11666_),
    .ZN(_11667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20590_ (.A1(_11665_),
    .A2(_11667_),
    .ZN(_11668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20591_ (.A1(_11664_),
    .A2(_11668_),
    .B(_11433_),
    .ZN(_11669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20592_ (.A1(_11659_),
    .A2(_11669_),
    .B(_11500_),
    .ZN(_11670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20593_ (.A1(_11650_),
    .A2(_11670_),
    .ZN(_11671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20594_ (.A1(_11627_),
    .A2(_11671_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20595_ (.A1(_11363_),
    .A2(_11370_),
    .Z(_11672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20596_ (.A1(_11588_),
    .A2(_11672_),
    .ZN(_11673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20597_ (.A1(_11518_),
    .A2(_15723_),
    .ZN(_11674_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20598_ (.I(_11516_),
    .ZN(_11675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20599_ (.A1(_11674_),
    .A2(_11675_),
    .ZN(_11676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20600_ (.A1(_11673_),
    .A2(_11676_),
    .A3(_11427_),
    .ZN(_11677_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20601_ (.I(_11245_),
    .ZN(_11678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20602_ (.A1(_11367_),
    .A2(_11678_),
    .ZN(_11679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20603_ (.A1(_11364_),
    .A2(_11679_),
    .A3(_11600_),
    .ZN(_11680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20604_ (.A1(_11677_),
    .A2(_11680_),
    .ZN(_11681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20605_ (.A1(_11681_),
    .A2(_11377_),
    .ZN(_11682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20606_ (.A1(_11318_),
    .A2(_11363_),
    .ZN(_11683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20607_ (.I(_11359_),
    .ZN(_11684_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20608_ (.A1(_11683_),
    .A2(_11684_),
    .ZN(_11685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20609_ (.A1(_11685_),
    .A2(_11408_),
    .B(_11376_),
    .ZN(_11686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20610_ (.A1(_11651_),
    .A2(_11424_),
    .ZN(_11687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20611_ (.A1(_11504_),
    .A2(_11687_),
    .ZN(_11688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20612_ (.A1(_11686_),
    .A2(_11688_),
    .B(_11433_),
    .ZN(_11689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20613_ (.A1(_11682_),
    .A2(_11689_),
    .B(_11442_),
    .ZN(_11690_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20614_ (.A1(_11672_),
    .A2(_11450_),
    .ZN(_11691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20615_ (.A1(_11327_),
    .A2(_11247_),
    .B(_11506_),
    .ZN(_11692_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20616_ (.A1(_11691_),
    .A2(_11427_),
    .A3(_11692_),
    .Z(_11693_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20617_ (.I(_11328_),
    .Z(_11694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20618_ (.A1(_11455_),
    .A2(_11395_),
    .A3(_11694_),
    .ZN(_11695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20619_ (.A1(_11632_),
    .A2(_11319_),
    .A3(_11695_),
    .ZN(_11696_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20620_ (.A1(_11693_),
    .A2(_11377_),
    .A3(_11696_),
    .ZN(_11697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20621_ (.A1(_11358_),
    .A2(_11537_),
    .Z(_11698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20622_ (.I(_11327_),
    .ZN(_11699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20623_ (.A1(_11699_),
    .A2(_11362_),
    .Z(_11700_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20624_ (.A1(_11698_),
    .A2(_11700_),
    .B(_11335_),
    .ZN(_11701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20625_ (.A1(_11358_),
    .A2(_11361_),
    .ZN(_11702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20626_ (.A1(_11298_),
    .A2(_11559_),
    .ZN(_11703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20627_ (.A1(_11702_),
    .A2(_11703_),
    .A3(_11374_),
    .ZN(_11704_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20628_ (.A1(_11701_),
    .A2(_11704_),
    .A3(_11354_),
    .ZN(_11705_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20629_ (.A1(_11697_),
    .A2(_11705_),
    .A3(_11390_),
    .ZN(_11706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20630_ (.A1(_11690_),
    .A2(_11706_),
    .ZN(_11707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20631_ (.I(_11493_),
    .ZN(_11708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20632_ (.A1(_11708_),
    .A2(_11694_),
    .B(_11353_),
    .ZN(_11709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20633_ (.A1(_11652_),
    .A2(_11709_),
    .B(_11600_),
    .ZN(_11710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20634_ (.A1(_15723_),
    .A2(_11607_),
    .ZN(_11711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20635_ (.A1(_11711_),
    .A2(_11328_),
    .ZN(_11712_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20636_ (.A1(_11712_),
    .A2(_11644_),
    .Z(_11713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20637_ (.A1(_11564_),
    .A2(_11293_),
    .ZN(_11714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20638_ (.A1(_11713_),
    .A2(_11714_),
    .A3(_11422_),
    .ZN(_11715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20639_ (.A1(_11710_),
    .A2(_11715_),
    .B(_11526_),
    .ZN(_11716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20640_ (.I(_11326_),
    .ZN(_11717_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20641_ (.A1(_11717_),
    .A2(_11376_),
    .B1(_11372_),
    .B2(_11462_),
    .ZN(_11718_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20642_ (.I(_11453_),
    .ZN(_11719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20643_ (.A1(_11468_),
    .A2(_11719_),
    .ZN(_11720_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20644_ (.A1(_11720_),
    .A2(_11700_),
    .B(_11353_),
    .ZN(_11721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20645_ (.A1(_11718_),
    .A2(_11721_),
    .ZN(_11722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20646_ (.A1(_11722_),
    .A2(_11335_),
    .ZN(_11723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20647_ (.A1(_11716_),
    .A2(_11723_),
    .B(_11500_),
    .ZN(_11724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20648_ (.A1(_11475_),
    .A2(_11711_),
    .ZN(_11725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20649_ (.A1(_11583_),
    .A2(_11725_),
    .B(_11600_),
    .ZN(_11726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20650_ (.I(_11656_),
    .ZN(_11727_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20651_ (.A1(_11726_),
    .A2(_11727_),
    .B(_11524_),
    .ZN(_11728_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20652_ (.A1(_11393_),
    .A2(_11708_),
    .B(_11450_),
    .ZN(_11729_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _20653_ (.I(_11334_),
    .Z(_11730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20654_ (.A1(_11426_),
    .A2(_11598_),
    .ZN(_11731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20655_ (.A1(_11729_),
    .A2(_11730_),
    .A3(_11731_),
    .ZN(_11732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20656_ (.A1(_11452_),
    .A2(_11530_),
    .ZN(_11733_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20657_ (.A1(_11732_),
    .A2(_11733_),
    .A3(_11377_),
    .ZN(_11734_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20658_ (.A1(_11728_),
    .A2(_11526_),
    .A3(_11734_),
    .ZN(_11735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20659_ (.A1(_11724_),
    .A2(_11735_),
    .ZN(_11736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20660_ (.A1(_11707_),
    .A2(_11736_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20661_ (.I(_11559_),
    .ZN(_11737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20662_ (.A1(_11466_),
    .A2(_11694_),
    .ZN(_11738_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20663_ (.A1(_11645_),
    .A2(_11427_),
    .ZN(_11739_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20664_ (.A1(_11737_),
    .A2(_11738_),
    .B(_11739_),
    .ZN(_11740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20665_ (.I(_11554_),
    .ZN(_11741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20666_ (.A1(_11741_),
    .A2(_11417_),
    .Z(_11742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20667_ (.A1(_11662_),
    .A2(_15730_),
    .ZN(_11743_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20668_ (.A1(_11542_),
    .A2(_11742_),
    .A3(_11743_),
    .ZN(_11744_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20669_ (.A1(_11740_),
    .A2(_11744_),
    .A3(_11354_),
    .ZN(_11745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20670_ (.A1(_11557_),
    .A2(_11493_),
    .Z(_11746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20671_ (.A1(_11492_),
    .A2(_11746_),
    .B(_11422_),
    .ZN(_11747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20672_ (.A1(_11544_),
    .A2(_11290_),
    .ZN(_11748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20673_ (.A1(_11476_),
    .A2(_11748_),
    .A3(_11319_),
    .ZN(_11749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20674_ (.A1(_11747_),
    .A2(_11749_),
    .B(_11526_),
    .ZN(_11750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20675_ (.A1(_11745_),
    .A2(_11750_),
    .ZN(_11751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20676_ (.A1(_11559_),
    .A2(_11356_),
    .ZN(_11752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20677_ (.A1(_11752_),
    .A2(_11372_),
    .ZN(_11753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20678_ (.A1(_11753_),
    .A2(_11575_),
    .A3(_11319_),
    .ZN(_11754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20679_ (.A1(_11451_),
    .A2(_11403_),
    .Z(_11755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20680_ (.A1(_11755_),
    .A2(_11474_),
    .B(_11422_),
    .ZN(_11756_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20681_ (.A1(_11754_),
    .A2(_11756_),
    .B(_11433_),
    .ZN(_11757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20682_ (.A1(_11602_),
    .A2(_11577_),
    .A3(_11319_),
    .ZN(_11758_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20683_ (.A1(_11400_),
    .A2(_11518_),
    .A3(_11397_),
    .ZN(_11759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20684_ (.A1(_11400_),
    .A2(_11694_),
    .A3(_11299_),
    .ZN(_11760_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20685_ (.A1(_11759_),
    .A2(_11760_),
    .A3(_11730_),
    .ZN(_11761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20686_ (.A1(_11758_),
    .A2(_11761_),
    .A3(_11354_),
    .ZN(_11762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20687_ (.A1(_11757_),
    .A2(_11762_),
    .ZN(_11763_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20688_ (.A1(_11751_),
    .A2(_11763_),
    .A3(_11500_),
    .ZN(_11764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20689_ (.A1(_11361_),
    .A2(_11559_),
    .A3(_11290_),
    .ZN(_11765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20690_ (.A1(_11475_),
    .A2(_11356_),
    .ZN(_11766_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20691_ (.A1(_11765_),
    .A2(_11766_),
    .A3(_11730_),
    .ZN(_11767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20692_ (.A1(_11486_),
    .A2(_11364_),
    .A3(_11374_),
    .ZN(_11768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20693_ (.A1(_11767_),
    .A2(_11768_),
    .A3(_11524_),
    .ZN(_11769_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20694_ (.A1(_11289_),
    .A2(_15723_),
    .Z(_11770_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20695_ (.A1(_11770_),
    .A2(_11361_),
    .B(_11417_),
    .ZN(_11771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20696_ (.A1(_11475_),
    .A2(_11400_),
    .ZN(_11772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20697_ (.A1(_11771_),
    .A2(_11772_),
    .ZN(_11773_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20698_ (.I(_15719_),
    .ZN(_11774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20699_ (.A1(_11289_),
    .A2(_11774_),
    .Z(_11775_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20700_ (.A1(_11591_),
    .A2(_11646_),
    .A3(_11775_),
    .Z(_11776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20701_ (.A1(_11773_),
    .A2(_11776_),
    .A3(_11514_),
    .ZN(_11777_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20702_ (.A1(_11769_),
    .A2(_11390_),
    .A3(_11777_),
    .ZN(_11778_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20703_ (.A1(_11730_),
    .A2(_11560_),
    .A3(_11613_),
    .A4(_11323_),
    .ZN(_11779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20704_ (.A1(_11358_),
    .A2(_11502_),
    .ZN(_11780_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20705_ (.A1(_11528_),
    .A2(_11646_),
    .ZN(_11781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20706_ (.A1(_11780_),
    .A2(_11781_),
    .B(_11376_),
    .ZN(_11782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20707_ (.A1(_11779_),
    .A2(_11782_),
    .ZN(_11783_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20708_ (.A1(_11643_),
    .A2(_11556_),
    .Z(_11784_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20709_ (.A1(_11413_),
    .A2(_11784_),
    .A3(_11374_),
    .ZN(_11785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20710_ (.A1(_11458_),
    .A2(_11289_),
    .ZN(_11786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20711_ (.A1(_11786_),
    .A2(_11334_),
    .Z(_11787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20712_ (.A1(_11787_),
    .A2(_11628_),
    .B(_11353_),
    .ZN(_11788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20713_ (.A1(_11785_),
    .A2(_11788_),
    .ZN(_11789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20714_ (.A1(_11783_),
    .A2(_11789_),
    .A3(_11526_),
    .ZN(_11790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20715_ (.A1(_11778_),
    .A2(_11790_),
    .A3(_11442_),
    .ZN(_11791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20716_ (.A1(_11764_),
    .A2(_11791_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20717_ (.A1(_11674_),
    .A2(_11450_),
    .A3(_11678_),
    .Z(_11792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20718_ (.A1(_11564_),
    .A2(_11518_),
    .Z(_11793_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20719_ (.A1(_11792_),
    .A2(_11793_),
    .B(_11335_),
    .ZN(_11794_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20720_ (.A1(_11662_),
    .A2(_11646_),
    .ZN(_11795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20721_ (.A1(_11759_),
    .A2(_11795_),
    .B(_11524_),
    .ZN(_11796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20722_ (.A1(_11794_),
    .A2(_11796_),
    .ZN(_11797_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20723_ (.A1(_11786_),
    .A2(_11719_),
    .ZN(_11798_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20724_ (.I(_11557_),
    .ZN(_11799_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20725_ (.A1(_11798_),
    .A2(_11799_),
    .B(_11646_),
    .ZN(_11800_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20726_ (.A1(_11297_),
    .A2(_11485_),
    .B(_11666_),
    .C(_11427_),
    .ZN(_11801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20727_ (.A1(_11800_),
    .A2(_11801_),
    .ZN(_11802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20728_ (.A1(_11802_),
    .A2(_11354_),
    .ZN(_11803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20729_ (.A1(_11797_),
    .A2(_11390_),
    .A3(_11803_),
    .ZN(_11804_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20730_ (.A1(_11367_),
    .A2(_11646_),
    .ZN(_11805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20731_ (.A1(_11729_),
    .A2(_11805_),
    .B(_11514_),
    .ZN(_11806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20732_ (.A1(_11528_),
    .A2(_11361_),
    .ZN(_11807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20733_ (.A1(_11807_),
    .A2(_11730_),
    .A3(_11643_),
    .ZN(_11808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20734_ (.A1(_11806_),
    .A2(_11808_),
    .B(_11433_),
    .ZN(_11809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20735_ (.A1(_11651_),
    .A2(_11466_),
    .ZN(_11810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20736_ (.A1(_11372_),
    .A2(net979),
    .ZN(_11811_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20737_ (.A1(_11464_),
    .A2(_11810_),
    .A3(_11811_),
    .ZN(_11812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20738_ (.A1(_11503_),
    .A2(_11532_),
    .ZN(_11813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20739_ (.A1(_11407_),
    .A2(_11813_),
    .A3(_11374_),
    .ZN(_11814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20740_ (.A1(_11812_),
    .A2(_11814_),
    .A3(_11377_),
    .ZN(_11815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20741_ (.A1(_11809_),
    .A2(_11815_),
    .B(_11442_),
    .ZN(_11816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20742_ (.A1(_11804_),
    .A2(_11816_),
    .ZN(_11817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20743_ (.I(_11503_),
    .ZN(_11818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20744_ (.A1(_11492_),
    .A2(_11818_),
    .B(_11524_),
    .ZN(_11819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20745_ (.A1(_11573_),
    .A2(_11290_),
    .ZN(_11820_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20746_ (.A1(_11820_),
    .A2(_11319_),
    .A3(_11712_),
    .ZN(_11821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20747_ (.A1(_11819_),
    .A2(_11821_),
    .ZN(_11822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20748_ (.A1(_11412_),
    .A2(_11598_),
    .ZN(_11823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20749_ (.A1(_11244_),
    .A2(_11694_),
    .B(_11451_),
    .ZN(_11824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20750_ (.A1(_11823_),
    .A2(_11824_),
    .B(_11514_),
    .ZN(_11825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20751_ (.A1(_11631_),
    .A2(_11502_),
    .ZN(_11826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20752_ (.A1(_11298_),
    .A2(_11467_),
    .ZN(_11827_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20753_ (.A1(_11826_),
    .A2(_11827_),
    .A3(_11730_),
    .ZN(_11828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20754_ (.A1(_11828_),
    .A2(_11825_),
    .ZN(_11829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20755_ (.A1(_11822_),
    .A2(_11829_),
    .A3(_11390_),
    .ZN(_11830_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20756_ (.A1(_11409_),
    .A2(_11417_),
    .Z(_11831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20757_ (.A1(_11360_),
    .A2(_11831_),
    .B(_11422_),
    .ZN(_11832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20758_ (.A1(_11651_),
    .A2(_11400_),
    .ZN(_11833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20759_ (.A1(_11298_),
    .A2(_11399_),
    .ZN(_11834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20760_ (.A1(_11833_),
    .A2(_11834_),
    .A3(_11600_),
    .ZN(_11835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20761_ (.A1(_11835_),
    .A2(_11832_),
    .B(_11433_),
    .ZN(_11836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20762_ (.A1(_11245_),
    .A2(_11694_),
    .B(_11417_),
    .ZN(_11837_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20763_ (.A1(_11823_),
    .A2(_11644_),
    .B(_11837_),
    .ZN(_11838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20764_ (.A1(_11540_),
    .A2(_11598_),
    .ZN(_11839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20765_ (.A1(_11413_),
    .A2(_11374_),
    .A3(_11839_),
    .ZN(_11840_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20766_ (.A1(_11838_),
    .A2(_11840_),
    .A3(_11524_),
    .ZN(_11841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20767_ (.A1(_11836_),
    .A2(_11841_),
    .ZN(_11842_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20768_ (.A1(_11842_),
    .A2(_11830_),
    .A3(_11442_),
    .ZN(_11843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20769_ (.A1(_11843_),
    .A2(_11817_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20770_ (.A1(_15724_),
    .A2(_15733_),
    .Z(_11844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20771_ (.A1(_11506_),
    .A2(_11844_),
    .ZN(_11845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20772_ (.A1(_11845_),
    .A2(_11417_),
    .ZN(_11846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20773_ (.A1(_11588_),
    .A2(_11361_),
    .B(_11846_),
    .ZN(_11847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20774_ (.A1(_11613_),
    .A2(_11451_),
    .ZN(_11848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20775_ (.A1(_11633_),
    .A2(_11493_),
    .B(_11397_),
    .ZN(_11849_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20776_ (.A1(_11848_),
    .A2(_11849_),
    .ZN(_11850_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20777_ (.A1(_11847_),
    .A2(_11850_),
    .B(_11388_),
    .ZN(_11851_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20778_ (.I(_11399_),
    .ZN(_11852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20779_ (.A1(_11400_),
    .A2(_11362_),
    .ZN(_11853_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20780_ (.A1(_11852_),
    .A2(_11853_),
    .B(_11786_),
    .ZN(_11854_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20781_ (.I(_11424_),
    .ZN(_11855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20782_ (.A1(_11855_),
    .A2(_11397_),
    .B(_11334_),
    .ZN(_11856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20783_ (.A1(_11854_),
    .A2(_11856_),
    .ZN(_11857_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20784_ (.A1(_11326_),
    .A2(_11334_),
    .Z(_11858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20785_ (.A1(_11623_),
    .A2(_11858_),
    .B(_11388_),
    .ZN(_11859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20786_ (.A1(_11859_),
    .A2(_11857_),
    .ZN(_11860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20787_ (.A1(_11851_),
    .A2(_11860_),
    .ZN(_11861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20788_ (.A1(_11861_),
    .A2(_11377_),
    .ZN(_11862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20789_ (.A1(_11473_),
    .A2(_11395_),
    .A3(_11506_),
    .ZN(_11863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20790_ (.A1(_11528_),
    .A2(_11518_),
    .ZN(_11864_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20791_ (.A1(_11863_),
    .A2(_11864_),
    .A3(_11463_),
    .ZN(_11865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20792_ (.A1(_11865_),
    .A2(_11374_),
    .ZN(_11866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20793_ (.A1(_11411_),
    .A2(_11289_),
    .Z(_11867_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20794_ (.A1(_11445_),
    .A2(_11867_),
    .ZN(_11868_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20795_ (.A1(_11450_),
    .A2(_11490_),
    .A3(_11633_),
    .A4(_11493_),
    .ZN(_11869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20796_ (.A1(_11868_),
    .A2(_11869_),
    .ZN(_11870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20797_ (.A1(_11866_),
    .A2(_11870_),
    .ZN(_11871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20798_ (.A1(_11871_),
    .A2(_11526_),
    .ZN(_11872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20799_ (.A1(_11245_),
    .A2(_11598_),
    .B(_11427_),
    .ZN(_11873_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20800_ (.A1(_11411_),
    .A2(net1),
    .B(_11694_),
    .ZN(_11874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20801_ (.A1(_11873_),
    .A2(_11874_),
    .B(_11388_),
    .ZN(_11875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20802_ (.A1(_11466_),
    .A2(_11372_),
    .A3(_11363_),
    .ZN(_11876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20803_ (.A1(_11675_),
    .A2(_11711_),
    .B(_11646_),
    .ZN(_11877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20804_ (.A1(_11876_),
    .A2(_11877_),
    .ZN(_11878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20805_ (.A1(_11875_),
    .A2(_11878_),
    .B(_11377_),
    .ZN(_11879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20806_ (.A1(_11872_),
    .A2(_11879_),
    .ZN(_11880_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20807_ (.A1(_11862_),
    .A2(_11880_),
    .A3(_11500_),
    .ZN(_11881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20808_ (.A1(_11855_),
    .A2(_11818_),
    .B(_11553_),
    .ZN(_11882_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20809_ (.I(_15725_),
    .ZN(_11883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20810_ (.A1(_11883_),
    .A2(_11694_),
    .B(_11451_),
    .ZN(_11884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20811_ (.A1(_11833_),
    .A2(_11884_),
    .ZN(_11885_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20812_ (.A1(_11882_),
    .A2(_11377_),
    .A3(_11885_),
    .ZN(_11886_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20813_ (.A1(_11474_),
    .A2(_11541_),
    .B(_11468_),
    .ZN(_11887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20814_ (.A1(_11887_),
    .A2(_11600_),
    .ZN(_11888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20815_ (.A1(_11888_),
    .A2(_11639_),
    .ZN(_11889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20816_ (.A1(_11889_),
    .A2(_11354_),
    .ZN(_11890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20817_ (.A1(_11886_),
    .A2(_11890_),
    .A3(_11390_),
    .ZN(_11891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20818_ (.A1(_11538_),
    .A2(_11431_),
    .ZN(_11892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20819_ (.A1(_11729_),
    .A2(_11856_),
    .ZN(_11893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20820_ (.A1(_11892_),
    .A2(_11893_),
    .A3(_11524_),
    .ZN(_11894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20821_ (.A1(_11685_),
    .A2(_11622_),
    .B(_11353_),
    .ZN(_11895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20822_ (.A1(_11359_),
    .A2(_11694_),
    .A3(_11363_),
    .ZN(_11896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20823_ (.A1(_11392_),
    .A2(_11543_),
    .ZN(_11897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20824_ (.A1(_11897_),
    .A2(_11598_),
    .ZN(_11898_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20825_ (.A1(_11896_),
    .A2(_11898_),
    .A3(_11600_),
    .ZN(_11899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20826_ (.A1(_11895_),
    .A2(_11899_),
    .ZN(_11900_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20827_ (.A1(_11894_),
    .A2(_11900_),
    .A3(_11526_),
    .ZN(_11901_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20828_ (.A1(_11891_),
    .A2(_11901_),
    .A3(_11442_),
    .ZN(_11902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20829_ (.A1(_11881_),
    .A2(_11902_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20830_ (.A1(_11589_),
    .A2(_11319_),
    .A3(_11863_),
    .ZN(_11903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20831_ (.A1(_11544_),
    .A2(_11372_),
    .ZN(_11904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20832_ (.A1(_11714_),
    .A2(_11904_),
    .A3(_11730_),
    .ZN(_11905_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20833_ (.A1(_11903_),
    .A2(_11354_),
    .A3(_11905_),
    .ZN(_11906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20834_ (.A1(_11552_),
    .A2(_11506_),
    .ZN(_11907_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20835_ (.A1(_11864_),
    .A2(_11907_),
    .A3(_11741_),
    .Z(_11908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20836_ (.A1(_11908_),
    .A2(_11771_),
    .ZN(_11909_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20837_ (.A1(_11568_),
    .A2(_11646_),
    .ZN(_11910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20838_ (.A1(_11910_),
    .A2(_11772_),
    .B(_11422_),
    .ZN(_11911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20839_ (.A1(_11909_),
    .A2(_11911_),
    .ZN(_11912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20840_ (.A1(_11906_),
    .A2(_11912_),
    .A3(_11526_),
    .ZN(_11913_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20841_ (.A1(_11417_),
    .A2(_11326_),
    .Z(_11914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20842_ (.A1(_11505_),
    .A2(_11372_),
    .ZN(_11915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20843_ (.A1(_11914_),
    .A2(_11915_),
    .B(_11514_),
    .ZN(_11916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20844_ (.A1(_11631_),
    .A2(_11366_),
    .ZN(_11917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20845_ (.A1(_11917_),
    .A2(_11738_),
    .A3(_11730_),
    .ZN(_11918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20846_ (.A1(_11916_),
    .A2(_11918_),
    .B(_11526_),
    .ZN(_11919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20847_ (.A1(_11719_),
    .A2(_11290_),
    .B(_11646_),
    .ZN(_11920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20848_ (.A1(_11920_),
    .A2(_11602_),
    .A3(_11759_),
    .ZN(_11921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20849_ (.A1(_11397_),
    .A2(_15714_),
    .ZN(_11922_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20850_ (.A1(_11752_),
    .A2(_11290_),
    .B(_11600_),
    .C(_11922_),
    .ZN(_11923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20851_ (.A1(_11921_),
    .A2(_11923_),
    .A3(_11377_),
    .ZN(_11924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20852_ (.A1(_11924_),
    .A2(_11919_),
    .ZN(_11925_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20853_ (.A1(_11925_),
    .A2(_11442_),
    .A3(_11913_),
    .ZN(_11926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20854_ (.A1(_11774_),
    .A2(_11694_),
    .B(_11451_),
    .ZN(_11927_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20855_ (.A1(_11633_),
    .A2(_11404_),
    .Z(_11928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20856_ (.A1(_11927_),
    .A2(_11928_),
    .B(_11353_),
    .ZN(_11929_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20857_ (.I(_11867_),
    .ZN(_11930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20858_ (.A1(_11622_),
    .A2(_11334_),
    .Z(_11931_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20859_ (.A1(_11930_),
    .A2(_11560_),
    .A3(_11931_),
    .ZN(_11932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20860_ (.A1(_11929_),
    .A2(_11932_),
    .B(_11388_),
    .ZN(_11933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20861_ (.A1(_11564_),
    .A2(_11400_),
    .ZN(_11934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20862_ (.A1(_11596_),
    .A2(_11424_),
    .ZN(_11935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20863_ (.A1(_11934_),
    .A2(_11935_),
    .A3(_11730_),
    .ZN(_11936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20864_ (.A1(_11362_),
    .A2(_15733_),
    .Z(_11937_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20865_ (.A1(_11937_),
    .A2(_11646_),
    .ZN(_11938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20866_ (.A1(_11699_),
    .A2(_11598_),
    .ZN(_11939_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20867_ (.A1(_11938_),
    .A2(_11495_),
    .A3(_11939_),
    .ZN(_11940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20868_ (.A1(_11936_),
    .A2(_11940_),
    .A3(_11524_),
    .ZN(_11941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20869_ (.A1(_11933_),
    .A2(_11941_),
    .B(_11442_),
    .ZN(_11942_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20870_ (.A1(_11518_),
    .A2(_15730_),
    .A3(_11290_),
    .Z(_11943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20871_ (.A1(_11482_),
    .A2(_11424_),
    .ZN(_11944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20872_ (.A1(_11614_),
    .A2(_11944_),
    .ZN(_11945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20873_ (.A1(_11393_),
    .A2(_11598_),
    .ZN(_11946_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20874_ (.A1(_11725_),
    .A2(_11931_),
    .A3(_11946_),
    .ZN(_11947_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20875_ (.A1(_11943_),
    .A2(_11945_),
    .B(_11947_),
    .C(_11514_),
    .ZN(_11948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20876_ (.A1(_11318_),
    .A2(_11247_),
    .Z(_11949_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20877_ (.A1(_11949_),
    .A2(_11928_),
    .Z(_11950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20878_ (.A1(_11528_),
    .A2(net1),
    .ZN(_11951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20879_ (.A1(_11950_),
    .A2(_11951_),
    .B(_11514_),
    .ZN(_11952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20880_ (.A1(_11588_),
    .A2(_11361_),
    .ZN(_11953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20881_ (.A1(_11290_),
    .A2(_15712_),
    .ZN(_11954_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20882_ (.A1(_11953_),
    .A2(_11954_),
    .A3(_11730_),
    .ZN(_11955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20883_ (.A1(_11952_),
    .A2(_11955_),
    .B(_11433_),
    .ZN(_11956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20884_ (.A1(_11948_),
    .A2(_11956_),
    .ZN(_11957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20885_ (.A1(_11942_),
    .A2(_11957_),
    .ZN(_11958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20886_ (.A1(_11926_),
    .A2(_11958_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20887_ (.I(\sa20_sub[1] ),
    .ZN(_11959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20888_ (.I(\sa31_sub[1] ),
    .ZN(_11960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20889_ (.A1(_11960_),
    .A2(_11959_),
    .ZN(_11961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20890_ (.A1(\sa20_sub[1] ),
    .A2(\sa31_sub[1] ),
    .ZN(_11962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20891_ (.A1(_11962_),
    .A2(_11961_),
    .ZN(_11963_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20892_ (.I(_11963_),
    .ZN(_11964_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20893_ (.I(\sa02_sr[7] ),
    .ZN(_11965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20894_ (.I(\sa02_sr[0] ),
    .ZN(_11966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20895_ (.A1(_11965_),
    .A2(_11966_),
    .ZN(_11967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20896_ (.A1(\sa02_sr[7] ),
    .A2(\sa02_sr[0] ),
    .ZN(_11968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20897_ (.A1(_11967_),
    .A2(_11968_),
    .ZN(_11969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20898_ (.A1(_11964_),
    .A2(_11969_),
    .ZN(_11970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20899_ (.A1(_11966_),
    .A2(\sa02_sr[7] ),
    .ZN(_11971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20900_ (.A1(_11965_),
    .A2(\sa02_sr[0] ),
    .ZN(_11972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20901_ (.A1(_11971_),
    .A2(_11972_),
    .ZN(_11973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20902_ (.A1(_11973_),
    .A2(_11963_),
    .ZN(_11974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20903_ (.A1(_11974_),
    .A2(_11970_),
    .ZN(_11975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20904_ (.I(_11975_),
    .ZN(_11976_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20905_ (.A1(\sa12_sr[7] ),
    .A2(\sa12_sr[0] ),
    .Z(_11977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20906_ (.I(\sa12_sr[1] ),
    .ZN(_11978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20907_ (.A1(_11977_),
    .A2(_11978_),
    .ZN(_11979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20908_ (.I(\sa12_sr[7] ),
    .ZN(_11980_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20909_ (.I(\sa12_sr[0] ),
    .ZN(_11981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20910_ (.A1(_11980_),
    .A2(_11981_),
    .ZN(_11982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20911_ (.A1(net1157),
    .A2(net1179),
    .ZN(_11983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20912_ (.A1(_11982_),
    .A2(_11983_),
    .ZN(_11984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20913_ (.A1(_11984_),
    .A2(net1190),
    .ZN(_11985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20914_ (.A1(_11979_),
    .A2(_11985_),
    .ZN(_11986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20915_ (.I(_11986_),
    .ZN(_11987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20916_ (.A1(_11987_),
    .A2(_11976_),
    .ZN(_11988_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _20917_ (.I(_10379_),
    .Z(_11989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20918_ (.A1(_11975_),
    .A2(_11986_),
    .ZN(_11990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20919_ (.A1(_11990_),
    .A2(_11989_),
    .A3(_11988_),
    .ZN(_11991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20920_ (.A1(_10586_),
    .A2(\text_in_r[57] ),
    .ZN(_11992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20921_ (.A1(_11991_),
    .A2(_11992_),
    .ZN(_11993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20922_ (.I(net622),
    .ZN(_11994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20923_ (.A1(_11993_),
    .A2(_11994_),
    .ZN(_11995_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20924_ (.A1(net1166),
    .A2(net623),
    .A3(_11992_),
    .ZN(_11996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20925_ (.A1(_11995_),
    .A2(_11996_),
    .ZN(_11997_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20926_ (.I(_11997_),
    .Z(_15743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20927_ (.A1(_11965_),
    .A2(_11980_),
    .ZN(_11998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20928_ (.A1(net1172),
    .A2(net1165),
    .ZN(_11999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20929_ (.A1(_11999_),
    .A2(_11998_),
    .ZN(_12000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20930_ (.A1(_12000_),
    .A2(net788),
    .ZN(_12001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20931_ (.I(\sa31_sub[0] ),
    .ZN(_12002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20932_ (.A1(_11998_),
    .A2(_12002_),
    .A3(_11999_),
    .ZN(_12003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20933_ (.A1(_12001_),
    .A2(_12003_),
    .ZN(_12004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20934_ (.A1(_11981_),
    .A2(\sa20_sub[0] ),
    .ZN(_12005_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20935_ (.I(\sa20_sub[0] ),
    .ZN(_12006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20936_ (.A1(_12006_),
    .A2(net1180),
    .ZN(_12007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20937_ (.A1(_12005_),
    .A2(_12007_),
    .ZN(_12008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20938_ (.A1(_12004_),
    .A2(_12008_),
    .ZN(_12009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20939_ (.I(_12008_),
    .ZN(_12010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20940_ (.A1(_12001_),
    .A2(_12003_),
    .A3(_12010_),
    .ZN(_12011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20941_ (.A1(_12009_),
    .A2(_12011_),
    .B(_10525_),
    .ZN(_12012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20942_ (.I(\text_in_r[56] ),
    .ZN(_12013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20943_ (.A1(_12013_),
    .A2(_10381_),
    .Z(_12014_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20944_ (.A1(_12012_),
    .A2(_12014_),
    .B(net488),
    .ZN(_12015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20945_ (.A1(_12009_),
    .A2(_12011_),
    .ZN(_12016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20946_ (.A1(_12016_),
    .A2(_10405_),
    .ZN(_12017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20947_ (.I(net488),
    .ZN(_12018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20948_ (.I(_12014_),
    .ZN(_12019_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20949_ (.A1(_12017_),
    .A2(_12018_),
    .A3(_12019_),
    .ZN(_12020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20950_ (.A1(_12020_),
    .A2(_12015_),
    .ZN(_15746_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20951_ (.I(\sa02_sr[1] ),
    .ZN(_12021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20952_ (.A1(_12021_),
    .A2(_11978_),
    .ZN(_12022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20953_ (.A1(\sa12_sr[1] ),
    .A2(\sa02_sr[1] ),
    .ZN(_12023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20954_ (.A1(_12022_),
    .A2(_12023_),
    .ZN(_12024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20955_ (.I(\sa20_sub[2] ),
    .ZN(_12025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20956_ (.A1(_12024_),
    .A2(_12025_),
    .ZN(_12026_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20957_ (.I(\sa20_sub[2] ),
    .Z(_12027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20958_ (.A1(_12022_),
    .A2(_12027_),
    .A3(_12023_),
    .ZN(_12028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20959_ (.A1(_12026_),
    .A2(_12028_),
    .ZN(_12029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20960_ (.I(\sa31_sub[2] ),
    .ZN(_12030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20961_ (.A1(_12030_),
    .A2(\sa12_sr[2] ),
    .ZN(_12031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20962_ (.I(\sa12_sr[2] ),
    .ZN(_12032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20963_ (.A1(_12032_),
    .A2(\sa31_sub[2] ),
    .ZN(_12033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20964_ (.A1(_12031_),
    .A2(_12033_),
    .ZN(_12034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20965_ (.I(_12034_),
    .ZN(_12035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20966_ (.A1(_12029_),
    .A2(_12035_),
    .ZN(_12036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20967_ (.A1(_12026_),
    .A2(_12028_),
    .A3(_12034_),
    .ZN(_12037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20968_ (.A1(_12036_),
    .A2(_12037_),
    .B(_10410_),
    .ZN(_12038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20969_ (.I(\text_in_r[58] ),
    .ZN(_12039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20970_ (.A1(_12039_),
    .A2(_11202_),
    .Z(_12040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20971_ (.I(net709),
    .ZN(_12041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20972_ (.A1(_12038_),
    .A2(_12040_),
    .B(_12041_),
    .ZN(_12042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20973_ (.A1(_12036_),
    .A2(_12037_),
    .ZN(_12043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20974_ (.A1(_12043_),
    .A2(_10522_),
    .ZN(_12044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20975_ (.I(_12040_),
    .ZN(_12045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20976_ (.A1(_12044_),
    .A2(net709),
    .A3(_12045_),
    .ZN(_12046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20977_ (.A1(_12042_),
    .A2(_12046_),
    .ZN(_12047_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _20978_ (.I(_12047_),
    .Z(_15762_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20979_ (.A1(_12012_),
    .A2(_12014_),
    .B(_12018_),
    .ZN(_12048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20980_ (.A1(net489),
    .A2(_12017_),
    .A3(_12019_),
    .ZN(_12049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20981_ (.A1(_12048_),
    .A2(_12049_),
    .ZN(_15737_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20982_ (.A1(_12038_),
    .A2(_12040_),
    .B(net709),
    .ZN(_12050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20983_ (.A1(_12044_),
    .A2(_12041_),
    .A3(_12045_),
    .ZN(_12051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20984_ (.A1(_12050_),
    .A2(_12051_),
    .ZN(_12052_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _20985_ (.I(_12052_),
    .Z(_15755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20986_ (.A1(_12047_),
    .A2(net1156),
    .ZN(_12053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20987_ (.I(_15753_),
    .ZN(_12054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20988_ (.A1(_12054_),
    .A2(_12052_),
    .ZN(_12055_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20989_ (.A1(\sa20_sub[3] ),
    .A2(\sa31_sub[3] ),
    .Z(_12056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20990_ (.I(\sa02_sr[2] ),
    .ZN(_12057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20991_ (.A1(_11965_),
    .A2(_12057_),
    .ZN(_12058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20992_ (.A1(net57),
    .A2(\sa02_sr[2] ),
    .ZN(_12059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20993_ (.A1(_12058_),
    .A2(_12059_),
    .ZN(_12060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20994_ (.A1(_12056_),
    .A2(_12060_),
    .ZN(_12061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20995_ (.A1(_12057_),
    .A2(net57),
    .ZN(_12062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20996_ (.A1(_11965_),
    .A2(\sa02_sr[2] ),
    .ZN(_12063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20997_ (.A1(_12062_),
    .A2(_12063_),
    .ZN(_12064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20998_ (.I(\sa20_sub[3] ),
    .ZN(_12065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20999_ (.I(\sa31_sub[3] ),
    .ZN(_12066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21000_ (.A1(_12065_),
    .A2(_12066_),
    .ZN(_12067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21001_ (.A1(\sa20_sub[3] ),
    .A2(\sa31_sub[3] ),
    .ZN(_12068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21002_ (.A1(_12067_),
    .A2(_12068_),
    .ZN(_12069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21003_ (.A1(_12064_),
    .A2(_12069_),
    .ZN(_12070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21004_ (.A1(_12061_),
    .A2(_12070_),
    .ZN(_12071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21005_ (.I(_12071_),
    .ZN(_12072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21006_ (.I(\sa12_sr[3] ),
    .ZN(_12073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21007_ (.A1(_12073_),
    .A2(net72),
    .ZN(_12074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21008_ (.A1(_11980_),
    .A2(\sa12_sr[3] ),
    .ZN(_12075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21009_ (.A1(_12074_),
    .A2(_12075_),
    .ZN(_12076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21010_ (.A1(_12076_),
    .A2(\sa12_sr[2] ),
    .ZN(_12077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21011_ (.A1(_11980_),
    .A2(_12073_),
    .ZN(_12078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21012_ (.A1(net72),
    .A2(\sa12_sr[3] ),
    .ZN(_12079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21013_ (.A1(_12078_),
    .A2(_12079_),
    .ZN(_12080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21014_ (.A1(_12080_),
    .A2(_12032_),
    .ZN(_12081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21015_ (.A1(_12077_),
    .A2(_12081_),
    .ZN(_12082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21016_ (.A1(_12072_),
    .A2(_12082_),
    .ZN(_12083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21017_ (.I(_12082_),
    .ZN(_12084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21018_ (.A1(_12084_),
    .A2(_12071_),
    .ZN(_12085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21019_ (.A1(_12083_),
    .A2(_12085_),
    .A3(_11279_),
    .ZN(_12086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21020_ (.A1(_10411_),
    .A2(\text_in_r[59] ),
    .ZN(_12087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21021_ (.A1(_12086_),
    .A2(\u0.w[2][27] ),
    .A3(_12087_),
    .ZN(_12088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21022_ (.A1(_12072_),
    .A2(_12084_),
    .ZN(_12089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21023_ (.A1(_12071_),
    .A2(_12082_),
    .ZN(_12090_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21024_ (.A1(_12089_),
    .A2(_12090_),
    .A3(_11279_),
    .ZN(_12091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21025_ (.I(\u0.w[2][27] ),
    .ZN(_12092_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21026_ (.A1(_10489_),
    .A2(\text_in_r[59] ),
    .Z(_12093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21027_ (.A1(_12091_),
    .A2(_12092_),
    .A3(_12093_),
    .ZN(_12094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21028_ (.A1(_12088_),
    .A2(_12094_),
    .ZN(_12095_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21029_ (.I(_12095_),
    .Z(_12096_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21030_ (.I(_12096_),
    .Z(_12097_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21031_ (.A1(_12053_),
    .A2(_12055_),
    .A3(_12097_),
    .Z(_12098_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21032_ (.A1(\sa12_sr[4] ),
    .A2(\sa31_sub[4] ),
    .Z(_12099_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21033_ (.A1(_12099_),
    .A2(_12076_),
    .Z(_12100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21034_ (.A1(_12099_),
    .A2(_12076_),
    .ZN(_12101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21035_ (.A1(_12100_),
    .A2(_12101_),
    .ZN(_12102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21036_ (.I(_12102_),
    .ZN(_12103_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21037_ (.A1(net57),
    .A2(\sa02_sr[3] ),
    .Z(_12104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21038_ (.I(\sa20_sub[4] ),
    .ZN(_12105_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21039_ (.A1(_12104_),
    .A2(_12105_),
    .ZN(_12106_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21040_ (.I(_12106_),
    .ZN(_12107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21041_ (.A1(_12104_),
    .A2(_12105_),
    .ZN(_12108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21042_ (.A1(_12107_),
    .A2(_12108_),
    .ZN(_12109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21043_ (.A1(_12103_),
    .A2(_12109_),
    .ZN(_12110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21044_ (.I(_12108_),
    .ZN(_12111_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21045_ (.A1(_12111_),
    .A2(_12106_),
    .ZN(_12112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21046_ (.A1(_12112_),
    .A2(_12102_),
    .ZN(_12113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21047_ (.A1(_12110_),
    .A2(_12113_),
    .A3(_10523_),
    .ZN(_12114_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _21048_ (.I(_11203_),
    .Z(_12115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21049_ (.A1(_12115_),
    .A2(\text_in_r[60] ),
    .ZN(_12116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21050_ (.A1(_12114_),
    .A2(_12116_),
    .ZN(_12117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21051_ (.A1(_12117_),
    .A2(\u0.w[2][28] ),
    .ZN(_12118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21052_ (.I(\u0.w[2][28] ),
    .ZN(_12119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21053_ (.A1(_12114_),
    .A2(_12119_),
    .A3(_12116_),
    .ZN(_12120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21054_ (.A1(_12118_),
    .A2(_12120_),
    .ZN(_12121_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21055_ (.I(_12121_),
    .Z(_12122_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21056_ (.A1(_12098_),
    .A2(_12122_),
    .ZN(_12123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21057_ (.I(_12053_),
    .ZN(_12124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21058_ (.A1(_12124_),
    .A2(net20),
    .ZN(_12125_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21059_ (.A1(_12086_),
    .A2(_12092_),
    .A3(_12087_),
    .ZN(_12126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21060_ (.A1(_12091_),
    .A2(\u0.w[2][27] ),
    .A3(_12093_),
    .ZN(_12127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21061_ (.A1(_12126_),
    .A2(_12127_),
    .ZN(_12128_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21062_ (.I(_12128_),
    .Z(_12129_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21063_ (.I(_12129_),
    .Z(_12130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21064_ (.A1(_11993_),
    .A2(net622),
    .ZN(_12131_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21065_ (.A1(net1166),
    .A2(_11994_),
    .A3(_11992_),
    .ZN(_12132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21066_ (.A1(_12131_),
    .A2(_12132_),
    .ZN(_15738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21067_ (.A1(_15738_),
    .A2(_12052_),
    .ZN(_12133_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21068_ (.I(_12133_),
    .Z(_12134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21069_ (.A1(_12125_),
    .A2(_12130_),
    .A3(_12134_),
    .ZN(_12135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21070_ (.A1(_12123_),
    .A2(_12135_),
    .ZN(_12136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21071_ (.I(_15741_),
    .ZN(_12137_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _21072_ (.A1(_12047_),
    .A2(_12137_),
    .ZN(_12138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21073_ (.A1(_12138_),
    .A2(_12128_),
    .ZN(_12139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21074_ (.A1(_12139_),
    .A2(_12121_),
    .ZN(_12140_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21075_ (.I(_12128_),
    .Z(_12141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21076_ (.A1(net17),
    .A2(_12141_),
    .A3(_15762_),
    .ZN(_12142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21077_ (.I(_12142_),
    .ZN(_12143_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21078_ (.A1(_12140_),
    .A2(_12143_),
    .ZN(_12144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21079_ (.A1(net1150),
    .A2(net1154),
    .A3(_12052_),
    .ZN(_12145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21080_ (.A1(_12053_),
    .A2(_12096_),
    .A3(_12145_),
    .ZN(_12146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21081_ (.A1(_12144_),
    .A2(_12146_),
    .ZN(_12147_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21082_ (.A1(\sa12_sr[4] ),
    .A2(\sa02_sr[4] ),
    .Z(_12148_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21083_ (.A1(\sa20_sub[5] ),
    .A2(\sa31_sub[5] ),
    .Z(_12149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21084_ (.A1(\sa20_sub[5] ),
    .A2(\sa31_sub[5] ),
    .ZN(_12150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21085_ (.A1(_12149_),
    .A2(_12150_),
    .ZN(_12151_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21086_ (.A1(\sa12_sr[5] ),
    .A2(_12151_),
    .Z(_12152_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21087_ (.A1(_12148_),
    .A2(_12152_),
    .Z(_12153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21088_ (.I(\u0.w[2][29] ),
    .ZN(_12154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21089_ (.A1(_10587_),
    .A2(\text_in_r[61] ),
    .ZN(_12155_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _21090_ (.A1(_12153_),
    .A2(_10639_),
    .B(_12154_),
    .C(_12155_),
    .ZN(_12156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21091_ (.A1(_12153_),
    .A2(_10585_),
    .ZN(_12157_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21092_ (.A1(_11348_),
    .A2(\text_in_r[61] ),
    .Z(_12158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21093_ (.A1(_12157_),
    .A2(\u0.w[2][29] ),
    .A3(_12158_),
    .ZN(_12159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21094_ (.A1(_12156_),
    .A2(_12159_),
    .ZN(_12160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21095_ (.I(_12160_),
    .Z(_12161_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21096_ (.A1(_12136_),
    .A2(_12147_),
    .A3(_12161_),
    .ZN(_12162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21097_ (.I(_15744_),
    .ZN(_12163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21098_ (.A1(_12163_),
    .A2(_12052_),
    .ZN(_12164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21099_ (.A1(_12164_),
    .A2(_12095_),
    .ZN(_12165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21100_ (.I(_12165_),
    .ZN(_12166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21101_ (.A1(_12125_),
    .A2(_12166_),
    .ZN(_12167_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21102_ (.I(_12121_),
    .Z(_12168_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21103_ (.I(_12168_),
    .Z(_12169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21104_ (.A1(_12053_),
    .A2(_12129_),
    .Z(_12170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21105_ (.I(_12170_),
    .ZN(_12171_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21106_ (.A1(_12167_),
    .A2(_12169_),
    .A3(_12171_),
    .ZN(_12172_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21107_ (.I(_12141_),
    .Z(_12173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21108_ (.A1(_12052_),
    .A2(_15737_),
    .ZN(_12174_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21109_ (.I(_12174_),
    .Z(_12175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21110_ (.A1(_12125_),
    .A2(_12173_),
    .A3(_12175_),
    .ZN(_12176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21111_ (.A1(_12052_),
    .A2(_15740_),
    .ZN(_12177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21112_ (.A1(_12050_),
    .A2(_12051_),
    .A3(_15753_),
    .ZN(_12178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21113_ (.A1(_12177_),
    .A2(_12178_),
    .ZN(_12179_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21114_ (.I(_12096_),
    .Z(_12180_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21115_ (.I(_12121_),
    .Z(_12181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21116_ (.A1(_12179_),
    .A2(_12180_),
    .B(_12181_),
    .ZN(_12182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21117_ (.A1(_12176_),
    .A2(_12182_),
    .ZN(_12183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21118_ (.I(_12160_),
    .ZN(_12184_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21119_ (.I(_12184_),
    .Z(_12185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21120_ (.A1(_12172_),
    .A2(_12183_),
    .A3(_12185_),
    .ZN(_12186_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21121_ (.A1(\sa12_sr[5] ),
    .A2(\sa02_sr[5] ),
    .ZN(_12187_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21122_ (.A1(\sa20_sub[6] ),
    .A2(\sa31_sub[6] ),
    .Z(_12188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21123_ (.A1(\sa20_sub[6] ),
    .A2(\sa31_sub[6] ),
    .ZN(_12189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21124_ (.A1(_12188_),
    .A2(_12189_),
    .ZN(_12190_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21125_ (.A1(\sa12_sr[6] ),
    .A2(_12190_),
    .Z(_12191_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21126_ (.A1(_12187_),
    .A2(_12191_),
    .Z(_12192_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _21127_ (.I(_10431_),
    .Z(_12193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21128_ (.A1(_12193_),
    .A2(\text_in_r[62] ),
    .Z(_12194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21129_ (.A1(_12192_),
    .A2(_11348_),
    .B(_12194_),
    .ZN(_12195_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21130_ (.A1(\u0.w[2][30] ),
    .A2(_12195_),
    .Z(_12196_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21131_ (.I(_12196_),
    .Z(_12197_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21132_ (.I(_12197_),
    .ZN(_12198_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21133_ (.I(_12198_),
    .Z(_12199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21134_ (.A1(_12162_),
    .A2(_12186_),
    .A3(_12199_),
    .ZN(_12200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21135_ (.A1(_12052_),
    .A2(net1150),
    .ZN(_12201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21136_ (.A1(_12201_),
    .A2(_12141_),
    .Z(_12202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21137_ (.A1(net17),
    .A2(net71),
    .ZN(_12203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21138_ (.A1(_12202_),
    .A2(_12203_),
    .ZN(_12204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21139_ (.A1(net71),
    .A2(net1152),
    .ZN(_12205_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21140_ (.I(_12095_),
    .Z(_12206_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21141_ (.I(_12047_),
    .Z(_12207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21142_ (.A1(_12207_),
    .A2(net1150),
    .ZN(_12208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21143_ (.A1(_12208_),
    .A2(_12206_),
    .A3(_12205_),
    .ZN(_12209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21144_ (.A1(_12117_),
    .A2(_12119_),
    .ZN(_12210_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21145_ (.A1(_12114_),
    .A2(\u0.w[2][28] ),
    .A3(_12116_),
    .ZN(_12211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21146_ (.A1(_12210_),
    .A2(_12211_),
    .ZN(_12212_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21147_ (.I(_12212_),
    .Z(_12213_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21148_ (.I(_12213_),
    .Z(_12214_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21149_ (.A1(_12204_),
    .A2(_12209_),
    .A3(_12214_),
    .ZN(_12215_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _21150_ (.I(_15739_),
    .ZN(_12216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21151_ (.A1(_12207_),
    .A2(_12216_),
    .ZN(_12217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21152_ (.I(_15747_),
    .ZN(_12218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21153_ (.A1(_15755_),
    .A2(_12218_),
    .ZN(_12219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21154_ (.A1(_12217_),
    .A2(_12219_),
    .ZN(_12220_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21155_ (.I(_12206_),
    .Z(_12221_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21156_ (.I(_12213_),
    .Z(_12222_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21157_ (.A1(_12220_),
    .A2(_12221_),
    .B(_12222_),
    .ZN(_12223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21158_ (.A1(_12047_),
    .A2(net1151),
    .Z(_12224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21159_ (.A1(net20),
    .A2(_12224_),
    .ZN(_12225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21160_ (.I(_15740_),
    .ZN(_12226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21161_ (.A1(_12226_),
    .A2(_12052_),
    .ZN(_12227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21162_ (.A1(_12227_),
    .A2(_12129_),
    .Z(_12228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21163_ (.A1(net1158),
    .A2(_12228_),
    .ZN(_12229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21164_ (.A1(_12223_),
    .A2(_12229_),
    .ZN(_12230_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21165_ (.A1(_12215_),
    .A2(_12230_),
    .A3(_12185_),
    .ZN(_12231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21166_ (.A1(_12129_),
    .A2(_12226_),
    .A3(_15755_),
    .ZN(_12232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21167_ (.A1(_12226_),
    .A2(_12207_),
    .ZN(_12233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21168_ (.A1(_12096_),
    .A2(_12233_),
    .ZN(_12234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21169_ (.A1(_12142_),
    .A2(_12232_),
    .A3(_12234_),
    .ZN(_12235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21170_ (.A1(_12235_),
    .A2(_12214_),
    .ZN(_12236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21171_ (.A1(_12052_),
    .A2(_12216_),
    .ZN(_12237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21172_ (.A1(_15762_),
    .A2(_12218_),
    .ZN(_12238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21173_ (.A1(_12237_),
    .A2(_12238_),
    .ZN(_12239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21174_ (.A1(_12239_),
    .A2(_12130_),
    .ZN(_12240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21175_ (.A1(_15762_),
    .A2(_15739_),
    .ZN(_12241_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21176_ (.I(_12096_),
    .Z(_12242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21177_ (.A1(_12227_),
    .A2(_12241_),
    .A3(_12242_),
    .ZN(_12243_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21178_ (.I(_12168_),
    .Z(_12244_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21179_ (.A1(_12240_),
    .A2(_12243_),
    .A3(_12244_),
    .ZN(_12245_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21180_ (.I(_12160_),
    .Z(_12246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21181_ (.A1(_12236_),
    .A2(_12245_),
    .A3(_12246_),
    .ZN(_12247_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21182_ (.I(_12197_),
    .Z(_12248_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21183_ (.A1(_12231_),
    .A2(_12247_),
    .A3(_12248_),
    .ZN(_12249_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21184_ (.I(\sa20_sub[7] ),
    .Z(_12250_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21185_ (.I(\sa31_sub[7] ),
    .Z(_12251_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21186_ (.A1(\sa12_sr[6] ),
    .A2(\sa02_sr[6] ),
    .Z(_12252_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21187_ (.A1(net72),
    .A2(_12252_),
    .Z(_12253_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _21188_ (.A1(net49),
    .A2(net642),
    .A3(_12253_),
    .Z(_12254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21189_ (.I0(_12254_),
    .I1(\text_in_r[63] ),
    .S(_10587_),
    .Z(_12255_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21190_ (.A1(\u0.w[2][31] ),
    .A2(_12255_),
    .ZN(_12256_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21191_ (.I(_12256_),
    .Z(_12257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21192_ (.A1(_12200_),
    .A2(_12249_),
    .A3(_12257_),
    .ZN(_12258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21193_ (.A1(_12207_),
    .A2(_15744_),
    .ZN(_12259_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21194_ (.I(_12259_),
    .ZN(_12260_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21195_ (.I(_12212_),
    .Z(_12261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21196_ (.A1(_12260_),
    .A2(_12173_),
    .B(_12261_),
    .ZN(_12262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21197_ (.A1(_12146_),
    .A2(_12262_),
    .ZN(_12263_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21198_ (.A1(_12042_),
    .A2(_12046_),
    .A3(_15749_),
    .ZN(_12264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21199_ (.A1(_12259_),
    .A2(_12264_),
    .B(_12097_),
    .ZN(_12265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21200_ (.A1(_12227_),
    .A2(_12096_),
    .ZN(_12266_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21201_ (.I(_12266_),
    .ZN(_12267_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21202_ (.A1(_12265_),
    .A2(_12267_),
    .ZN(_12268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21203_ (.A1(_12268_),
    .A2(_12214_),
    .ZN(_12269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21204_ (.A1(_12263_),
    .A2(_12269_),
    .A3(_12199_),
    .ZN(_12270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21205_ (.A1(_12208_),
    .A2(_12237_),
    .ZN(_12271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21206_ (.A1(_12271_),
    .A2(_12242_),
    .B(_12261_),
    .ZN(_12272_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21207_ (.A1(_15755_),
    .A2(net71),
    .A3(net20),
    .ZN(_12273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21208_ (.A1(_12050_),
    .A2(_12051_),
    .A3(_12163_),
    .ZN(_12274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21209_ (.A1(_12273_),
    .A2(_12173_),
    .A3(_12274_),
    .ZN(_12275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21210_ (.A1(_12207_),
    .A2(_15741_),
    .Z(_12276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21211_ (.A1(_12276_),
    .A2(_12129_),
    .ZN(_12277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21212_ (.A1(_12272_),
    .A2(_12275_),
    .A3(_12277_),
    .ZN(_12278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21213_ (.A1(_12050_),
    .A2(net1161),
    .A3(_12051_),
    .ZN(_12279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21214_ (.I(_12279_),
    .ZN(_12280_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21215_ (.I(_12141_),
    .Z(_12281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21216_ (.A1(_12280_),
    .A2(_12281_),
    .B(_12121_),
    .ZN(_12282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21217_ (.A1(_12221_),
    .A2(_15760_),
    .ZN(_12283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21218_ (.A1(_12282_),
    .A2(_12283_),
    .B(_12198_),
    .ZN(_12284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21219_ (.A1(_12278_),
    .A2(_12284_),
    .ZN(_12285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21220_ (.A1(_12270_),
    .A2(_12285_),
    .A3(_12161_),
    .ZN(_12286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21221_ (.A1(_12138_),
    .A2(_12206_),
    .ZN(_12287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21222_ (.A1(_12287_),
    .A2(_12213_),
    .Z(_12288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21223_ (.A1(_12207_),
    .A2(_15747_),
    .ZN(_12289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21224_ (.A1(_12289_),
    .A2(_12141_),
    .Z(_12290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21225_ (.A1(_12290_),
    .A2(net1155),
    .ZN(_12291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21226_ (.A1(_12288_),
    .A2(_12291_),
    .B(_12198_),
    .ZN(_12292_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21227_ (.I(_12140_),
    .ZN(_12293_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21228_ (.I(_15749_),
    .ZN(_12294_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21229_ (.A1(_12050_),
    .A2(_12051_),
    .A3(_12294_),
    .ZN(_12295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21230_ (.A1(_12095_),
    .A2(_12295_),
    .Z(_12296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21231_ (.A1(_12273_),
    .A2(_12296_),
    .ZN(_12297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21232_ (.A1(_12293_),
    .A2(_12297_),
    .ZN(_12298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21233_ (.A1(_12292_),
    .A2(_12298_),
    .B(_12246_),
    .ZN(_12299_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21234_ (.A1(_12139_),
    .A2(_12165_),
    .Z(_12300_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21235_ (.I(_12217_),
    .ZN(_12301_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21236_ (.I(_12128_),
    .Z(_12302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21237_ (.A1(_12301_),
    .A2(_12302_),
    .ZN(_12303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21238_ (.A1(_12300_),
    .A2(_12303_),
    .B(_12122_),
    .ZN(_12304_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _21239_ (.I(_12201_),
    .ZN(_12305_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21240_ (.I(_12238_),
    .ZN(_12306_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21241_ (.A1(_12305_),
    .A2(_12306_),
    .B(_12242_),
    .ZN(_12307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21242_ (.A1(_15755_),
    .A2(net20),
    .ZN(_12308_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21243_ (.A1(_12308_),
    .A2(_12302_),
    .A3(_12279_),
    .ZN(_12309_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21244_ (.I(_12213_),
    .Z(_12310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21245_ (.A1(_12307_),
    .A2(_12309_),
    .B(_12310_),
    .ZN(_12311_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21246_ (.A1(_12304_),
    .A2(_12311_),
    .B(_12198_),
    .ZN(_12312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21247_ (.A1(_12299_),
    .A2(_12312_),
    .ZN(_12313_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21248_ (.I(_12257_),
    .ZN(_12314_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21249_ (.A1(_12286_),
    .A2(_12313_),
    .A3(_12314_),
    .ZN(_12315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21250_ (.A1(_12258_),
    .A2(_12315_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21251_ (.A1(_15738_),
    .A2(_12207_),
    .ZN(_12316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21252_ (.A1(_12166_),
    .A2(_12316_),
    .ZN(_12317_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21253_ (.A1(_12201_),
    .A2(_12241_),
    .A3(_12173_),
    .ZN(_12318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21254_ (.A1(_12317_),
    .A2(_12169_),
    .A3(_12318_),
    .ZN(_12319_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21255_ (.I(_12129_),
    .Z(_12320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21256_ (.A1(net1149),
    .A2(_12320_),
    .B(_12181_),
    .ZN(_12321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21257_ (.A1(_12237_),
    .A2(net1163),
    .ZN(_12322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21258_ (.A1(_12322_),
    .A2(_12180_),
    .ZN(_12323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21259_ (.A1(_12224_),
    .A2(_12281_),
    .ZN(_12324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21260_ (.A1(_12321_),
    .A2(_12323_),
    .A3(_12324_),
    .ZN(_12325_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21261_ (.I(_12184_),
    .Z(_12326_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21262_ (.A1(_12319_),
    .A2(_12325_),
    .A3(_12326_),
    .ZN(_12327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21263_ (.A1(_12170_),
    .A2(_12145_),
    .ZN(_12328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21264_ (.A1(_12266_),
    .A2(_12168_),
    .Z(_12329_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21265_ (.A1(_12329_),
    .A2(_12328_),
    .B(_12184_),
    .ZN(_12330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21266_ (.A1(_12055_),
    .A2(_12129_),
    .Z(_12331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21267_ (.A1(_12207_),
    .A2(_12137_),
    .ZN(_12332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21268_ (.A1(_12331_),
    .A2(_12332_),
    .B(_12181_),
    .ZN(_12333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21269_ (.A1(_12225_),
    .A2(_12242_),
    .A3(_12177_),
    .ZN(_12334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21270_ (.A1(_12333_),
    .A2(_12334_),
    .ZN(_12335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21271_ (.A1(_12330_),
    .A2(_12335_),
    .ZN(_12336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21272_ (.A1(_12336_),
    .A2(_12327_),
    .B(_12248_),
    .ZN(_12337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21273_ (.A1(_15743_),
    .A2(_15762_),
    .ZN(_12338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21274_ (.A1(_12202_),
    .A2(_12338_),
    .ZN(_12339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21275_ (.A1(_12339_),
    .A2(_12317_),
    .ZN(_12340_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21276_ (.A1(_12340_),
    .A2(_12246_),
    .B(_12169_),
    .ZN(_12341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21277_ (.A1(_12305_),
    .A2(net20),
    .B(_12302_),
    .ZN(_12342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21278_ (.A1(_12342_),
    .A2(_12125_),
    .ZN(_12343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21279_ (.A1(_12175_),
    .A2(_12241_),
    .A3(_12281_),
    .ZN(_12344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21280_ (.A1(_12343_),
    .A2(_12344_),
    .ZN(_12345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21281_ (.A1(_12345_),
    .A2(_12185_),
    .ZN(_12346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21282_ (.A1(_12156_),
    .A2(_12159_),
    .B(_15763_),
    .ZN(_12347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21283_ (.A1(_12347_),
    .A2(_12221_),
    .ZN(_12348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21284_ (.A1(_12290_),
    .A2(_12145_),
    .ZN(_12349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21285_ (.A1(_12348_),
    .A2(_12349_),
    .A3(_12122_),
    .ZN(_12350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21286_ (.A1(_12350_),
    .A2(_12197_),
    .ZN(_12351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21287_ (.A1(_12341_),
    .A2(_12346_),
    .B(_12351_),
    .ZN(_12352_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21288_ (.A1(_12337_),
    .A2(_12352_),
    .B(_12257_),
    .ZN(_12353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21289_ (.A1(_12207_),
    .A2(_12054_),
    .ZN(_12354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21290_ (.A1(_12354_),
    .A2(_12096_),
    .ZN(_12355_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21291_ (.I(_12355_),
    .ZN(_12356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21292_ (.A1(_12356_),
    .A2(_12134_),
    .B(_12181_),
    .ZN(_12357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21293_ (.A1(_12134_),
    .A2(_12175_),
    .ZN(_12358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21294_ (.A1(_12358_),
    .A2(_12130_),
    .ZN(_12359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21295_ (.A1(_12357_),
    .A2(_12359_),
    .ZN(_12360_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21296_ (.A1(_15755_),
    .A2(net1159),
    .Z(_12361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21297_ (.A1(_12361_),
    .A2(_12320_),
    .B(_12222_),
    .ZN(_12362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21298_ (.A1(_12334_),
    .A2(_12362_),
    .ZN(_12363_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21299_ (.A1(_12360_),
    .A2(_12363_),
    .A3(_12185_),
    .ZN(_12364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21300_ (.A1(_15743_),
    .A2(net1150),
    .ZN(_12365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21301_ (.A1(_12365_),
    .A2(_12175_),
    .ZN(_12366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21302_ (.A1(_12366_),
    .A2(_12221_),
    .ZN(_12367_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21303_ (.A1(_12141_),
    .A2(_12279_),
    .Z(_12368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21304_ (.A1(_12368_),
    .A2(_12175_),
    .ZN(_12369_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21305_ (.A1(_12367_),
    .A2(_12244_),
    .A3(_12369_),
    .ZN(_12370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21306_ (.A1(_12259_),
    .A2(net13),
    .ZN(_12371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21307_ (.A1(_12371_),
    .A2(_12221_),
    .ZN(_12372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21308_ (.A1(_12271_),
    .A2(_12320_),
    .ZN(_12373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21309_ (.A1(_12372_),
    .A2(_12373_),
    .A3(_12310_),
    .ZN(_12374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21310_ (.A1(_12370_),
    .A2(_12374_),
    .A3(_12246_),
    .ZN(_12375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21311_ (.A1(_12364_),
    .A2(_12375_),
    .A3(_12199_),
    .ZN(_12376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21312_ (.A1(_12338_),
    .A2(_12206_),
    .ZN(_12377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21313_ (.A1(_12377_),
    .A2(_12134_),
    .Z(_12378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21314_ (.A1(_12260_),
    .A2(_12281_),
    .B(_12168_),
    .ZN(_12379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21315_ (.A1(_12378_),
    .A2(_12379_),
    .B(_12184_),
    .ZN(_12380_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21316_ (.I(_12234_),
    .ZN(_12381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21317_ (.A1(_12055_),
    .A2(_12381_),
    .ZN(_12382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21318_ (.A1(_12275_),
    .A2(_12169_),
    .A3(_12382_),
    .ZN(_12383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21319_ (.A1(_12380_),
    .A2(_12383_),
    .ZN(_12384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21320_ (.A1(_12164_),
    .A2(_12128_),
    .Z(_12385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21321_ (.A1(_12385_),
    .A2(_12208_),
    .ZN(_12386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21322_ (.I(_12213_),
    .Z(_12387_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21323_ (.I(_12096_),
    .Z(_12388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21324_ (.A1(_12053_),
    .A2(_12227_),
    .A3(_12388_),
    .ZN(_12389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21325_ (.A1(_12386_),
    .A2(_12387_),
    .A3(_12389_),
    .ZN(_12390_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21326_ (.A1(_12096_),
    .A2(_12207_),
    .Z(_12391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21327_ (.A1(_12391_),
    .A2(_12205_),
    .B(_12222_),
    .ZN(_12392_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21328_ (.A1(_12308_),
    .A2(_12203_),
    .A3(_12281_),
    .ZN(_12393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21329_ (.A1(_12392_),
    .A2(_12393_),
    .ZN(_12394_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21330_ (.A1(_12390_),
    .A2(_12326_),
    .A3(_12394_),
    .ZN(_12395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21331_ (.A1(_12384_),
    .A2(_12395_),
    .A3(_12248_),
    .ZN(_12396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21332_ (.A1(_12376_),
    .A2(_12396_),
    .A3(_12314_),
    .ZN(_12397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21333_ (.A1(_12353_),
    .A2(_12397_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21334_ (.A1(net20),
    .A2(_15762_),
    .ZN(_12398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21335_ (.A1(_12274_),
    .A2(_12097_),
    .ZN(_12399_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21336_ (.A1(_12398_),
    .A2(_12399_),
    .ZN(_12400_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21337_ (.A1(_12400_),
    .A2(_12265_),
    .B(_12122_),
    .ZN(_12401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21338_ (.A1(_12264_),
    .A2(_12178_),
    .ZN(_12402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21339_ (.A1(_12402_),
    .A2(_12302_),
    .ZN(_12403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21340_ (.A1(_12175_),
    .A2(_12097_),
    .A3(_12274_),
    .ZN(_12404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21341_ (.A1(_12403_),
    .A2(_12404_),
    .ZN(_12405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21342_ (.A1(_12405_),
    .A2(_12310_),
    .ZN(_12406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21343_ (.A1(_12401_),
    .A2(_12406_),
    .A3(_12246_),
    .ZN(_12407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21344_ (.A1(_12316_),
    .A2(_12388_),
    .A3(_12264_),
    .ZN(_12408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21345_ (.A1(_12201_),
    .A2(_12302_),
    .A3(_12178_),
    .ZN(_12409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21346_ (.A1(_12408_),
    .A2(_12310_),
    .A3(_12409_),
    .ZN(_12410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21347_ (.A1(_12175_),
    .A2(_12129_),
    .A3(_12295_),
    .ZN(_12411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21348_ (.A1(_12227_),
    .A2(_12279_),
    .A3(_12206_),
    .ZN(_12412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21349_ (.A1(_12411_),
    .A2(_12412_),
    .ZN(_12413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21350_ (.A1(_12413_),
    .A2(_12122_),
    .ZN(_12414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21351_ (.A1(_12410_),
    .A2(_12414_),
    .A3(_12326_),
    .ZN(_12415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21352_ (.A1(_12407_),
    .A2(_12415_),
    .ZN(_12416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21353_ (.A1(_12416_),
    .A2(_12199_),
    .B(_12314_),
    .ZN(_12417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21354_ (.A1(_12308_),
    .A2(_12205_),
    .A3(_12206_),
    .ZN(_12418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21355_ (.A1(_12385_),
    .A2(_12354_),
    .ZN(_12419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21356_ (.A1(_12418_),
    .A2(_12419_),
    .ZN(_12420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21357_ (.A1(_12420_),
    .A2(_12310_),
    .ZN(_12421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21358_ (.A1(_12174_),
    .A2(_12274_),
    .ZN(_12422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21359_ (.A1(_12422_),
    .A2(_12097_),
    .A3(_12133_),
    .ZN(_12423_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21360_ (.A1(_12423_),
    .A2(_12122_),
    .A3(_12309_),
    .ZN(_12424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21361_ (.A1(_12421_),
    .A2(_12424_),
    .ZN(_12425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21362_ (.A1(_12425_),
    .A2(_12161_),
    .ZN(_12426_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21363_ (.A1(_12225_),
    .A2(_12221_),
    .A3(_12055_),
    .ZN(_12427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21364_ (.A1(_12125_),
    .A2(_12173_),
    .ZN(_12428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21365_ (.A1(_12427_),
    .A2(_12169_),
    .A3(_12428_),
    .ZN(_12429_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21366_ (.A1(_12305_),
    .A2(_12276_),
    .B(_12180_),
    .ZN(_12430_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21367_ (.A1(_12338_),
    .A2(_12320_),
    .A3(net13),
    .ZN(_12431_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21368_ (.A1(_12430_),
    .A2(_12431_),
    .A3(_12387_),
    .ZN(_12432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21369_ (.A1(_12429_),
    .A2(_12185_),
    .A3(_12432_),
    .ZN(_12433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21370_ (.A1(_12426_),
    .A2(_12433_),
    .A3(_12248_),
    .ZN(_12434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21371_ (.A1(_12417_),
    .A2(_12434_),
    .ZN(_12435_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21372_ (.A1(_12308_),
    .A2(_12281_),
    .A3(_12217_),
    .Z(_12436_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21373_ (.A1(_12219_),
    .A2(_12388_),
    .A3(_12279_),
    .Z(_12437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21374_ (.A1(_12436_),
    .A2(_12437_),
    .B(_12214_),
    .ZN(_12438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21375_ (.A1(_12308_),
    .A2(_12203_),
    .A3(_12388_),
    .ZN(_12439_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21376_ (.A1(_12388_),
    .A2(_15763_),
    .Z(_12440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21377_ (.A1(_12439_),
    .A2(_12169_),
    .A3(_12440_),
    .ZN(_12441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21378_ (.A1(_12438_),
    .A2(_12161_),
    .A3(_12441_),
    .ZN(_12442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21379_ (.A1(_12381_),
    .A2(_12273_),
    .ZN(_12443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21380_ (.A1(_15760_),
    .A2(_12173_),
    .B(_12261_),
    .ZN(_12444_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21381_ (.I(_12160_),
    .Z(_12445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21382_ (.A1(_12443_),
    .A2(_12444_),
    .B(_12445_),
    .ZN(_12446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21383_ (.A1(net17),
    .A2(_15762_),
    .B(_12141_),
    .ZN(_12447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21384_ (.A1(_12447_),
    .A2(_12175_),
    .ZN(_12448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21385_ (.A1(_12448_),
    .A2(_12309_),
    .A3(_12387_),
    .ZN(_12449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21386_ (.A1(_12446_),
    .A2(_12449_),
    .B(_12197_),
    .ZN(_12450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21387_ (.A1(_12442_),
    .A2(_12450_),
    .ZN(_12451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21388_ (.A1(_12391_),
    .A2(_12365_),
    .ZN(_12452_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21389_ (.A1(_12452_),
    .A2(_12261_),
    .Z(_12453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21390_ (.A1(_12137_),
    .A2(_12163_),
    .Z(_12454_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21391_ (.A1(_12302_),
    .A2(_15762_),
    .A3(_12454_),
    .Z(_12455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21392_ (.A1(_12453_),
    .A2(_12349_),
    .A3(_12455_),
    .ZN(_12456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21393_ (.A1(_12267_),
    .A2(_12274_),
    .ZN(_12457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21394_ (.I(_12237_),
    .ZN(_12458_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21395_ (.A1(_12458_),
    .A2(_12173_),
    .B(_12213_),
    .ZN(_12459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21396_ (.A1(_12457_),
    .A2(_12459_),
    .B(_12445_),
    .ZN(_12460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21397_ (.A1(_12456_),
    .A2(_12460_),
    .ZN(_12461_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21398_ (.A1(_15767_),
    .A2(_12173_),
    .B(_12168_),
    .ZN(_12462_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21399_ (.A1(_12418_),
    .A2(_12462_),
    .B(_12184_),
    .ZN(_12463_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21400_ (.A1(_12302_),
    .A2(_15758_),
    .Z(_12464_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21401_ (.A1(_12428_),
    .A2(_12244_),
    .A3(_12464_),
    .ZN(_12465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21402_ (.A1(_12463_),
    .A2(_12465_),
    .ZN(_12466_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21403_ (.A1(_12461_),
    .A2(_12466_),
    .A3(_12248_),
    .ZN(_12467_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21404_ (.A1(_12451_),
    .A2(_12467_),
    .A3(_12314_),
    .ZN(_12468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21405_ (.A1(_12435_),
    .A2(_12468_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21406_ (.A1(_12208_),
    .A2(_12219_),
    .Z(_12469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21407_ (.A1(_12447_),
    .A2(_12469_),
    .ZN(_12470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21408_ (.A1(_12365_),
    .A2(_15755_),
    .ZN(_12471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21409_ (.A1(_12471_),
    .A2(_12368_),
    .ZN(_12472_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _21410_ (.A1(_12470_),
    .A2(_12472_),
    .A3(_12122_),
    .Z(_12473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21411_ (.A1(_12228_),
    .A2(_12238_),
    .ZN(_12474_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21412_ (.A1(_12474_),
    .A2(_12209_),
    .A3(_12222_),
    .Z(_12475_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21413_ (.A1(_12473_),
    .A2(_12475_),
    .B(_12185_),
    .ZN(_12476_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21414_ (.A1(_12203_),
    .A2(_12168_),
    .A3(_12208_),
    .Z(_12477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21415_ (.A1(_12096_),
    .A2(_15755_),
    .ZN(_12478_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21416_ (.A1(_12477_),
    .A2(_12478_),
    .B(_12326_),
    .ZN(_12479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21417_ (.A1(_12295_),
    .A2(_12141_),
    .Z(_12480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21418_ (.A1(_12480_),
    .A2(_12177_),
    .ZN(_12481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21419_ (.A1(_12357_),
    .A2(_12481_),
    .ZN(_12482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21420_ (.A1(_12479_),
    .A2(_12482_),
    .B(_12197_),
    .ZN(_12483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21421_ (.A1(_12476_),
    .A2(_12483_),
    .ZN(_12484_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21422_ (.A1(_12234_),
    .A2(_12213_),
    .Z(_12485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21423_ (.A1(_12316_),
    .A2(_12320_),
    .A3(_12175_),
    .ZN(_12486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21424_ (.A1(_12485_),
    .A2(_12486_),
    .B(_12184_),
    .ZN(_12487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21425_ (.A1(_12202_),
    .A2(_12205_),
    .ZN(_12488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21426_ (.A1(_12267_),
    .A2(_12316_),
    .ZN(_12489_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21427_ (.A1(_12488_),
    .A2(_12489_),
    .A3(_12244_),
    .ZN(_12490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21428_ (.A1(_12487_),
    .A2(_12490_),
    .B(_12198_),
    .ZN(_12491_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21429_ (.A1(_12469_),
    .A2(_12388_),
    .Z(_12492_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21430_ (.I(_12478_),
    .ZN(_12493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21431_ (.A1(_12493_),
    .A2(_12216_),
    .B(_12168_),
    .ZN(_12494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21432_ (.I(_12233_),
    .ZN(_12495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21433_ (.A1(_12495_),
    .A2(_12206_),
    .Z(_12496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21434_ (.I(_12496_),
    .ZN(_12497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21435_ (.A1(_12492_),
    .A2(_12494_),
    .A3(_12497_),
    .ZN(_12498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21436_ (.A1(_12316_),
    .A2(_12320_),
    .A3(_12177_),
    .ZN(_12499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21437_ (.A1(_12055_),
    .A2(_12274_),
    .A3(_12242_),
    .ZN(_12500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21438_ (.A1(_12499_),
    .A2(_12244_),
    .A3(_12500_),
    .ZN(_12501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21439_ (.A1(_12498_),
    .A2(_12185_),
    .A3(_12501_),
    .ZN(_12502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21440_ (.A1(_12491_),
    .A2(_12502_),
    .ZN(_12503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21441_ (.A1(_12484_),
    .A2(_12314_),
    .A3(_12503_),
    .ZN(_12504_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21442_ (.I(_12264_),
    .ZN(_12505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21443_ (.A1(_12180_),
    .A2(_12505_),
    .B(_12160_),
    .ZN(_12506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21444_ (.A1(_12506_),
    .A2(_12411_),
    .B(_12310_),
    .ZN(_12507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21445_ (.A1(_12170_),
    .A2(net13),
    .ZN(_12508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21446_ (.A1(_15755_),
    .A2(_12454_),
    .ZN(_12509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21447_ (.A1(_12509_),
    .A2(_12206_),
    .ZN(_12510_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21448_ (.I(_12354_),
    .ZN(_12511_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21449_ (.A1(_12510_),
    .A2(_12511_),
    .Z(_12512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21450_ (.A1(_12508_),
    .A2(_12512_),
    .A3(_12246_),
    .ZN(_12513_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21451_ (.A1(_12507_),
    .A2(_12513_),
    .B(_12198_),
    .ZN(_12514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21452_ (.A1(_12133_),
    .A2(_12238_),
    .B(_12097_),
    .ZN(_12515_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21453_ (.A1(_12515_),
    .A2(_12496_),
    .B(_12445_),
    .ZN(_12516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21454_ (.I(_12232_),
    .ZN(_12517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21455_ (.A1(_12517_),
    .A2(_12184_),
    .B1(_12180_),
    .B2(net1149),
    .ZN(_12518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21456_ (.A1(_12516_),
    .A2(_12518_),
    .ZN(_12519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21457_ (.A1(_12519_),
    .A2(_12214_),
    .ZN(_12520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21458_ (.A1(_12520_),
    .A2(_12514_),
    .B(_12314_),
    .ZN(_12521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21459_ (.A1(_12296_),
    .A2(_12509_),
    .ZN(_12522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21460_ (.A1(_12349_),
    .A2(_12522_),
    .B(_12310_),
    .ZN(_12523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21461_ (.A1(_12409_),
    .A2(_12310_),
    .ZN(_12524_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21462_ (.I(_12524_),
    .ZN(_12525_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21463_ (.A1(_12523_),
    .A2(_12525_),
    .B(_12161_),
    .ZN(_12526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _21464_ (.A1(_12124_),
    .A2(_12505_),
    .B(_12388_),
    .ZN(_12527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21465_ (.A1(_12179_),
    .A2(_12130_),
    .ZN(_12528_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21466_ (.A1(_12527_),
    .A2(_12387_),
    .A3(_12528_),
    .ZN(_12529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21467_ (.A1(_12272_),
    .A2(_12393_),
    .ZN(_12530_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21468_ (.A1(_12529_),
    .A2(_12530_),
    .A3(_12326_),
    .ZN(_12531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21469_ (.A1(_12526_),
    .A2(_12531_),
    .A3(_12199_),
    .ZN(_12532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21470_ (.A1(_12521_),
    .A2(_12532_),
    .ZN(_12533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21471_ (.A1(_12504_),
    .A2(_12533_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21472_ (.A1(_12332_),
    .A2(_12141_),
    .Z(_12534_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21473_ (.A1(_12534_),
    .A2(_12121_),
    .ZN(_12535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21474_ (.A1(_12225_),
    .A2(_12097_),
    .ZN(_12536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21475_ (.A1(_12535_),
    .A2(_12536_),
    .B(_12160_),
    .ZN(_12537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21476_ (.A1(_12385_),
    .A2(net1164),
    .B(_12213_),
    .ZN(_12538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21477_ (.A1(_12538_),
    .A2(_12146_),
    .ZN(_12539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21478_ (.A1(_12537_),
    .A2(_12539_),
    .ZN(_12540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21479_ (.A1(_12202_),
    .A2(_12354_),
    .ZN(_12541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21480_ (.A1(_12391_),
    .A2(_12213_),
    .ZN(_12542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21481_ (.A1(_12541_),
    .A2(_12542_),
    .B(_12184_),
    .ZN(_12543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21482_ (.A1(_12458_),
    .A2(_12129_),
    .B(_12121_),
    .ZN(_12544_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21483_ (.A1(_12317_),
    .A2(_12544_),
    .A3(_12142_),
    .ZN(_12545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21484_ (.A1(_12543_),
    .A2(_12545_),
    .ZN(_12546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21485_ (.A1(_12540_),
    .A2(_12546_),
    .ZN(_12547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21486_ (.A1(_12547_),
    .A2(_12199_),
    .ZN(_12548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21487_ (.A1(_12133_),
    .A2(_12201_),
    .B(_12097_),
    .ZN(_12549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21488_ (.A1(_12296_),
    .A2(_12133_),
    .ZN(_12550_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21489_ (.I(_12550_),
    .ZN(_12551_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21490_ (.A1(_12549_),
    .A2(_12551_),
    .B(_12310_),
    .ZN(_12552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21491_ (.A1(_15751_),
    .A2(_12281_),
    .B(_12213_),
    .ZN(_12553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21492_ (.A1(_12206_),
    .A2(_12280_),
    .ZN(_12554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21493_ (.A1(_12553_),
    .A2(_12554_),
    .B(_12160_),
    .ZN(_12555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21494_ (.A1(_12552_),
    .A2(_12555_),
    .B(_12198_),
    .ZN(_12556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21495_ (.A1(_12293_),
    .A2(_12209_),
    .A3(_12303_),
    .ZN(_12557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21496_ (.A1(_12205_),
    .A2(_12316_),
    .A3(_12302_),
    .ZN(_12558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21497_ (.A1(_12296_),
    .A2(_12201_),
    .ZN(_12559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21498_ (.A1(_12558_),
    .A2(_12559_),
    .A3(_12261_),
    .ZN(_12560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21499_ (.A1(_12557_),
    .A2(_12560_),
    .ZN(_12561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21500_ (.A1(_12561_),
    .A2(_12246_),
    .ZN(_12562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21501_ (.A1(_12556_),
    .A2(_12562_),
    .ZN(_12563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21502_ (.A1(_12548_),
    .A2(_12563_),
    .ZN(_12564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21503_ (.A1(_12564_),
    .A2(_12257_),
    .ZN(_12565_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21504_ (.A1(_12377_),
    .A2(_12458_),
    .B(_12181_),
    .ZN(_12566_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21505_ (.A1(_12422_),
    .A2(_12281_),
    .A3(_12133_),
    .Z(_12567_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21506_ (.A1(_12566_),
    .A2(_12567_),
    .ZN(_12568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21507_ (.A1(_12447_),
    .A2(_12273_),
    .ZN(_12569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21508_ (.A1(_12569_),
    .A2(_12419_),
    .B(_12122_),
    .ZN(_12570_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21509_ (.A1(_12568_),
    .A2(_12570_),
    .B(_12161_),
    .ZN(_12571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21510_ (.A1(_12554_),
    .A2(_12264_),
    .Z(_12572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21511_ (.A1(_12379_),
    .A2(_12572_),
    .B(_12445_),
    .ZN(_12573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21512_ (.A1(_12331_),
    .A2(_12233_),
    .ZN(_12574_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21513_ (.A1(_12574_),
    .A2(_12297_),
    .A3(_12244_),
    .ZN(_12575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21514_ (.A1(_12573_),
    .A2(_12575_),
    .B(_12198_),
    .ZN(_12576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21515_ (.A1(_12576_),
    .A2(_12571_),
    .ZN(_12577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21516_ (.A1(_12439_),
    .A2(_12339_),
    .A3(_12169_),
    .ZN(_12578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21517_ (.A1(_12365_),
    .A2(_12134_),
    .A3(_12320_),
    .ZN(_12579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21518_ (.A1(_12134_),
    .A2(_12242_),
    .A3(_12241_),
    .ZN(_12580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21519_ (.A1(_12579_),
    .A2(_12580_),
    .A3(_12387_),
    .ZN(_12581_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21520_ (.A1(_12578_),
    .A2(_12581_),
    .A3(_12161_),
    .ZN(_12582_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21521_ (.A1(_12338_),
    .A2(_12097_),
    .A3(_12175_),
    .ZN(_12583_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21522_ (.A1(_12583_),
    .A2(_12244_),
    .A3(_12344_),
    .ZN(_12584_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21523_ (.I(_12296_),
    .ZN(_12585_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21524_ (.A1(_12138_),
    .A2(_12181_),
    .ZN(_12586_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21525_ (.A1(_12585_),
    .A2(_12586_),
    .B(_12445_),
    .ZN(_12587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21526_ (.A1(_12584_),
    .A2(_12587_),
    .B(_12197_),
    .ZN(_12588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21527_ (.A1(_12582_),
    .A2(_12588_),
    .ZN(_12589_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21528_ (.A1(_12589_),
    .A2(_12314_),
    .A3(_12577_),
    .ZN(_12590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21529_ (.A1(_12565_),
    .A2(_12590_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21530_ (.A1(_12471_),
    .A2(_12388_),
    .A3(_12238_),
    .ZN(_12591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21531_ (.A1(_12170_),
    .A2(_12365_),
    .ZN(_12592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21532_ (.A1(_12591_),
    .A2(_12592_),
    .ZN(_12593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21533_ (.A1(_12593_),
    .A2(_12326_),
    .ZN(_12594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21534_ (.A1(_12554_),
    .A2(_12160_),
    .Z(_12595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21535_ (.A1(_12534_),
    .A2(_12308_),
    .ZN(_12596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21536_ (.A1(_12595_),
    .A2(_12596_),
    .B(_12244_),
    .ZN(_12597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21537_ (.A1(_12594_),
    .A2(_12597_),
    .ZN(_12598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21538_ (.A1(_12178_),
    .A2(_12281_),
    .ZN(_12599_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21539_ (.A1(_12266_),
    .A2(_12301_),
    .B(_12160_),
    .C(_12599_),
    .ZN(_12600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21540_ (.A1(net17),
    .A2(_12388_),
    .B(_12160_),
    .ZN(_12601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21541_ (.A1(_12601_),
    .A2(_12558_),
    .ZN(_12602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21542_ (.A1(_12600_),
    .A2(_12602_),
    .ZN(_12603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21543_ (.A1(_12603_),
    .A2(_12169_),
    .ZN(_12604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21544_ (.A1(_12598_),
    .A2(_12248_),
    .A3(_12604_),
    .ZN(_12605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21545_ (.A1(_12356_),
    .A2(_12164_),
    .ZN(_12606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21546_ (.A1(_12144_),
    .A2(_12606_),
    .ZN(_12607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21547_ (.A1(net1155),
    .A2(_12480_),
    .ZN(_12608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21548_ (.A1(net1160),
    .A2(_12180_),
    .B(_12181_),
    .ZN(_12609_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21549_ (.A1(_12608_),
    .A2(_12609_),
    .A3(_12287_),
    .ZN(_12610_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21550_ (.A1(_12607_),
    .A2(_12610_),
    .A3(_12185_),
    .ZN(_12611_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21551_ (.A1(_12228_),
    .A2(_12222_),
    .ZN(_12612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21552_ (.A1(_12612_),
    .A2(_12527_),
    .ZN(_12613_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21553_ (.A1(_12385_),
    .A2(_12181_),
    .ZN(_12614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21554_ (.A1(_12391_),
    .A2(_12205_),
    .ZN(_12615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21555_ (.A1(_12614_),
    .A2(_12615_),
    .ZN(_12616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21556_ (.A1(_12613_),
    .A2(_12616_),
    .A3(_12246_),
    .ZN(_12617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21557_ (.A1(_12611_),
    .A2(_12199_),
    .A3(_12617_),
    .ZN(_12618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21558_ (.A1(_12605_),
    .A2(_12618_),
    .A3(_12314_),
    .ZN(_12619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21559_ (.A1(_12145_),
    .A2(_12320_),
    .ZN(_12620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21560_ (.A1(_12306_),
    .A2(_12180_),
    .ZN(_12621_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21561_ (.A1(_12620_),
    .A2(_12511_),
    .B(_12387_),
    .C(_12621_),
    .ZN(_12622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21562_ (.A1(_12305_),
    .A2(_12281_),
    .ZN(_12623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21563_ (.A1(_12146_),
    .A2(_12262_),
    .A3(_12623_),
    .ZN(_12624_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21564_ (.A1(_12622_),
    .A2(_12624_),
    .A3(_12161_),
    .ZN(_12625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21565_ (.A1(net1150),
    .A2(_12242_),
    .B(_12261_),
    .ZN(_12626_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21566_ (.A1(_12204_),
    .A2(_12626_),
    .B(_12445_),
    .ZN(_12627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21567_ (.A1(_12125_),
    .A2(_12267_),
    .ZN(_12628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21568_ (.A1(_12480_),
    .A2(_12134_),
    .ZN(_12629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21569_ (.A1(_12628_),
    .A2(_12387_),
    .A3(_12629_),
    .ZN(_12630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21570_ (.A1(_12627_),
    .A2(_12630_),
    .B(_12197_),
    .ZN(_12631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21571_ (.A1(_12625_),
    .A2(_12631_),
    .ZN(_12632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21572_ (.I(_12177_),
    .ZN(_12633_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21573_ (.A1(_12633_),
    .A2(_12511_),
    .A3(_12097_),
    .Z(_12634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21574_ (.A1(_12267_),
    .A2(_12289_),
    .ZN(_12635_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21575_ (.A1(_12634_),
    .A2(_12214_),
    .A3(_12635_),
    .ZN(_12636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21576_ (.A1(_12218_),
    .A2(_12242_),
    .B(_12261_),
    .ZN(_12637_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21577_ (.A1(_12620_),
    .A2(_12637_),
    .B(_12184_),
    .ZN(_12638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21578_ (.A1(_12636_),
    .A2(_12638_),
    .ZN(_12639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21579_ (.I(_12145_),
    .ZN(_12640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21580_ (.A1(_12510_),
    .A2(_12168_),
    .Z(_12641_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21581_ (.A1(_12428_),
    .A2(_12640_),
    .B(_12641_),
    .ZN(_12642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21582_ (.A1(_12379_),
    .A2(_12355_),
    .B(_12445_),
    .ZN(_12643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21583_ (.A1(_12642_),
    .A2(_12643_),
    .ZN(_12644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21584_ (.A1(_12639_),
    .A2(_12644_),
    .A3(_12248_),
    .ZN(_12645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21585_ (.A1(_12632_),
    .A2(_12645_),
    .A3(_12257_),
    .ZN(_12646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21586_ (.A1(_12619_),
    .A2(_12646_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21587_ (.A1(_12125_),
    .A2(_12130_),
    .A3(net13),
    .ZN(_12647_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21588_ (.A1(_12647_),
    .A2(_12214_),
    .A3(_12464_),
    .ZN(_12648_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21589_ (.A1(_12125_),
    .A2(_12221_),
    .A3(_12134_),
    .ZN(_12649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21590_ (.A1(_12534_),
    .A2(_12177_),
    .ZN(_12650_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21591_ (.A1(_12649_),
    .A2(_12169_),
    .A3(_12650_),
    .ZN(_12651_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21592_ (.A1(_12648_),
    .A2(_12651_),
    .A3(_12185_),
    .ZN(_12652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21593_ (.A1(_12306_),
    .A2(_12130_),
    .B(_12181_),
    .ZN(_12653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21594_ (.A1(_12201_),
    .A2(net20),
    .ZN(_12654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21595_ (.A1(_12654_),
    .A2(_12221_),
    .ZN(_12655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21596_ (.A1(_12653_),
    .A2(_12655_),
    .B(_12326_),
    .ZN(_12656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21597_ (.A1(_12368_),
    .A2(_12509_),
    .B(_12222_),
    .ZN(_12657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21598_ (.A1(_12273_),
    .A2(_12221_),
    .A3(_12208_),
    .ZN(_12658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21599_ (.A1(_12657_),
    .A2(_12658_),
    .ZN(_12659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21600_ (.A1(_12656_),
    .A2(_12659_),
    .B(_12199_),
    .ZN(_12660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21601_ (.A1(_12652_),
    .A2(_12660_),
    .ZN(_12661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21602_ (.A1(_15762_),
    .A2(_15741_),
    .ZN(_12662_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _21603_ (.A1(_12388_),
    .A2(_12259_),
    .A3(_12662_),
    .A4(_12264_),
    .ZN(_12663_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21604_ (.A1(_12663_),
    .A2(_12282_),
    .A3(_12623_),
    .ZN(_12664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21605_ (.A1(_12055_),
    .A2(_12295_),
    .A3(_12129_),
    .ZN(_12665_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21606_ (.A1(_12452_),
    .A2(_12665_),
    .A3(_12287_),
    .ZN(_12666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21607_ (.A1(_12666_),
    .A2(_12122_),
    .ZN(_12667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21608_ (.A1(_12664_),
    .A2(_12667_),
    .ZN(_12668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21609_ (.A1(_12668_),
    .A2(_12161_),
    .ZN(_12669_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21610_ (.A1(_12276_),
    .A2(_12505_),
    .B(_12242_),
    .ZN(_12670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21611_ (.A1(_12544_),
    .A2(_12670_),
    .B(_12445_),
    .ZN(_12671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21612_ (.A1(_12447_),
    .A2(_12205_),
    .ZN(_12672_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21613_ (.A1(_15756_),
    .A2(_15765_),
    .B(_12173_),
    .ZN(_12673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21614_ (.A1(_12672_),
    .A2(_12244_),
    .A3(_12673_),
    .ZN(_12674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21615_ (.A1(_12671_),
    .A2(_12674_),
    .B(_12197_),
    .ZN(_12675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21616_ (.A1(_12669_),
    .A2(_12675_),
    .ZN(_12676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21617_ (.A1(_12661_),
    .A2(_12676_),
    .A3(_12314_),
    .ZN(_12677_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21618_ (.A1(_15755_),
    .A2(_15753_),
    .Z(_12678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21619_ (.A1(_12124_),
    .A2(_12678_),
    .B(_12320_),
    .ZN(_12679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21620_ (.A1(_12203_),
    .A2(_12180_),
    .A3(_12208_),
    .ZN(_12680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21621_ (.A1(_12679_),
    .A2(_12680_),
    .A3(_12387_),
    .ZN(_12681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21622_ (.A1(net17),
    .A2(_12302_),
    .ZN(_12682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21623_ (.A1(_12477_),
    .A2(_12682_),
    .ZN(_12683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21624_ (.A1(_12681_),
    .A2(_12683_),
    .A3(_12185_),
    .ZN(_12684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21625_ (.A1(_12633_),
    .A2(_12173_),
    .B(_12222_),
    .ZN(_12685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21626_ (.A1(_12527_),
    .A2(_12685_),
    .B(_12184_),
    .ZN(_12686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21627_ (.A1(_12377_),
    .A2(_12261_),
    .Z(_12687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21628_ (.A1(_12176_),
    .A2(_12687_),
    .ZN(_12688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21629_ (.A1(_12686_),
    .A2(_12688_),
    .ZN(_12689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21630_ (.A1(_12684_),
    .A2(_12199_),
    .A3(_12689_),
    .ZN(_12690_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21631_ (.A1(_12551_),
    .A2(_12290_),
    .B(_12222_),
    .ZN(_12691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21632_ (.A1(_12423_),
    .A2(_12122_),
    .ZN(_12692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21633_ (.A1(_12691_),
    .A2(_12692_),
    .ZN(_12693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21634_ (.A1(_12693_),
    .A2(_12161_),
    .ZN(_12694_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21635_ (.A1(_12633_),
    .A2(_12355_),
    .B(_12324_),
    .C(_12310_),
    .ZN(_12695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21636_ (.I(_15757_),
    .ZN(_12696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21637_ (.A1(_12696_),
    .A2(_12242_),
    .B(_12261_),
    .ZN(_12697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21638_ (.A1(_12697_),
    .A2(_12629_),
    .B(_12445_),
    .ZN(_12698_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21639_ (.A1(_12695_),
    .A2(_12698_),
    .B(_12198_),
    .ZN(_12699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21640_ (.A1(_12694_),
    .A2(_12699_),
    .ZN(_12700_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21641_ (.A1(_12690_),
    .A2(_12700_),
    .A3(_12257_),
    .ZN(_12701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21642_ (.A1(_12677_),
    .A2(_12701_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21643_ (.A1(_12121_),
    .A2(_12237_),
    .Z(_12702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21644_ (.A1(_12702_),
    .A2(_12277_),
    .Z(_12703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21645_ (.A1(_12391_),
    .A2(net17),
    .ZN(_12704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21646_ (.A1(_12703_),
    .A2(_12704_),
    .B(_12326_),
    .ZN(_12705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21647_ (.A1(_12130_),
    .A2(net1160),
    .ZN(_12706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21648_ (.A1(_12672_),
    .A2(_12706_),
    .A3(_12214_),
    .ZN(_12707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21649_ (.A1(_12705_),
    .A2(_12707_),
    .B(_12248_),
    .ZN(_12708_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21650_ (.A1(_12141_),
    .A2(net71),
    .Z(_12709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21651_ (.A1(_12709_),
    .A2(_15762_),
    .Z(_12710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21652_ (.A1(_12682_),
    .A2(_12261_),
    .ZN(_12711_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21653_ (.A1(_12710_),
    .A2(_12711_),
    .ZN(_12712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21654_ (.A1(_12712_),
    .A2(_12522_),
    .B(_12246_),
    .ZN(_12713_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21655_ (.A1(_12710_),
    .A2(_12143_),
    .ZN(_12714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21656_ (.A1(_12289_),
    .A2(_12177_),
    .A3(_12221_),
    .ZN(_12715_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21657_ (.A1(_12714_),
    .A2(_12459_),
    .A3(_12715_),
    .ZN(_12716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21658_ (.A1(_12713_),
    .A2(_12716_),
    .ZN(_12717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21659_ (.A1(_12708_),
    .A2(_12717_),
    .ZN(_12718_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21660_ (.A1(_12505_),
    .A2(_12302_),
    .Z(_12719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21661_ (.A1(_12206_),
    .A2(_15765_),
    .ZN(_12720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21662_ (.A1(_12720_),
    .A2(_12168_),
    .ZN(_12721_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21663_ (.A1(_12719_),
    .A2(_12721_),
    .ZN(_12722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21664_ (.A1(_12495_),
    .A2(_12130_),
    .ZN(_12723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21665_ (.A1(_12722_),
    .A2(_12723_),
    .B(_12326_),
    .ZN(_12724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21666_ (.A1(_12170_),
    .A2(_12134_),
    .ZN(_12725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21667_ (.A1(_12381_),
    .A2(_12177_),
    .ZN(_12726_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21668_ (.A1(_12725_),
    .A2(_12726_),
    .A3(_12214_),
    .ZN(_12727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21669_ (.A1(_12724_),
    .A2(_12727_),
    .ZN(_12728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21670_ (.I(_15751_),
    .ZN(_12729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21671_ (.A1(_12729_),
    .A2(_12180_),
    .B(_12222_),
    .ZN(_12730_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21672_ (.A1(_12730_),
    .A2(_12277_),
    .B(_12445_),
    .ZN(_12731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21673_ (.A1(_12654_),
    .A2(_12320_),
    .ZN(_12732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21674_ (.A1(_12317_),
    .A2(_12387_),
    .A3(_12732_),
    .ZN(_12733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21675_ (.A1(_12731_),
    .A2(_12733_),
    .ZN(_12734_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21676_ (.A1(_12728_),
    .A2(_12248_),
    .A3(_12734_),
    .ZN(_12735_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21677_ (.A1(_12735_),
    .A2(_12314_),
    .A3(_12718_),
    .ZN(_12736_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21678_ (.A1(_12331_),
    .A2(_12222_),
    .ZN(_12737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21679_ (.A1(_12737_),
    .A2(_12550_),
    .B(_12197_),
    .ZN(_12738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21680_ (.A1(_12170_),
    .A2(net1155),
    .ZN(_12739_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21681_ (.A1(_12494_),
    .A2(_12739_),
    .A3(_12452_),
    .ZN(_12740_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21682_ (.A1(_12738_),
    .A2(_12740_),
    .B(_12246_),
    .ZN(_12741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21683_ (.A1(net1158),
    .A2(_12130_),
    .A3(_12134_),
    .ZN(_12742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21684_ (.A1(_12742_),
    .A2(_12169_),
    .A3(_12439_),
    .ZN(_12743_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21685_ (.I(_12709_),
    .ZN(_12744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21686_ (.A1(_12583_),
    .A2(_12744_),
    .ZN(_12745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21687_ (.A1(_12745_),
    .A2(_12214_),
    .ZN(_12746_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21688_ (.A1(_12743_),
    .A2(_12746_),
    .A3(_12248_),
    .ZN(_12747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21689_ (.A1(_12741_),
    .A2(_12747_),
    .ZN(_12748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21690_ (.A1(_12232_),
    .A2(_12168_),
    .Z(_12749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21691_ (.A1(_12493_),
    .A2(_12365_),
    .ZN(_12750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21692_ (.A1(_12749_),
    .A2(_12750_),
    .B(_12198_),
    .ZN(_12751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21693_ (.A1(net1155),
    .A2(_12180_),
    .B(_12181_),
    .ZN(_12752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21694_ (.A1(_12225_),
    .A2(_12130_),
    .A3(_12177_),
    .ZN(_12753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21695_ (.A1(_12752_),
    .A2(_12753_),
    .ZN(_12754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21696_ (.A1(_12751_),
    .A2(_12754_),
    .B(_12326_),
    .ZN(_12755_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21697_ (.A1(_12508_),
    .A2(_12387_),
    .A3(_12382_),
    .ZN(_12756_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21698_ (.A1(_12448_),
    .A2(_12244_),
    .A3(_12665_),
    .ZN(_12757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21699_ (.A1(_12199_),
    .A2(_12757_),
    .A3(_12756_),
    .ZN(_12758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21700_ (.A1(_12758_),
    .A2(_12755_),
    .ZN(_12759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21701_ (.A1(_12759_),
    .A2(_12748_),
    .A3(_12257_),
    .ZN(_12760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21702_ (.A1(_12760_),
    .A2(_12736_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21703_ (.I(\sa03_sr[7] ),
    .ZN(_12761_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21704_ (.I(net726),
    .ZN(_12762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21705_ (.A1(_12761_),
    .A2(_12762_),
    .ZN(_12763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21706_ (.A1(\sa03_sr[7] ),
    .A2(net720),
    .ZN(_12764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21707_ (.A1(_12763_),
    .A2(_12764_),
    .ZN(_12765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _21708_ (.I(\sa32_sub[1] ),
    .ZN(_12766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21709_ (.A1(net777),
    .A2(_12766_),
    .ZN(_12767_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21710_ (.I(\sa21_sub[1] ),
    .ZN(_12768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21711_ (.A1(_12768_),
    .A2(\sa32_sub[1] ),
    .ZN(_12769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21712_ (.A1(_12769_),
    .A2(_12767_),
    .ZN(_12770_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21713_ (.A1(_12770_),
    .A2(_12765_),
    .ZN(_12771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21714_ (.A1(_12762_),
    .A2(\sa03_sr[7] ),
    .ZN(_12772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21715_ (.A1(_12761_),
    .A2(net721),
    .ZN(_12773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21716_ (.A1(_12772_),
    .A2(_12773_),
    .ZN(_12774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21717_ (.A1(_12768_),
    .A2(_12766_),
    .ZN(_12775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21718_ (.A1(\sa21_sub[1] ),
    .A2(\sa32_sub[1] ),
    .ZN(_12776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21719_ (.A1(_12776_),
    .A2(_12775_),
    .ZN(_12777_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21720_ (.A1(_12774_),
    .A2(_12777_),
    .ZN(_12778_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21721_ (.A1(_12778_),
    .A2(_12771_),
    .ZN(_12779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21722_ (.I(\sa10_sub[0] ),
    .ZN(_12780_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21723_ (.I(\sa10_sub[7] ),
    .Z(_12781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21724_ (.A1(_12781_),
    .A2(_12780_),
    .ZN(_12782_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21725_ (.I(\sa10_sub[7] ),
    .ZN(_12783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21726_ (.A1(_12783_),
    .A2(net722),
    .ZN(_12784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21727_ (.A1(_12784_),
    .A2(_12782_),
    .ZN(_12785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21728_ (.A1(net736),
    .A2(_12785_),
    .ZN(_12786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21729_ (.A1(_12783_),
    .A2(_12780_),
    .ZN(_12787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21730_ (.A1(_12781_),
    .A2(net722),
    .ZN(_12788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21731_ (.A1(_12787_),
    .A2(_12788_),
    .ZN(_12789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21732_ (.I(\sa10_sub[1] ),
    .ZN(_12790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21733_ (.A1(_12789_),
    .A2(_12790_),
    .ZN(_12791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21734_ (.A1(_12791_),
    .A2(_12786_),
    .ZN(_12792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21735_ (.A1(_12779_),
    .A2(_12792_),
    .ZN(_12793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21736_ (.A1(_12774_),
    .A2(_12777_),
    .ZN(_12794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21737_ (.A1(_12765_),
    .A2(_12770_),
    .ZN(_12795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21738_ (.A1(_12794_),
    .A2(_12795_),
    .ZN(_12796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21739_ (.A1(_12789_),
    .A2(net736),
    .ZN(_12797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21740_ (.A1(_12785_),
    .A2(_12790_),
    .ZN(_12798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21741_ (.A1(_12797_),
    .A2(_12798_),
    .ZN(_12799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21742_ (.A1(_12796_),
    .A2(_12799_),
    .ZN(_12800_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21743_ (.A1(_12793_),
    .A2(_12800_),
    .A3(_10402_),
    .ZN(_12801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21744_ (.A1(_10410_),
    .A2(\text_in_r[25] ),
    .ZN(_12802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21745_ (.A1(_12801_),
    .A2(_12802_),
    .ZN(_12803_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21746_ (.I(net626),
    .ZN(_12804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21747_ (.A1(_12804_),
    .A2(_12803_),
    .ZN(_12805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21748_ (.A1(net771),
    .A2(net627),
    .A3(_12802_),
    .ZN(_12806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21749_ (.A1(_12805_),
    .A2(_12806_),
    .ZN(_15775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21750_ (.A1(_12783_),
    .A2(_12761_),
    .ZN(_12807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21751_ (.A1(\sa03_sr[7] ),
    .A2(\sa10_sub[7] ),
    .ZN(_12808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21752_ (.A1(_12808_),
    .A2(_12807_),
    .ZN(_12809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21753_ (.A1(net746),
    .A2(_12809_),
    .ZN(_12810_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21754_ (.I(\sa32_sub[0] ),
    .ZN(_12811_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21755_ (.A1(net971),
    .A2(_12811_),
    .A3(_12808_),
    .ZN(_12812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21756_ (.A1(_12812_),
    .A2(_12810_),
    .ZN(_12813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21757_ (.A1(net532),
    .A2(_12780_),
    .ZN(_12814_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21758_ (.I(\sa21_sub[0] ),
    .ZN(_12815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21759_ (.A1(_12815_),
    .A2(\sa10_sub[0] ),
    .ZN(_12816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21760_ (.A1(_12816_),
    .A2(_12814_),
    .ZN(_12817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21761_ (.A1(_12817_),
    .A2(_12813_),
    .ZN(_12818_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21762_ (.I(_12817_),
    .ZN(_12819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21763_ (.A1(net974),
    .A2(_12812_),
    .A3(_12819_),
    .ZN(_12820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21764_ (.A1(_12818_),
    .A2(_12820_),
    .B(_10410_),
    .ZN(_12821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21765_ (.I(\text_in_r[24] ),
    .ZN(_12822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21766_ (.A1(_12822_),
    .A2(_10431_),
    .Z(_12823_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21767_ (.A1(_12821_),
    .A2(_12823_),
    .B(\u0.tmp_w[24] ),
    .ZN(_12824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21768_ (.A1(_12818_),
    .A2(_12820_),
    .ZN(_12825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21769_ (.A1(_12825_),
    .A2(_11989_),
    .ZN(_12826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21770_ (.I(\u0.tmp_w[24] ),
    .ZN(_12827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21771_ (.I(_12823_),
    .ZN(_12828_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21772_ (.A1(net964),
    .A2(_12827_),
    .A3(_12828_),
    .ZN(_12829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21773_ (.A1(_12829_),
    .A2(_12824_),
    .ZN(_15778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21774_ (.I(\sa03_sr[1] ),
    .ZN(_12830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21775_ (.A1(_12790_),
    .A2(_12830_),
    .ZN(_12831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21776_ (.A1(net734),
    .A2(\sa03_sr[1] ),
    .ZN(_12832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21777_ (.A1(_12831_),
    .A2(_12832_),
    .ZN(_12833_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21778_ (.I(\sa21_sub[2] ),
    .ZN(_12834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21779_ (.A1(_12833_),
    .A2(_12834_),
    .ZN(_12835_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _21780_ (.I(\sa21_sub[2] ),
    .Z(_12836_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21781_ (.A1(_12831_),
    .A2(_12836_),
    .A3(_12832_),
    .ZN(_12837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21782_ (.A1(_12835_),
    .A2(_12837_),
    .ZN(_12838_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21783_ (.I(\sa32_sub[2] ),
    .ZN(_12839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21784_ (.A1(_12839_),
    .A2(\sa10_sub[2] ),
    .ZN(_12840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21785_ (.I(\sa10_sub[2] ),
    .ZN(_12841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21786_ (.A1(_12841_),
    .A2(\sa32_sub[2] ),
    .ZN(_12842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21787_ (.A1(_12840_),
    .A2(_12842_),
    .ZN(_12843_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21788_ (.I(_12843_),
    .ZN(_12844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21789_ (.A1(_12838_),
    .A2(_12844_),
    .ZN(_12845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21790_ (.A1(_12835_),
    .A2(_12837_),
    .A3(_12843_),
    .ZN(_12846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21791_ (.A1(_12845_),
    .A2(_12846_),
    .B(_10381_),
    .ZN(_12847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21792_ (.I(\text_in_r[26] ),
    .ZN(_12848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21793_ (.A1(_12848_),
    .A2(net596),
    .Z(_12849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21794_ (.I(\u0.tmp_w[26] ),
    .ZN(_12850_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _21795_ (.A1(_12847_),
    .A2(_12849_),
    .B(_12850_),
    .ZN(_12851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21796_ (.A1(_12845_),
    .A2(_12846_),
    .ZN(_12852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21797_ (.A1(_12852_),
    .A2(_10402_),
    .ZN(_12853_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21798_ (.I(_12849_),
    .ZN(_12854_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21799_ (.A1(_12854_),
    .A2(\u0.tmp_w[26] ),
    .A3(_12853_),
    .ZN(_12855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21800_ (.A1(_12851_),
    .A2(_12855_),
    .ZN(_12856_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _21801_ (.I(_12856_),
    .Z(_15794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _21802_ (.A1(_12823_),
    .A2(_12821_),
    .B(_12827_),
    .ZN(_12857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21803_ (.A1(_12826_),
    .A2(\u0.tmp_w[24] ),
    .A3(_12828_),
    .ZN(_12858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21804_ (.A1(_12857_),
    .A2(_12858_),
    .ZN(_15769_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21805_ (.A1(_12847_),
    .A2(_12849_),
    .B(\u0.tmp_w[26] ),
    .ZN(_12859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21806_ (.A1(_12853_),
    .A2(_12850_),
    .A3(_12854_),
    .ZN(_12860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21807_ (.A1(_12859_),
    .A2(_12860_),
    .ZN(_12861_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21808_ (.I(_12861_),
    .Z(_15787_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _21809_ (.I(_12856_),
    .Z(_12862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21810_ (.A1(net41),
    .A2(_12862_),
    .A3(net12),
    .ZN(_12863_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21811_ (.I(\sa03_sr[2] ),
    .ZN(_12864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21812_ (.A1(_12761_),
    .A2(_12864_),
    .ZN(_12865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21813_ (.A1(net39),
    .A2(\sa03_sr[2] ),
    .ZN(_12866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21814_ (.A1(_12865_),
    .A2(_12866_),
    .ZN(_12867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21815_ (.I(\sa32_sub[3] ),
    .ZN(_12868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21816_ (.A1(_12868_),
    .A2(\sa21_sub[3] ),
    .ZN(_12869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21817_ (.I(\sa21_sub[3] ),
    .ZN(_12870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21818_ (.A1(_12870_),
    .A2(\sa32_sub[3] ),
    .ZN(_12871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21819_ (.A1(_12869_),
    .A2(_12871_),
    .ZN(_12872_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21820_ (.A1(_12867_),
    .A2(_12872_),
    .ZN(_12873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21821_ (.A1(_12864_),
    .A2(net39),
    .ZN(_12874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21822_ (.A1(_12761_),
    .A2(\sa03_sr[2] ),
    .ZN(_12875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21823_ (.A1(_12874_),
    .A2(_12875_),
    .ZN(_12876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21824_ (.A1(_12870_),
    .A2(_12868_),
    .ZN(_12877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21825_ (.A1(\sa21_sub[3] ),
    .A2(\sa32_sub[3] ),
    .ZN(_12878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21826_ (.A1(_12877_),
    .A2(_12878_),
    .ZN(_12879_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21827_ (.A1(_12876_),
    .A2(_12879_),
    .ZN(_12880_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21828_ (.A1(_12873_),
    .A2(_12880_),
    .ZN(_12881_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21829_ (.I(\sa10_sub[3] ),
    .ZN(_12882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21830_ (.A1(_12882_),
    .A2(net772),
    .ZN(_12883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21831_ (.A1(net932),
    .A2(\sa10_sub[3] ),
    .ZN(_12884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21832_ (.A1(_12883_),
    .A2(_12884_),
    .ZN(_12885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21833_ (.A1(_12885_),
    .A2(\sa10_sub[2] ),
    .ZN(_12886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21834_ (.A1(net932),
    .A2(_12882_),
    .ZN(_12887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21835_ (.A1(net772),
    .A2(\sa10_sub[3] ),
    .ZN(_12888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21836_ (.A1(_12887_),
    .A2(_12888_),
    .ZN(_12889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21837_ (.A1(_12889_),
    .A2(_12841_),
    .ZN(_12890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21838_ (.A1(_12886_),
    .A2(_12890_),
    .ZN(_12891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21839_ (.A1(_12881_),
    .A2(_12891_),
    .ZN(_12892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21840_ (.A1(_12876_),
    .A2(_12879_),
    .ZN(_12893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21841_ (.A1(_12867_),
    .A2(_12872_),
    .ZN(_12894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21842_ (.A1(_12893_),
    .A2(_12894_),
    .ZN(_12895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21843_ (.A1(net932),
    .A2(_12841_),
    .ZN(_12896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21844_ (.A1(net772),
    .A2(\sa10_sub[2] ),
    .ZN(_12897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21845_ (.A1(_12896_),
    .A2(_12897_),
    .ZN(_12898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21846_ (.A1(_12898_),
    .A2(\sa10_sub[3] ),
    .ZN(_12899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21847_ (.A1(_12896_),
    .A2(_12882_),
    .A3(_12897_),
    .ZN(_12900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21848_ (.A1(_12899_),
    .A2(_12900_),
    .ZN(_12901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21849_ (.A1(_12895_),
    .A2(_12901_),
    .ZN(_12902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21850_ (.A1(_12892_),
    .A2(_12902_),
    .A3(_10405_),
    .ZN(_12903_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21851_ (.I(\u0.tmp_w[27] ),
    .ZN(_12904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21852_ (.A1(_12193_),
    .A2(\text_in_r[27] ),
    .ZN(_12905_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21853_ (.A1(_12903_),
    .A2(_12904_),
    .A3(_12905_),
    .ZN(_12906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21854_ (.A1(_12881_),
    .A2(_12901_),
    .ZN(_12907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21855_ (.A1(_12895_),
    .A2(_12891_),
    .ZN(_12908_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21856_ (.A1(_12907_),
    .A2(_12908_),
    .A3(_10405_),
    .ZN(_12909_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21857_ (.A1(_10522_),
    .A2(\text_in_r[27] ),
    .Z(_12910_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21858_ (.A1(_12909_),
    .A2(\u0.tmp_w[27] ),
    .A3(_12910_),
    .ZN(_12911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21859_ (.A1(_12906_),
    .A2(_12911_),
    .ZN(_12912_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21860_ (.I(_12912_),
    .Z(_12913_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _21861_ (.I(_12913_),
    .Z(_12914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21862_ (.A1(_12863_),
    .A2(_12914_),
    .ZN(_12915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21863_ (.A1(net626),
    .A2(_12803_),
    .ZN(_12916_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21864_ (.A1(net779),
    .A2(_12804_),
    .A3(_12802_),
    .ZN(_12917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21865_ (.A1(_12916_),
    .A2(_12917_),
    .ZN(_15770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21866_ (.A1(_12861_),
    .A2(net487),
    .ZN(_12918_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21867_ (.I(_12918_),
    .ZN(_12919_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21868_ (.A1(_12915_),
    .A2(_12919_),
    .Z(_12920_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21869_ (.A1(\sa10_sub[4] ),
    .A2(\sa32_sub[4] ),
    .ZN(_12921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21870_ (.A1(_12921_),
    .A2(_12889_),
    .ZN(_12922_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21871_ (.A1(\sa10_sub[4] ),
    .A2(\sa32_sub[4] ),
    .Z(_12923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21872_ (.A1(_12923_),
    .A2(_12885_),
    .ZN(_12924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21873_ (.A1(_12922_),
    .A2(_12924_),
    .ZN(_12925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21874_ (.I(_12925_),
    .ZN(_12926_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21875_ (.A1(\sa03_sr[7] ),
    .A2(\sa03_sr[3] ),
    .Z(_12927_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21876_ (.I(\sa21_sub[4] ),
    .ZN(_12928_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21877_ (.A1(_12927_),
    .A2(_12928_),
    .Z(_12929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21878_ (.A1(_12927_),
    .A2(_12928_),
    .ZN(_12930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21879_ (.A1(_12929_),
    .A2(_12930_),
    .ZN(_12931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21880_ (.A1(_12926_),
    .A2(_12931_),
    .ZN(_12932_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21881_ (.A1(_12927_),
    .A2(_12928_),
    .Z(_12933_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21882_ (.A1(_12927_),
    .A2(_12928_),
    .ZN(_12934_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21883_ (.A1(_12933_),
    .A2(_12934_),
    .ZN(_12935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21884_ (.A1(_12935_),
    .A2(_12925_),
    .ZN(_12936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21885_ (.A1(_12932_),
    .A2(_12936_),
    .A3(_10523_),
    .ZN(_12937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21886_ (.A1(_10526_),
    .A2(\text_in_r[28] ),
    .ZN(_12938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21887_ (.A1(_12937_),
    .A2(_12938_),
    .ZN(_12939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21888_ (.I(\u0.tmp_w[28] ),
    .ZN(_12940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21889_ (.A1(_12939_),
    .A2(_12940_),
    .ZN(_12941_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21890_ (.A1(_12937_),
    .A2(\u0.tmp_w[28] ),
    .A3(_12938_),
    .ZN(_12942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21891_ (.A1(_12942_),
    .A2(_12941_),
    .ZN(_12943_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _21892_ (.I(_12943_),
    .Z(_12944_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _21893_ (.I(_12944_),
    .Z(_12945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21894_ (.A1(net550),
    .A2(_12856_),
    .ZN(_12946_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21895_ (.I(_12912_),
    .ZN(_12947_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _21896_ (.I(_12947_),
    .Z(_12948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21897_ (.A1(_12946_),
    .A2(_12948_),
    .ZN(_12949_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21898_ (.I(_15785_),
    .ZN(_12950_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21899_ (.A1(_12851_),
    .A2(_12950_),
    .A3(_12855_),
    .ZN(_12951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21900_ (.I(_12951_),
    .ZN(_12952_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21901_ (.A1(_12949_),
    .A2(_12952_),
    .Z(_12953_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21902_ (.A1(_12920_),
    .A2(_12945_),
    .A3(_12953_),
    .ZN(_12954_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21903_ (.A1(\sa10_sub[4] ),
    .A2(\sa03_sr[4] ),
    .Z(_12955_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21904_ (.A1(\sa21_sub[5] ),
    .A2(\sa32_sub[5] ),
    .Z(_12956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21905_ (.A1(\sa21_sub[5] ),
    .A2(\sa32_sub[5] ),
    .ZN(_12957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21906_ (.A1(_12956_),
    .A2(_12957_),
    .ZN(_12958_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21907_ (.A1(\sa10_sub[5] ),
    .A2(_12958_),
    .Z(_12959_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21908_ (.A1(_12955_),
    .A2(_12959_),
    .Z(_12960_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21909_ (.I(_11385_),
    .Z(_12961_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21910_ (.I(\u0.tmp_w[29] ),
    .ZN(_12962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21911_ (.A1(_12961_),
    .A2(\text_in_r[29] ),
    .ZN(_12963_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21912_ (.A1(_12960_),
    .A2(_12961_),
    .B(_12962_),
    .C(_12963_),
    .ZN(_12964_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _21913_ (.I(_11348_),
    .Z(_12965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21914_ (.A1(_12960_),
    .A2(_12965_),
    .ZN(_12966_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21915_ (.A1(_10585_),
    .A2(\text_in_r[29] ),
    .Z(_12967_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21916_ (.A1(_12966_),
    .A2(\u0.tmp_w[29] ),
    .A3(_12967_),
    .ZN(_12968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21917_ (.A1(_12964_),
    .A2(_12968_),
    .ZN(_12969_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21918_ (.I(_12969_),
    .Z(_12970_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21919_ (.I(_12970_),
    .Z(_12971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21920_ (.A1(_15787_),
    .A2(_15773_),
    .Z(_12972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21921_ (.A1(_12972_),
    .A2(_12914_),
    .ZN(_12973_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21922_ (.I(_12943_),
    .ZN(_12974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21923_ (.A1(_12973_),
    .A2(_12974_),
    .ZN(_12975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21924_ (.A1(net486),
    .A2(_12862_),
    .ZN(_12976_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21925_ (.I(_12976_),
    .ZN(_12977_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _21926_ (.I(_12913_),
    .Z(_12978_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21927_ (.A1(_12977_),
    .A2(_12978_),
    .Z(_12979_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21928_ (.A1(_12975_),
    .A2(_12979_),
    .ZN(_12980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21929_ (.A1(net541),
    .A2(_12861_),
    .ZN(_12981_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _21930_ (.A1(net4),
    .A2(_12981_),
    .ZN(_12982_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21931_ (.A1(net966),
    .A2(_12949_),
    .Z(_12983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21932_ (.A1(_12980_),
    .A2(_12983_),
    .ZN(_12984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21933_ (.A1(_12954_),
    .A2(_12971_),
    .A3(_12984_),
    .ZN(_12985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21934_ (.A1(_12946_),
    .A2(net776),
    .ZN(_12986_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21935_ (.A1(_12986_),
    .A2(_12974_),
    .Z(_12987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21936_ (.I(_15776_),
    .ZN(_12988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21937_ (.A1(_12861_),
    .A2(_12988_),
    .ZN(_12989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21938_ (.A1(_12947_),
    .A2(_12989_),
    .Z(_12990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21939_ (.A1(_12990_),
    .A2(_12863_),
    .ZN(_12991_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21940_ (.I(_12969_),
    .Z(_12992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21941_ (.A1(_12987_),
    .A2(_12991_),
    .B(_12992_),
    .ZN(_12993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21942_ (.A1(net12),
    .A2(_15787_),
    .ZN(_12994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21943_ (.A1(_12863_),
    .A2(_12978_),
    .A3(_12994_),
    .ZN(_12995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21944_ (.I(_15772_),
    .ZN(_12996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21945_ (.A1(_12851_),
    .A2(_12855_),
    .A3(_12996_),
    .ZN(_12997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21946_ (.A1(_12997_),
    .A2(_12947_),
    .ZN(_12998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21947_ (.I(_12998_),
    .ZN(_12999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21948_ (.A1(_12862_),
    .A2(_12950_),
    .ZN(_13000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21949_ (.A1(_12999_),
    .A2(net965),
    .ZN(_13001_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21950_ (.I(_12944_),
    .Z(_13002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21951_ (.A1(_12995_),
    .A2(_13001_),
    .A3(_13002_),
    .ZN(_13003_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21952_ (.A1(\sa10_sub[5] ),
    .A2(\sa03_sr[5] ),
    .ZN(_13004_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21953_ (.A1(\sa21_sub[6] ),
    .A2(\sa32_sub[6] ),
    .Z(_13005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21954_ (.A1(\sa21_sub[6] ),
    .A2(\sa32_sub[6] ),
    .ZN(_13006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21955_ (.A1(_13005_),
    .A2(_13006_),
    .ZN(_13007_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21956_ (.A1(\sa10_sub[6] ),
    .A2(_13007_),
    .Z(_13008_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21957_ (.A1(_13004_),
    .A2(_13008_),
    .Z(_13009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _21958_ (.I(_11989_),
    .Z(_13010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21959_ (.A1(_10586_),
    .A2(\text_in_r[30] ),
    .Z(_13011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21960_ (.A1(_13009_),
    .A2(_13010_),
    .B(_13011_),
    .ZN(_13012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21961_ (.A1(_13012_),
    .A2(\u0.tmp_w[30] ),
    .Z(_13013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21962_ (.A1(_13012_),
    .A2(\u0.tmp_w[30] ),
    .ZN(_13014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21963_ (.A1(_13013_),
    .A2(_13014_),
    .Z(_13015_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21964_ (.I(_13015_),
    .Z(_13016_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21965_ (.I(_13016_),
    .Z(_13017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21966_ (.A1(_12993_),
    .A2(_13003_),
    .B(_13017_),
    .ZN(_13018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21967_ (.A1(_12985_),
    .A2(_13018_),
    .ZN(_13019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21968_ (.A1(_12981_),
    .A2(_12913_),
    .ZN(_13020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21969_ (.I(_13020_),
    .ZN(_13021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21970_ (.A1(net4),
    .A2(net12),
    .ZN(_13022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21971_ (.A1(_13021_),
    .A2(_13022_),
    .ZN(_13023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21972_ (.A1(_15775_),
    .A2(net556),
    .ZN(_13024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21973_ (.A1(_12862_),
    .A2(net542),
    .ZN(_13025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21974_ (.I(_12947_),
    .Z(_13026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21975_ (.A1(_13024_),
    .A2(_13025_),
    .A3(_13026_),
    .ZN(_13027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21976_ (.A1(_13023_),
    .A2(_12945_),
    .A3(_13027_),
    .ZN(_13028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21977_ (.A1(_12997_),
    .A2(_12914_),
    .Z(_13029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21978_ (.A1(net41),
    .A2(_15794_),
    .A3(net542),
    .ZN(_13030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21979_ (.A1(_13029_),
    .A2(_13030_),
    .ZN(_13031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21980_ (.I(_15771_),
    .ZN(_13032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21981_ (.A1(_15794_),
    .A2(_13032_),
    .ZN(_13033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21982_ (.I(_15779_),
    .ZN(_13034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21983_ (.A1(_15787_),
    .A2(net775),
    .ZN(_13035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21984_ (.A1(_13033_),
    .A2(_13035_),
    .ZN(_13036_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21985_ (.I(_12948_),
    .Z(_13037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21986_ (.A1(_13036_),
    .A2(_13037_),
    .ZN(_13038_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21987_ (.I(_12974_),
    .Z(_13039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21988_ (.A1(_13031_),
    .A2(_13038_),
    .A3(_13039_),
    .ZN(_13040_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21989_ (.A1(_12960_),
    .A2(_12961_),
    .B(\u0.tmp_w[29] ),
    .C(_12963_),
    .ZN(_13041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21990_ (.A1(_12966_),
    .A2(_12962_),
    .A3(_12967_),
    .ZN(_13042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21991_ (.A1(_13041_),
    .A2(_13042_),
    .ZN(_13043_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21992_ (.I(_13043_),
    .Z(_13044_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21993_ (.A1(_13028_),
    .A2(_13040_),
    .A3(_13044_),
    .ZN(_13045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21994_ (.A1(_12851_),
    .A2(_13032_),
    .A3(_12855_),
    .ZN(_13046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21995_ (.I(_13046_),
    .ZN(_13047_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _21996_ (.I(net776),
    .Z(_13048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21997_ (.A1(_13047_),
    .A2(_13048_),
    .B(_12944_),
    .ZN(_13049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21998_ (.A1(_15794_),
    .A2(_15771_),
    .ZN(_13050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21999_ (.A1(_12999_),
    .A2(_13050_),
    .ZN(_13051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22000_ (.A1(_15794_),
    .A2(_13034_),
    .Z(_13052_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22001_ (.I(_12914_),
    .Z(_13053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22002_ (.A1(_13052_),
    .A2(_13053_),
    .ZN(_13054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22003_ (.A1(_13049_),
    .A2(_13051_),
    .A3(_13054_),
    .ZN(_13055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22004_ (.A1(_12861_),
    .A2(_15772_),
    .ZN(_13056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22005_ (.A1(_13056_),
    .A2(net776),
    .ZN(_13057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22006_ (.A1(net769),
    .A2(_12862_),
    .ZN(_13058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22007_ (.I(_13058_),
    .ZN(_13059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22008_ (.A1(net972),
    .A2(_12862_),
    .ZN(_13060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22009_ (.A1(_13060_),
    .A2(_12948_),
    .ZN(_13061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22010_ (.A1(_13057_),
    .A2(_13059_),
    .B(_13061_),
    .ZN(_13062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22011_ (.A1(_13062_),
    .A2(_12945_),
    .ZN(_13063_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22012_ (.I(_12970_),
    .Z(_13064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22013_ (.A1(_13055_),
    .A2(_13063_),
    .A3(_13064_),
    .ZN(_13065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22014_ (.A1(_13045_),
    .A2(_13065_),
    .A3(_13017_),
    .ZN(_13066_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22015_ (.I(\sa32_sub[7] ),
    .Z(_13067_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22016_ (.A1(\sa03_sr[6] ),
    .A2(net50),
    .Z(_13068_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22017_ (.A1(net772),
    .A2(\sa10_sub[6] ),
    .Z(_13069_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22018_ (.A1(net54),
    .A2(_13068_),
    .A3(_13069_),
    .Z(_13070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22019_ (.I0(_13070_),
    .I1(\text_in_r[31] ),
    .S(_12961_),
    .Z(_13071_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _22020_ (.A1(_07739_),
    .A2(_13071_),
    .Z(_13072_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22021_ (.I(_13072_),
    .Z(_13073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22022_ (.A1(_13019_),
    .A2(_13066_),
    .A3(_13073_),
    .ZN(_13074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22023_ (.A1(_15794_),
    .A2(_12988_),
    .ZN(_13075_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _22024_ (.A1(_13024_),
    .A2(_15794_),
    .B(_13075_),
    .C(_13048_),
    .ZN(_13076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22025_ (.A1(_12862_),
    .A2(_15773_),
    .ZN(_13077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22026_ (.I(_13077_),
    .ZN(_13078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22027_ (.A1(_13078_),
    .A2(_12914_),
    .Z(_13079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22028_ (.I(_13079_),
    .ZN(_13080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22029_ (.I(_13025_),
    .ZN(_13081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _22030_ (.I(_12948_),
    .Z(_13082_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22031_ (.A1(_13081_),
    .A2(_13047_),
    .B(_13082_),
    .ZN(_13083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22032_ (.A1(_13076_),
    .A2(_13080_),
    .A3(_13083_),
    .ZN(_13084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22033_ (.A1(_12862_),
    .A2(net774),
    .ZN(_13085_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22034_ (.A1(_13085_),
    .A2(_13026_),
    .B(_12944_),
    .ZN(_13086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22035_ (.A1(_13026_),
    .A2(_15792_),
    .Z(_13087_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22036_ (.A1(_13086_),
    .A2(_13087_),
    .Z(_13088_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22037_ (.A1(_13084_),
    .A2(_12945_),
    .B(_13064_),
    .C(_13088_),
    .ZN(_13089_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22038_ (.I(_12975_),
    .ZN(_13090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22039_ (.A1(net769),
    .A2(_12861_),
    .ZN(_13091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22040_ (.I(_13091_),
    .ZN(_13092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22041_ (.A1(_13092_),
    .A2(net12),
    .ZN(_13093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22042_ (.I(_15781_),
    .ZN(_13094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22043_ (.A1(_13094_),
    .A2(_12862_),
    .ZN(_13095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22044_ (.A1(_12947_),
    .A2(_13095_),
    .ZN(_13096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22045_ (.I(_13096_),
    .ZN(_13097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22046_ (.A1(_13093_),
    .A2(_13097_),
    .ZN(_13098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22047_ (.A1(_13090_),
    .A2(_13098_),
    .B(_13064_),
    .ZN(_13099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22048_ (.A1(_12862_),
    .A2(_15779_),
    .ZN(_13100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22049_ (.A1(_12913_),
    .A2(_13100_),
    .ZN(_13101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22050_ (.I(_13101_),
    .ZN(_13102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22051_ (.A1(_13093_),
    .A2(_13102_),
    .ZN(_13103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22052_ (.A1(_12972_),
    .A2(_13026_),
    .ZN(_13104_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22053_ (.A1(_13103_),
    .A2(_13002_),
    .A3(_13104_),
    .ZN(_13105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _22054_ (.I(_13016_),
    .ZN(_13106_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22055_ (.I(_13106_),
    .Z(_13107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22056_ (.A1(_13099_),
    .A2(_13105_),
    .B(_13107_),
    .ZN(_13108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22057_ (.A1(_13089_),
    .A2(_13108_),
    .ZN(_13109_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22058_ (.I(_12944_),
    .Z(_13110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22059_ (.A1(net773),
    .A2(_13110_),
    .Z(_13111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22060_ (.A1(_15794_),
    .A2(_15776_),
    .ZN(_13112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22061_ (.A1(_12861_),
    .A2(_15781_),
    .ZN(_13113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22062_ (.A1(_13112_),
    .A2(_13113_),
    .ZN(_13114_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22063_ (.I(_12914_),
    .Z(_13115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22064_ (.A1(_13114_),
    .A2(_13115_),
    .ZN(_13116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22065_ (.A1(_13111_),
    .A2(_13116_),
    .B(_13043_),
    .ZN(_13117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22066_ (.I(_13112_),
    .ZN(_13118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _22067_ (.A1(_13118_),
    .A2(_13115_),
    .B(_13110_),
    .ZN(_13119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22068_ (.A1(_12983_),
    .A2(_13119_),
    .ZN(_13120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22069_ (.A1(_13117_),
    .A2(_13120_),
    .B(_13016_),
    .ZN(_13121_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22070_ (.I(_12974_),
    .Z(_13122_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22071_ (.A1(_12990_),
    .A2(_13122_),
    .ZN(_13123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22072_ (.I(_13033_),
    .ZN(_13124_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22073_ (.A1(_12972_),
    .A2(_13124_),
    .B(_13048_),
    .ZN(_13125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22074_ (.A1(_13123_),
    .A2(_13125_),
    .B(_12992_),
    .ZN(_13126_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22075_ (.A1(_13091_),
    .A2(net776),
    .Z(_13127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22076_ (.A1(_13127_),
    .A2(_13085_),
    .ZN(_13128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22077_ (.A1(_15787_),
    .A2(net538),
    .Z(_13129_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22078_ (.I(_12948_),
    .Z(_13130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22079_ (.A1(_13129_),
    .A2(_13052_),
    .B(_13130_),
    .ZN(_13131_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22080_ (.A1(_13128_),
    .A2(_13131_),
    .A3(_13039_),
    .ZN(_13132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22081_ (.A1(_13126_),
    .A2(_13132_),
    .ZN(_13133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22082_ (.A1(_13121_),
    .A2(_13133_),
    .B(_13072_),
    .ZN(_13134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22083_ (.A1(_13109_),
    .A2(_13134_),
    .ZN(_13135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22084_ (.A1(_13074_),
    .A2(_13135_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22085_ (.A1(_13000_),
    .A2(_12948_),
    .ZN(_13136_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22086_ (.A1(_13136_),
    .A2(_12919_),
    .ZN(_13137_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22087_ (.A1(_13122_),
    .A2(_13137_),
    .ZN(_13138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22088_ (.A1(net542),
    .A2(net770),
    .ZN(_13139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22089_ (.A1(_13139_),
    .A2(_15787_),
    .ZN(_13140_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _22090_ (.I(_12948_),
    .Z(_13141_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22091_ (.A1(_13140_),
    .A2(_13141_),
    .Z(_13142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22092_ (.A1(_13138_),
    .A2(_13142_),
    .ZN(_13143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22093_ (.A1(_13030_),
    .A2(_13141_),
    .A3(_13056_),
    .ZN(_13144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22094_ (.A1(_15787_),
    .A2(_15776_),
    .Z(_13145_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _22095_ (.I(_12944_),
    .Z(_13146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22096_ (.A1(_13145_),
    .A2(_13053_),
    .B(_13146_),
    .ZN(_13147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22097_ (.A1(_13144_),
    .A2(_13147_),
    .ZN(_13148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22098_ (.A1(_13143_),
    .A2(_13044_),
    .A3(_13148_),
    .ZN(_13149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22099_ (.A1(_12994_),
    .A2(net927),
    .ZN(_13150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22100_ (.A1(_13150_),
    .A2(_13037_),
    .ZN(_13151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22101_ (.A1(_12994_),
    .A2(_13085_),
    .A3(_13115_),
    .ZN(_13152_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22102_ (.A1(_13151_),
    .A2(_13152_),
    .A3(_13039_),
    .ZN(_13153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22103_ (.A1(_13025_),
    .A2(_13048_),
    .A3(_13046_),
    .ZN(_13154_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22104_ (.A1(_13112_),
    .A2(_12997_),
    .A3(_13026_),
    .ZN(_13155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22105_ (.A1(_13154_),
    .A2(_13155_),
    .ZN(_13156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22106_ (.A1(_13156_),
    .A2(_13002_),
    .ZN(_13157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22107_ (.A1(_13153_),
    .A2(_13157_),
    .A3(_13064_),
    .ZN(_13158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22108_ (.A1(_13149_),
    .A2(_13158_),
    .A3(_13107_),
    .ZN(_13159_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22109_ (.I(_12974_),
    .Z(_13160_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22110_ (.I(_13061_),
    .ZN(_13161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22111_ (.A1(_13161_),
    .A2(_12951_),
    .ZN(_13162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22112_ (.A1(_13076_),
    .A2(_13160_),
    .A3(_13162_),
    .ZN(_13163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22113_ (.A1(_13058_),
    .A2(_12947_),
    .ZN(_13164_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22114_ (.A1(_13164_),
    .A2(net970),
    .Z(_13165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _22115_ (.A1(_13118_),
    .A2(_13048_),
    .B(_12974_),
    .ZN(_13166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22116_ (.A1(_13165_),
    .A2(_13166_),
    .B(_13043_),
    .ZN(_13167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22117_ (.A1(_13163_),
    .A2(_13167_),
    .ZN(_13168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22118_ (.A1(_12999_),
    .A2(_12946_),
    .ZN(_13169_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22119_ (.A1(_13025_),
    .A2(_12989_),
    .A3(_13115_),
    .ZN(_13170_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22120_ (.I(_12944_),
    .Z(_13171_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22121_ (.A1(_13169_),
    .A2(_13170_),
    .A3(_13171_),
    .ZN(_13172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22122_ (.I(_13043_),
    .Z(_13173_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22123_ (.A1(_12861_),
    .A2(_12913_),
    .ZN(_13174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22124_ (.A1(_13024_),
    .A2(net933),
    .B(_13146_),
    .ZN(_13175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22125_ (.A1(_13091_),
    .A2(_13022_),
    .A3(_13048_),
    .ZN(_13176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22126_ (.A1(_13175_),
    .A2(_13176_),
    .ZN(_13177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22127_ (.A1(_13172_),
    .A2(_13173_),
    .A3(_13177_),
    .ZN(_13178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22128_ (.A1(_13178_),
    .A2(_13168_),
    .A3(_13017_),
    .ZN(_13179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22129_ (.A1(_13179_),
    .A2(_13159_),
    .B(_13073_),
    .ZN(_13180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22130_ (.A1(_13024_),
    .A2(_13174_),
    .ZN(_13181_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _22131_ (.A1(_13048_),
    .A2(_13140_),
    .B(_13181_),
    .ZN(_13182_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22132_ (.A1(_12994_),
    .A2(_13050_),
    .A3(_12978_),
    .ZN(_13183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22133_ (.I(_13183_),
    .ZN(_13184_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22134_ (.I(_12944_),
    .Z(_13185_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22135_ (.A1(_13182_),
    .A2(_13184_),
    .B(_13185_),
    .ZN(_13186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22136_ (.I(_12982_),
    .ZN(_13187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22137_ (.A1(_13187_),
    .A2(_13102_),
    .ZN(_13188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22138_ (.I(_13188_),
    .ZN(_13189_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22139_ (.I(_12974_),
    .Z(_13190_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22140_ (.I(_15795_),
    .ZN(_13191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22141_ (.A1(_13026_),
    .A2(_13191_),
    .ZN(_13192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22142_ (.A1(_12974_),
    .A2(_13192_),
    .B(_13043_),
    .ZN(_13193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22143_ (.A1(_13189_),
    .A2(_13190_),
    .B(_13193_),
    .ZN(_13194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22144_ (.A1(_13186_),
    .A2(_13194_),
    .ZN(_13195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22145_ (.A1(_13021_),
    .A2(_13058_),
    .ZN(_13196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22146_ (.A1(_13196_),
    .A2(_12970_),
    .Z(_13197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22147_ (.A1(_12990_),
    .A2(_12976_),
    .ZN(_13198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22148_ (.A1(_13198_),
    .A2(_12944_),
    .Z(_13199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22149_ (.A1(_13197_),
    .A2(_13199_),
    .B(_13106_),
    .ZN(_13200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22150_ (.A1(_13195_),
    .A2(_13200_),
    .ZN(_13201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22151_ (.A1(_13201_),
    .A2(_13073_),
    .ZN(_13202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22152_ (.A1(_13021_),
    .A2(_13050_),
    .ZN(_13203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22153_ (.A1(_13203_),
    .A2(_13198_),
    .A3(_13039_),
    .ZN(_13204_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22154_ (.A1(_13081_),
    .A2(_12972_),
    .B(_13115_),
    .ZN(_13205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22155_ (.A1(_13085_),
    .A2(_13046_),
    .ZN(_13206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22156_ (.A1(_13206_),
    .A2(_13130_),
    .ZN(_13207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22157_ (.A1(_13205_),
    .A2(_13171_),
    .A3(_13207_),
    .ZN(_13208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22158_ (.A1(_13204_),
    .A2(_13208_),
    .A3(_13173_),
    .ZN(_13209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22159_ (.A1(_12951_),
    .A2(_12914_),
    .Z(_13210_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22160_ (.I(_15773_),
    .ZN(_13211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22161_ (.A1(_15794_),
    .A2(_13211_),
    .ZN(_13212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22162_ (.A1(_13210_),
    .A2(_13212_),
    .ZN(_13213_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22163_ (.A1(_13144_),
    .A2(_13213_),
    .A3(_13171_),
    .ZN(_13214_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _22164_ (.A1(_12982_),
    .A2(_12986_),
    .B(_13190_),
    .C(net773),
    .ZN(_13215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22165_ (.A1(_13214_),
    .A2(_13064_),
    .A3(_13215_),
    .ZN(_13216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22166_ (.A1(_13216_),
    .A2(_13209_),
    .B(_13017_),
    .ZN(_13217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22167_ (.A1(_13217_),
    .A2(_13202_),
    .ZN(_13218_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22168_ (.A1(_13218_),
    .A2(_13180_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22169_ (.A1(_12994_),
    .A2(_13075_),
    .ZN(_13219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22170_ (.A1(_13219_),
    .A2(_13141_),
    .A3(_12918_),
    .ZN(_13220_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22171_ (.A1(_13220_),
    .A2(_13128_),
    .A3(_13190_),
    .Z(_13221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22172_ (.A1(_12989_),
    .A2(_12914_),
    .Z(_13222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22173_ (.A1(_13222_),
    .A2(net965),
    .ZN(_13223_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22174_ (.A1(_13024_),
    .A2(_13091_),
    .A3(_13141_),
    .ZN(_13224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22175_ (.A1(_13223_),
    .A2(_13224_),
    .B(_13039_),
    .ZN(_13225_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22176_ (.A1(_13221_),
    .A2(_13225_),
    .B(_12971_),
    .ZN(_13226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22177_ (.A1(_12863_),
    .A2(_13053_),
    .B(_13146_),
    .ZN(_13227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22178_ (.A1(_13030_),
    .A2(_13037_),
    .A3(_12951_),
    .ZN(_13228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22179_ (.A1(_13227_),
    .A2(_13228_),
    .B(_12992_),
    .ZN(_13229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22180_ (.I(_13057_),
    .ZN(_13230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22181_ (.A1(_13230_),
    .A2(_12976_),
    .ZN(_13231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22182_ (.I(_13231_),
    .ZN(_13232_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22183_ (.A1(_12981_),
    .A2(_13077_),
    .A3(_13026_),
    .Z(_13233_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22184_ (.A1(_13232_),
    .A2(_13233_),
    .B(_13002_),
    .ZN(_13234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22185_ (.A1(_13229_),
    .A2(_13234_),
    .B(_13106_),
    .ZN(_13235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22186_ (.A1(_13226_),
    .A2(_13235_),
    .ZN(_13236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22187_ (.A1(_15794_),
    .A2(_15785_),
    .ZN(_13237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22188_ (.I(_13237_),
    .ZN(_13238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22189_ (.A1(_13020_),
    .A2(_13238_),
    .B(_13146_),
    .ZN(_13239_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22190_ (.A1(_12976_),
    .A2(_13141_),
    .A3(_13113_),
    .Z(_13240_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22191_ (.A1(_13239_),
    .A2(_13240_),
    .ZN(_13241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22192_ (.A1(_12994_),
    .A2(_13095_),
    .A3(_13048_),
    .ZN(_13242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22193_ (.A1(_13085_),
    .A2(_12997_),
    .A3(_13082_),
    .ZN(_13243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22194_ (.A1(_13242_),
    .A2(_13243_),
    .B(_13185_),
    .ZN(_13244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22195_ (.A1(_13241_),
    .A2(_13244_),
    .B(_13044_),
    .ZN(_13245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22196_ (.A1(_13075_),
    .A2(_13026_),
    .ZN(_13246_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22197_ (.A1(_13246_),
    .A2(_12919_),
    .Z(_13247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22198_ (.A1(_13247_),
    .A2(_13160_),
    .A3(_13116_),
    .ZN(_13248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22199_ (.A1(_13113_),
    .A2(_13237_),
    .ZN(_13249_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22200_ (.I(_12978_),
    .Z(_13250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22201_ (.A1(_13249_),
    .A2(_13250_),
    .ZN(_13251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22202_ (.A1(_12994_),
    .A2(_13075_),
    .A3(_13082_),
    .ZN(_13252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22203_ (.A1(_13251_),
    .A2(_13252_),
    .A3(_13171_),
    .ZN(_13253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22204_ (.A1(_13248_),
    .A2(_13253_),
    .A3(_13064_),
    .ZN(_13254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22205_ (.A1(_13245_),
    .A2(_13254_),
    .A3(_13107_),
    .ZN(_13255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22206_ (.A1(_13236_),
    .A2(_13255_),
    .A3(_13073_),
    .ZN(_13256_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22207_ (.A1(_13211_),
    .A2(_12988_),
    .Z(_13257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22208_ (.A1(_15787_),
    .A2(_13257_),
    .ZN(_13258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22209_ (.A1(_13030_),
    .A2(_13130_),
    .A3(_13258_),
    .ZN(_13259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22210_ (.A1(_13188_),
    .A2(_13259_),
    .A3(_13002_),
    .ZN(_13260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22211_ (.A1(_12999_),
    .A2(_13075_),
    .ZN(_13261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22212_ (.A1(_13261_),
    .A2(_13049_),
    .B(_13106_),
    .ZN(_13262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22213_ (.A1(_13262_),
    .A2(_13260_),
    .B(_13064_),
    .ZN(_13263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22214_ (.A1(_13093_),
    .A2(_13161_),
    .ZN(_13264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22215_ (.A1(_15792_),
    .A2(_13053_),
    .B(_13146_),
    .ZN(_13265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22216_ (.A1(_13264_),
    .A2(_13265_),
    .B(_13016_),
    .ZN(_13266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22217_ (.A1(_13058_),
    .A2(net967),
    .ZN(_13267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22218_ (.A1(_13267_),
    .A2(_13130_),
    .ZN(_13268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22219_ (.A1(_13128_),
    .A2(_12945_),
    .A3(_13268_),
    .ZN(_13269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22220_ (.A1(_13266_),
    .A2(_13269_),
    .ZN(_13270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22221_ (.A1(_13270_),
    .A2(_13263_),
    .B(_13073_),
    .ZN(_13271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22222_ (.A1(_13127_),
    .A2(_13033_),
    .Z(_13272_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22223_ (.A1(_13085_),
    .A2(_13035_),
    .A3(_13141_),
    .Z(_13273_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22224_ (.A1(_13272_),
    .A2(_13273_),
    .B(_13002_),
    .ZN(_13274_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22225_ (.A1(_13091_),
    .A2(_13022_),
    .A3(_12948_),
    .Z(_13275_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22226_ (.A1(_13275_),
    .A2(_13110_),
    .ZN(_13276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22227_ (.A1(_13250_),
    .A2(_13191_),
    .ZN(_13277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22228_ (.A1(_13276_),
    .A2(_13277_),
    .ZN(_13278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22229_ (.A1(_13274_),
    .A2(_13278_),
    .A3(_13107_),
    .ZN(_13279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22230_ (.A1(_13053_),
    .A2(_15799_),
    .ZN(_13280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22231_ (.A1(_13224_),
    .A2(_13280_),
    .B(_13190_),
    .ZN(_13281_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22232_ (.A1(_12978_),
    .A2(_15790_),
    .Z(_13282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22233_ (.A1(_12915_),
    .A2(_13282_),
    .B(_13185_),
    .ZN(_13283_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22234_ (.A1(_13281_),
    .A2(_13283_),
    .B(_13017_),
    .ZN(_13284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22235_ (.A1(_13279_),
    .A2(_13284_),
    .A3(_12971_),
    .ZN(_13285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22236_ (.A1(_13285_),
    .A2(_13271_),
    .ZN(_13286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22237_ (.A1(_13286_),
    .A2(_13256_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _22238_ (.A1(_13141_),
    .A2(_12976_),
    .A3(_13025_),
    .A4(_13035_),
    .ZN(_13287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22239_ (.A1(_13085_),
    .A2(_12914_),
    .Z(_13288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22240_ (.A1(_13288_),
    .A2(_13140_),
    .ZN(_13289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22241_ (.A1(_13287_),
    .A2(_13190_),
    .A3(_13289_),
    .ZN(_13290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22242_ (.I(_13052_),
    .ZN(_13291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22243_ (.A1(_13029_),
    .A2(_13291_),
    .ZN(_13292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22244_ (.A1(_13292_),
    .A2(_13027_),
    .A3(_13185_),
    .ZN(_13293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22245_ (.A1(_13290_),
    .A2(_13293_),
    .ZN(_13294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22246_ (.A1(_13294_),
    .A2(_13044_),
    .ZN(_13295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22247_ (.A1(_12947_),
    .A2(_15787_),
    .Z(_13296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22248_ (.I(_13296_),
    .ZN(_13297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22249_ (.A1(_13024_),
    .A2(net967),
    .ZN(_13298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22250_ (.A1(_13297_),
    .A2(_13298_),
    .Z(_13299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22251_ (.A1(_13299_),
    .A2(_13160_),
    .B(_13173_),
    .ZN(_13300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22252_ (.A1(_13230_),
    .A2(_13095_),
    .ZN(_13301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22253_ (.A1(_13138_),
    .A2(_13301_),
    .ZN(_13302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22254_ (.A1(_13300_),
    .A2(_13302_),
    .B(_13017_),
    .ZN(_13303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22255_ (.A1(_13295_),
    .A2(_13303_),
    .ZN(_13304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22256_ (.A1(_13296_),
    .A2(_13032_),
    .B(_12970_),
    .ZN(_13305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22257_ (.A1(_13174_),
    .A2(net972),
    .Z(_13306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22258_ (.I(_13306_),
    .ZN(_13307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22259_ (.A1(_13025_),
    .A2(_13035_),
    .ZN(_13308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22260_ (.A1(_13308_),
    .A2(_13250_),
    .ZN(_13309_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22261_ (.A1(_13305_),
    .A2(_13307_),
    .A3(_13309_),
    .ZN(_13310_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22262_ (.A1(_13061_),
    .A2(_12970_),
    .Z(_13311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22263_ (.A1(_13267_),
    .A2(_13250_),
    .ZN(_13312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22264_ (.A1(_13311_),
    .A2(_13312_),
    .B(_13039_),
    .ZN(_13313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22265_ (.A1(_13310_),
    .A2(_13313_),
    .B(_13106_),
    .ZN(_13314_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22266_ (.A1(_13246_),
    .A2(_12952_),
    .Z(_13315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22267_ (.A1(_13315_),
    .A2(_13231_),
    .A3(_13173_),
    .ZN(_13316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22268_ (.A1(_13021_),
    .A2(_13024_),
    .ZN(_13317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22269_ (.A1(_12999_),
    .A2(_12976_),
    .ZN(_13318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22270_ (.A1(_13317_),
    .A2(_13318_),
    .A3(_13064_),
    .ZN(_13319_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22271_ (.A1(_13316_),
    .A2(_13319_),
    .A3(_13160_),
    .ZN(_13320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22272_ (.A1(_13320_),
    .A2(_13314_),
    .ZN(_13321_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22273_ (.I(_13072_),
    .ZN(_13322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22274_ (.A1(_13304_),
    .A2(_13321_),
    .A3(_13322_),
    .ZN(_13323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22275_ (.I(_13113_),
    .ZN(_13324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22276_ (.A1(_13130_),
    .A2(_13324_),
    .B(_12970_),
    .ZN(_13325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22277_ (.A1(_13325_),
    .A2(_13242_),
    .B(_13185_),
    .ZN(_13326_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22278_ (.I(_12986_),
    .ZN(_13327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22279_ (.A1(_13327_),
    .A2(_12997_),
    .ZN(_13328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22280_ (.A1(_13258_),
    .A2(_12948_),
    .Z(_13329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22281_ (.A1(_13329_),
    .A2(_13000_),
    .ZN(_13330_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22282_ (.A1(_13328_),
    .A2(_13330_),
    .A3(_12992_),
    .ZN(_13331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22283_ (.A1(_13326_),
    .A2(_13331_),
    .B(_13106_),
    .ZN(_13332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22284_ (.I(_12997_),
    .ZN(_13333_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22285_ (.A1(_13333_),
    .A2(_12978_),
    .Z(_13334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22286_ (.A1(_13334_),
    .A2(_13043_),
    .B1(_13037_),
    .B2(_12972_),
    .ZN(_13335_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22287_ (.A1(net973),
    .A2(_13092_),
    .ZN(_13336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22288_ (.A1(_13336_),
    .A2(_13306_),
    .B(_12970_),
    .ZN(_13337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22289_ (.A1(_13335_),
    .A2(_13337_),
    .ZN(_13338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22290_ (.A1(_13338_),
    .A2(_12945_),
    .ZN(_13339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22291_ (.A1(_13332_),
    .A2(_13339_),
    .B(_13322_),
    .ZN(_13340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22292_ (.A1(_13329_),
    .A2(_13095_),
    .ZN(_13341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22293_ (.A1(_13188_),
    .A2(_13341_),
    .B(_13185_),
    .ZN(_13342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22294_ (.I(_13239_),
    .ZN(_13343_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22295_ (.A1(_13342_),
    .A2(_13343_),
    .B(_12971_),
    .ZN(_13344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22296_ (.A1(_13083_),
    .A2(_13176_),
    .A3(_13160_),
    .ZN(_13345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22297_ (.A1(_13029_),
    .A2(_13000_),
    .ZN(_13346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22298_ (.A1(_12946_),
    .A2(_13113_),
    .ZN(_13347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22299_ (.A1(_13347_),
    .A2(_13026_),
    .ZN(_13348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22300_ (.A1(_13346_),
    .A2(_13348_),
    .A3(_13171_),
    .ZN(_13349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22301_ (.A1(_13345_),
    .A2(_13349_),
    .A3(_13173_),
    .ZN(_13350_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22302_ (.A1(_13344_),
    .A2(_13350_),
    .A3(_13107_),
    .ZN(_13351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22303_ (.A1(_13340_),
    .A2(_13351_),
    .ZN(_13352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22304_ (.A1(_13323_),
    .A2(_13352_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22305_ (.A1(_13093_),
    .A2(_13037_),
    .A3(_12976_),
    .ZN(_13353_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22306_ (.A1(_13353_),
    .A2(_12945_),
    .A3(_13223_),
    .ZN(_13354_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22307_ (.A1(_13059_),
    .A2(_13047_),
    .B(_13130_),
    .ZN(_13355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22308_ (.A1(_13076_),
    .A2(_13160_),
    .A3(_13355_),
    .ZN(_13356_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22309_ (.A1(_13354_),
    .A2(_13356_),
    .A3(_12971_),
    .ZN(_13357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22310_ (.A1(_13174_),
    .A2(_15772_),
    .Z(_13358_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22311_ (.A1(_13358_),
    .A2(_13324_),
    .ZN(_13359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22312_ (.A1(_13359_),
    .A2(_13166_),
    .B(_12992_),
    .ZN(_13360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22313_ (.A1(_13210_),
    .A2(_13060_),
    .ZN(_13361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22314_ (.A1(_13098_),
    .A2(_13361_),
    .A3(_13160_),
    .ZN(_13362_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22315_ (.A1(_13360_),
    .A2(_13362_),
    .B(_13106_),
    .ZN(_13363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22316_ (.A1(_13363_),
    .A2(_13357_),
    .ZN(_13364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22317_ (.A1(_12918_),
    .A2(_13139_),
    .ZN(_13365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22318_ (.A1(net970),
    .A2(_13050_),
    .A3(_13082_),
    .ZN(_13366_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22319_ (.A1(_13037_),
    .A2(_13365_),
    .B(_13366_),
    .C(_13171_),
    .ZN(_13367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22320_ (.A1(_13276_),
    .A2(_13196_),
    .ZN(_13368_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22321_ (.A1(_13367_),
    .A2(_13368_),
    .A3(_12971_),
    .ZN(_13369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22322_ (.I(_13164_),
    .ZN(_13370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22323_ (.A1(_13370_),
    .A2(_12994_),
    .ZN(_13371_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22324_ (.A1(_13371_),
    .A2(_13183_),
    .A3(_13160_),
    .ZN(_13372_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22325_ (.A1(_12972_),
    .A2(_13122_),
    .ZN(_13373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22326_ (.A1(_13373_),
    .A2(_13096_),
    .B(_12970_),
    .ZN(_13374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22327_ (.A1(_13372_),
    .A2(_13374_),
    .B(_13016_),
    .ZN(_13375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22328_ (.A1(_13369_),
    .A2(_13375_),
    .ZN(_13376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22329_ (.A1(_13364_),
    .A2(_13376_),
    .A3(_13322_),
    .ZN(_13377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22330_ (.A1(_12976_),
    .A2(_13046_),
    .Z(_13378_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22331_ (.A1(_13378_),
    .A2(_13082_),
    .Z(_13379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22332_ (.A1(_13199_),
    .A2(_13379_),
    .ZN(_13380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22333_ (.A1(_13021_),
    .A2(net965),
    .ZN(_13381_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22334_ (.A1(_13174_),
    .A2(_13146_),
    .ZN(_13382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22335_ (.A1(_13381_),
    .A2(_13382_),
    .B(_13173_),
    .ZN(_13383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22336_ (.A1(_13380_),
    .A2(_13383_),
    .ZN(_13384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22337_ (.A1(_13250_),
    .A2(_13212_),
    .B(_13122_),
    .ZN(_13385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22338_ (.A1(_13030_),
    .A2(_13037_),
    .ZN(_13386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22339_ (.A1(_13385_),
    .A2(_13386_),
    .B(_12992_),
    .ZN(_13387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22340_ (.A1(_13222_),
    .A2(_13085_),
    .ZN(_13388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22341_ (.A1(_12983_),
    .A2(_13388_),
    .A3(_13039_),
    .ZN(_13389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22342_ (.A1(_13387_),
    .A2(_13389_),
    .ZN(_13390_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22343_ (.A1(_13384_),
    .A2(_13390_),
    .A3(_13107_),
    .ZN(_13391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22344_ (.A1(_13129_),
    .A2(net776),
    .ZN(_13392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22345_ (.A1(_13392_),
    .A2(_13110_),
    .Z(_13393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22346_ (.A1(_13097_),
    .A2(net970),
    .ZN(_13394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22347_ (.A1(_12919_),
    .A2(_13250_),
    .ZN(_13395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22348_ (.A1(_13394_),
    .A2(_13393_),
    .A3(_13395_),
    .ZN(_13396_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22349_ (.I(_15783_),
    .ZN(_13397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22350_ (.A1(_13397_),
    .A2(_13115_),
    .B(_13110_),
    .ZN(_13398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22351_ (.A1(_13085_),
    .A2(_13130_),
    .ZN(_13399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22352_ (.A1(_13398_),
    .A2(_13399_),
    .B(_12970_),
    .ZN(_13400_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22353_ (.A1(_13396_),
    .A2(_13400_),
    .B(_13106_),
    .ZN(_13401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22354_ (.A1(_13097_),
    .A2(net967),
    .ZN(_13402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22355_ (.A1(_13048_),
    .A2(_13365_),
    .ZN(_13403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22356_ (.A1(_13402_),
    .A2(net930),
    .A3(_13002_),
    .ZN(_13404_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22357_ (.A1(_13125_),
    .A2(_13039_),
    .A3(_13027_),
    .ZN(_13405_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22358_ (.A1(_13404_),
    .A2(_13405_),
    .A3(_13064_),
    .ZN(_13406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22359_ (.A1(_13406_),
    .A2(_13401_),
    .ZN(_13407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22360_ (.A1(_13391_),
    .A2(_13407_),
    .A3(_13073_),
    .ZN(_13408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22361_ (.A1(_13377_),
    .A2(_13408_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22362_ (.A1(_13140_),
    .A2(_13141_),
    .A3(_13291_),
    .Z(_13409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22363_ (.A1(_13327_),
    .A2(net927),
    .ZN(_13410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22364_ (.A1(_13410_),
    .A2(_13185_),
    .ZN(_13411_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22365_ (.A1(_13409_),
    .A2(_13411_),
    .ZN(_13412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22366_ (.A1(_13141_),
    .A2(net928),
    .ZN(_13413_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22367_ (.A1(_13403_),
    .A2(_13190_),
    .A3(_13413_),
    .Z(_13414_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22368_ (.A1(_13412_),
    .A2(_13414_),
    .B(_13044_),
    .ZN(_13415_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22369_ (.A1(_13091_),
    .A2(_12978_),
    .A3(_13212_),
    .Z(_13416_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22370_ (.A1(_13416_),
    .A2(_13358_),
    .B(_13185_),
    .ZN(_13417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22371_ (.A1(_13237_),
    .A2(_13048_),
    .ZN(_13418_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22372_ (.A1(_13124_),
    .A2(net773),
    .B(_13418_),
    .C(_13190_),
    .ZN(_13419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22373_ (.A1(_13417_),
    .A2(_13419_),
    .ZN(_13420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22374_ (.A1(_13420_),
    .A2(_12971_),
    .ZN(_13421_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22375_ (.A1(_13415_),
    .A2(_13421_),
    .A3(_13017_),
    .ZN(_13422_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22376_ (.A1(_13222_),
    .A2(_13122_),
    .ZN(_13423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22377_ (.A1(_13423_),
    .A2(_13181_),
    .B(_13043_),
    .ZN(_13424_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22378_ (.I(_13029_),
    .ZN(_13425_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22379_ (.A1(_13348_),
    .A2(_13039_),
    .A3(_13425_),
    .ZN(_13426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22380_ (.A1(_13424_),
    .A2(_13426_),
    .B(_13016_),
    .ZN(_13427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22381_ (.I(_13136_),
    .ZN(_13428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22382_ (.A1(_13428_),
    .A2(_12989_),
    .ZN(_13429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22383_ (.A1(_12980_),
    .A2(_13429_),
    .ZN(_13430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22384_ (.A1(_13095_),
    .A2(_12914_),
    .Z(_13431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22385_ (.A1(_13093_),
    .A2(_13431_),
    .ZN(_13432_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22386_ (.A1(_13246_),
    .A2(_13257_),
    .Z(_13433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22387_ (.A1(_13432_),
    .A2(_13433_),
    .A3(_13171_),
    .ZN(_13434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22388_ (.A1(_13430_),
    .A2(_13434_),
    .A3(_13044_),
    .ZN(_13435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22389_ (.A1(_13427_),
    .A2(_13435_),
    .B(_13073_),
    .ZN(_13436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22390_ (.A1(_13422_),
    .A2(_13436_),
    .ZN(_13437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22391_ (.I(_13329_),
    .ZN(_13438_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22392_ (.A1(_12915_),
    .A2(net966),
    .B(_13438_),
    .C(_13039_),
    .ZN(_13439_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22393_ (.A1(_13166_),
    .A2(_13136_),
    .B(_12992_),
    .ZN(_13440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22394_ (.A1(_13439_),
    .A2(_13440_),
    .ZN(_13441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22395_ (.A1(_13187_),
    .A2(_13250_),
    .ZN(_13442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22396_ (.A1(net775),
    .A2(_13130_),
    .B(_13146_),
    .ZN(_13443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22397_ (.A1(_13442_),
    .A2(_13443_),
    .B(_13173_),
    .ZN(_13444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22398_ (.A1(_13230_),
    .A2(_13000_),
    .ZN(_13445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22399_ (.A1(_12999_),
    .A2(_13100_),
    .ZN(_13446_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22400_ (.A1(_13445_),
    .A2(_13446_),
    .A3(_13002_),
    .ZN(_13447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22401_ (.A1(_13444_),
    .A2(_13447_),
    .ZN(_13448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22402_ (.A1(_13441_),
    .A2(_13448_),
    .A3(_13017_),
    .ZN(_13449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22403_ (.A1(net539),
    .A2(_13082_),
    .B(_13110_),
    .ZN(_13450_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22404_ (.A1(_13023_),
    .A2(_13450_),
    .B(_12992_),
    .ZN(_13451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22405_ (.A1(_13431_),
    .A2(_12918_),
    .ZN(_13452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22406_ (.A1(_12999_),
    .A2(_12863_),
    .ZN(_13453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22407_ (.A1(_13452_),
    .A2(_13453_),
    .A3(_13171_),
    .ZN(_13454_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22408_ (.A1(_13454_),
    .A2(_13451_),
    .B(_13016_),
    .ZN(_13455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22409_ (.A1(_12983_),
    .A2(_13119_),
    .A3(_13392_),
    .ZN(_13456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22410_ (.A1(_13187_),
    .A2(_13250_),
    .A3(net965),
    .ZN(_13457_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22411_ (.A1(_13052_),
    .A2(_13130_),
    .B(_13122_),
    .ZN(_13458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22412_ (.A1(_13457_),
    .A2(_13458_),
    .ZN(_13459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22413_ (.A1(_13456_),
    .A2(_13459_),
    .A3(_13064_),
    .ZN(_13460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22414_ (.A1(_13455_),
    .A2(_13460_),
    .ZN(_13461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22415_ (.A1(_13461_),
    .A2(_13449_),
    .A3(_13073_),
    .ZN(_13462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22416_ (.A1(_13462_),
    .A2(_13437_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22417_ (.A1(_13095_),
    .A2(_12951_),
    .A3(_12978_),
    .ZN(_13463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22418_ (.A1(net926),
    .A2(_13174_),
    .ZN(_13464_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22419_ (.A1(_13463_),
    .A2(_13104_),
    .A3(_13464_),
    .ZN(_13465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22420_ (.A1(_13465_),
    .A2(_13190_),
    .ZN(_13466_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _22421_ (.A1(_13141_),
    .A2(_13112_),
    .A3(_13077_),
    .A4(_13113_),
    .ZN(_13467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22422_ (.I(_13392_),
    .ZN(_13468_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22423_ (.A1(_13086_),
    .A2(_13468_),
    .ZN(_13469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22424_ (.A1(_13467_),
    .A2(_13469_),
    .ZN(_13470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22425_ (.A1(_13466_),
    .A2(_13470_),
    .ZN(_13471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22426_ (.A1(_13471_),
    .A2(_12971_),
    .ZN(_13472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22427_ (.A1(_13077_),
    .A2(_13113_),
    .Z(_13473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22428_ (.A1(_13047_),
    .A2(_13115_),
    .ZN(_13474_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22429_ (.A1(_13473_),
    .A2(_13250_),
    .B(_13171_),
    .C(_13474_),
    .ZN(_13475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22430_ (.A1(_13365_),
    .A2(_13082_),
    .ZN(_13476_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22431_ (.A1(_15788_),
    .A2(_15797_),
    .B(_13115_),
    .ZN(_13477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22432_ (.A1(_13476_),
    .A2(_13160_),
    .A3(_13477_),
    .ZN(_13478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22433_ (.A1(_13475_),
    .A2(_13478_),
    .A3(_13044_),
    .ZN(_13479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22434_ (.A1(_13472_),
    .A2(_13479_),
    .A3(_13107_),
    .ZN(_13480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22435_ (.A1(net4),
    .A2(_15787_),
    .B(_12978_),
    .ZN(_13481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22436_ (.A1(_13481_),
    .A2(_12863_),
    .ZN(_13482_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22437_ (.A1(_13056_),
    .A2(_13212_),
    .A3(_13115_),
    .ZN(_13483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22438_ (.A1(_13482_),
    .A2(_13483_),
    .B(_13185_),
    .ZN(_13484_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22439_ (.A1(_13082_),
    .A2(_12997_),
    .B(_13110_),
    .ZN(_13485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22440_ (.A1(_12915_),
    .A2(_13282_),
    .B(_13485_),
    .ZN(_13486_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22441_ (.A1(_13484_),
    .A2(_13486_),
    .B(_13044_),
    .ZN(_13487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22442_ (.A1(_13370_),
    .A2(_13024_),
    .ZN(_13488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22443_ (.A1(_13052_),
    .A2(_13053_),
    .B(_13122_),
    .ZN(_13489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22444_ (.A1(_13488_),
    .A2(_13489_),
    .B(_13043_),
    .ZN(_13490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22445_ (.A1(_13288_),
    .A2(_13258_),
    .B(_13146_),
    .ZN(_13491_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22446_ (.A1(_13093_),
    .A2(_13037_),
    .A3(_13025_),
    .ZN(_13492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22447_ (.A1(_13491_),
    .A2(_13492_),
    .ZN(_13493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22448_ (.A1(_13490_),
    .A2(_13493_),
    .ZN(_13494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22449_ (.A1(_13487_),
    .A2(_13017_),
    .A3(_13494_),
    .ZN(_13495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22450_ (.A1(_13480_),
    .A2(_13495_),
    .A3(_13322_),
    .ZN(_13496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22451_ (.A1(_13164_),
    .A2(_12944_),
    .Z(_13497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22452_ (.A1(_12995_),
    .A2(_13497_),
    .ZN(_13498_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22453_ (.A1(_13056_),
    .A2(_12948_),
    .Z(_13499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22454_ (.A1(_13348_),
    .A2(_13122_),
    .A3(_13499_),
    .ZN(_13500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22455_ (.A1(_13498_),
    .A2(_13500_),
    .ZN(_13501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22456_ (.A1(_13501_),
    .A2(_13106_),
    .ZN(_13502_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22457_ (.A1(_13096_),
    .A2(_12919_),
    .B(net973),
    .ZN(_13503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22458_ (.A1(_13503_),
    .A2(_13185_),
    .ZN(_13504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22459_ (.A1(_13220_),
    .A2(_13190_),
    .ZN(_13505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22460_ (.A1(_13504_),
    .A2(_13505_),
    .A3(_13016_),
    .ZN(_13506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22461_ (.A1(_13502_),
    .A2(_13506_),
    .ZN(_13507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22462_ (.A1(_13507_),
    .A2(_12971_),
    .ZN(_13508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22463_ (.A1(net929),
    .A2(_12978_),
    .ZN(_13509_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22464_ (.A1(_13298_),
    .A2(_12974_),
    .A3(_13509_),
    .Z(_13510_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22465_ (.A1(_13510_),
    .A2(_13016_),
    .ZN(_13511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22466_ (.A1(_13022_),
    .A2(_13026_),
    .Z(_13512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22467_ (.A1(_13512_),
    .A2(_13210_),
    .B(_13025_),
    .ZN(_13513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22468_ (.A1(_13513_),
    .A2(_12945_),
    .ZN(_13514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22469_ (.A1(_13511_),
    .A2(_13514_),
    .ZN(_13515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22470_ (.A1(_13081_),
    .A2(_13053_),
    .B(_13122_),
    .ZN(_13516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22471_ (.A1(_13428_),
    .A2(_13056_),
    .ZN(_13517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22472_ (.A1(_13516_),
    .A2(_13517_),
    .ZN(_13518_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22473_ (.I(_15789_),
    .ZN(_13519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22474_ (.A1(_13519_),
    .A2(_13082_),
    .B(_13110_),
    .ZN(_13520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22475_ (.A1(_13452_),
    .A2(_13520_),
    .ZN(_13521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22476_ (.A1(_13518_),
    .A2(_13521_),
    .A3(_13016_),
    .ZN(_13522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22477_ (.A1(_13515_),
    .A2(_13522_),
    .A3(_13044_),
    .ZN(_13523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22478_ (.A1(_13508_),
    .A2(_13073_),
    .A3(_13523_),
    .ZN(_13524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22479_ (.A1(_13496_),
    .A2(_13524_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22480_ (.A1(_13296_),
    .A2(net926),
    .B(_13146_),
    .ZN(_13525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22481_ (.I(_13334_),
    .ZN(_13526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22482_ (.A1(_13525_),
    .A2(_13526_),
    .B(_13173_),
    .ZN(_13527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22483_ (.A1(_13093_),
    .A2(_13037_),
    .ZN(_13528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22484_ (.A1(_13230_),
    .A2(_13030_),
    .ZN(_13529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22485_ (.A1(_13528_),
    .A2(_13529_),
    .A3(_12945_),
    .ZN(_13530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22486_ (.A1(_13527_),
    .A2(_13530_),
    .B(_13107_),
    .ZN(_13531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22487_ (.A1(_13030_),
    .A2(_13250_),
    .A3(net969),
    .ZN(_13532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22488_ (.A1(_13276_),
    .A2(_13532_),
    .ZN(_13533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22489_ (.A1(_13115_),
    .A2(net12),
    .ZN(_13534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22490_ (.A1(_13371_),
    .A2(_13534_),
    .ZN(_13535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22491_ (.A1(_13535_),
    .A2(_12945_),
    .ZN(_13536_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22492_ (.A1(_13533_),
    .A2(_13536_),
    .A3(_13044_),
    .ZN(_13537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22493_ (.A1(_13531_),
    .A2(_13537_),
    .ZN(_13538_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22494_ (.A1(_13328_),
    .A2(_13162_),
    .A3(_13002_),
    .ZN(_13539_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22495_ (.A1(_13268_),
    .A2(_13160_),
    .A3(_13463_),
    .ZN(_13540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22496_ (.A1(_13539_),
    .A2(_13540_),
    .A3(_12971_),
    .ZN(_13541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22497_ (.A1(_13093_),
    .A2(_13327_),
    .B(_13122_),
    .ZN(_13542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22498_ (.A1(_12976_),
    .A2(_12946_),
    .ZN(_13543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22499_ (.A1(_13543_),
    .A2(_13047_),
    .B(_13037_),
    .ZN(_13544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22500_ (.A1(_13542_),
    .A2(_13544_),
    .ZN(_13545_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22501_ (.A1(_13210_),
    .A2(_13146_),
    .ZN(_13546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22502_ (.A1(_13394_),
    .A2(_13546_),
    .B(_12992_),
    .ZN(_13547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22503_ (.A1(_13545_),
    .A2(_13547_),
    .ZN(_13548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22504_ (.A1(_13541_),
    .A2(_13548_),
    .A3(_13107_),
    .ZN(_13549_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22505_ (.A1(_13538_),
    .A2(_13549_),
    .A3(_13073_),
    .ZN(_13550_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22506_ (.A1(_13378_),
    .A2(_13327_),
    .Z(_13551_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22507_ (.A1(_12999_),
    .A2(_13291_),
    .Z(_13552_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22508_ (.A1(_13552_),
    .A2(_13551_),
    .B(_13173_),
    .ZN(_13553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22509_ (.A1(_12970_),
    .A2(_13046_),
    .ZN(_13554_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22510_ (.A1(_13079_),
    .A2(_13554_),
    .ZN(_13555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22511_ (.A1(net933),
    .A2(net4),
    .ZN(_13556_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22512_ (.A1(_13555_),
    .A2(_13556_),
    .B(_13171_),
    .ZN(_13557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22513_ (.A1(_13557_),
    .A2(_13553_),
    .ZN(_13558_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22514_ (.A1(_13543_),
    .A2(_12919_),
    .B(_13053_),
    .ZN(_13559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22515_ (.A1(_13559_),
    .A2(_13173_),
    .A3(_13341_),
    .ZN(_13560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22516_ (.A1(_15776_),
    .A2(_13053_),
    .B(_13043_),
    .ZN(_13561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22517_ (.A1(_13561_),
    .A2(_13476_),
    .B(_13190_),
    .ZN(_13562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22518_ (.A1(_13560_),
    .A2(_13562_),
    .ZN(_13563_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22519_ (.A1(_13563_),
    .A2(_13558_),
    .A3(_13107_),
    .ZN(_13564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22520_ (.A1(_13392_),
    .A2(_13509_),
    .Z(_13565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22521_ (.A1(_13199_),
    .A2(_13565_),
    .ZN(_13566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22522_ (.A1(_13397_),
    .A2(_13130_),
    .B(_13110_),
    .ZN(_13567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22523_ (.A1(_13080_),
    .A2(_13567_),
    .B(_12992_),
    .ZN(_13568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22524_ (.A1(_13566_),
    .A2(_13568_),
    .ZN(_13569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22525_ (.A1(_13327_),
    .A2(net970),
    .ZN(_13570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22526_ (.A1(_13161_),
    .A2(_13056_),
    .ZN(_13571_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22527_ (.A1(_13570_),
    .A2(_13571_),
    .A3(_13002_),
    .ZN(_13572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22528_ (.A1(_15797_),
    .A2(_13082_),
    .B(_13110_),
    .ZN(_13573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22529_ (.A1(_13060_),
    .A2(_13113_),
    .ZN(_13574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22530_ (.A1(_13574_),
    .A2(_13053_),
    .ZN(_13575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22531_ (.A1(_13573_),
    .A2(_13575_),
    .B(_13043_),
    .ZN(_13576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22532_ (.A1(_13572_),
    .A2(_13576_),
    .ZN(_13577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22533_ (.A1(_13569_),
    .A2(_13577_),
    .A3(_13017_),
    .ZN(_13578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22534_ (.A1(_13322_),
    .A2(_13578_),
    .A3(_13564_),
    .ZN(_13579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22535_ (.A1(_13550_),
    .A2(_13579_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22536_ (.I(\sa20_sr[7] ),
    .ZN(_13580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22537_ (.A1(_13580_),
    .A2(net1073),
    .ZN(_13581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22538_ (.A1(_10394_),
    .A2(_10634_),
    .ZN(_13582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22539_ (.A1(_13581_),
    .A2(_13582_),
    .ZN(_13583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22540_ (.A1(_10354_),
    .A2(_13583_),
    .ZN(_13584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22541_ (.A1(_10394_),
    .A2(_13580_),
    .ZN(_13585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22542_ (.A1(\sa20_sr[0] ),
    .A2(_10634_),
    .ZN(_13586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22543_ (.A1(_13585_),
    .A2(_13586_),
    .ZN(_13587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22544_ (.A1(_10347_),
    .A2(_13587_),
    .ZN(_13588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22545_ (.A1(_13584_),
    .A2(_13588_),
    .Z(_13589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22546_ (.A1(_10362_),
    .A2(_10414_),
    .ZN(_13590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22547_ (.A1(_10366_),
    .A2(\sa00_sr[1] ),
    .ZN(_13591_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22548_ (.A1(_13591_),
    .A2(_13590_),
    .Z(_13592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22549_ (.A1(_13589_),
    .A2(_13592_),
    .ZN(_13593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22550_ (.A1(_13584_),
    .A2(_13588_),
    .ZN(_13594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22551_ (.A1(_13590_),
    .A2(_13591_),
    .ZN(_13595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22552_ (.A1(_13595_),
    .A2(_13594_),
    .ZN(_13596_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22553_ (.A1(_13593_),
    .A2(_13596_),
    .A3(net811),
    .ZN(_13597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22554_ (.A1(_10381_),
    .A2(\text_in_r[113] ),
    .ZN(_13598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22555_ (.A1(_13597_),
    .A2(_13598_),
    .ZN(_13599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22556_ (.I(\u0.w[0][17] ),
    .ZN(_13600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22557_ (.A1(_13599_),
    .A2(_13600_),
    .ZN(_13601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22558_ (.A1(net673),
    .A2(\u0.w[0][17] ),
    .A3(_13598_),
    .ZN(_13602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22559_ (.A1(_13602_),
    .A2(_13601_),
    .ZN(_15807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22560_ (.A1(net681),
    .A2(net581),
    .ZN(_13603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22561_ (.A1(_10391_),
    .A2(_10358_),
    .ZN(_13604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22562_ (.A1(_13603_),
    .A2(_13604_),
    .ZN(_13605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22563_ (.A1(_13605_),
    .A2(net75),
    .ZN(_13606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22564_ (.A1(_13603_),
    .A2(_13604_),
    .A3(_10339_),
    .ZN(_13607_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22565_ (.A1(_13606_),
    .A2(_13607_),
    .A3(net1138),
    .ZN(_13608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22566_ (.A1(net75),
    .A2(_10358_),
    .ZN(_13609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22567_ (.I(_13609_),
    .ZN(_13610_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22568_ (.A1(net75),
    .A2(_10358_),
    .ZN(_13611_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22569_ (.A1(_13610_),
    .A2(_13611_),
    .B(net582),
    .ZN(_13612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22570_ (.A1(_10339_),
    .A2(net681),
    .ZN(_13613_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22571_ (.A1(_13613_),
    .A2(_10391_),
    .A3(_13609_),
    .ZN(_13614_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22572_ (.A1(_13587_),
    .A2(_13614_),
    .A3(_13612_),
    .ZN(_13615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _22573_ (.A1(_13608_),
    .A2(net868),
    .B(_11203_),
    .ZN(_13616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22574_ (.I(\text_in_r[112] ),
    .ZN(_13617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22575_ (.A1(_13617_),
    .A2(_10431_),
    .Z(_13618_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22576_ (.A1(_13616_),
    .A2(_13618_),
    .B(\u0.w[0][16] ),
    .ZN(_13619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22577_ (.A1(net869),
    .A2(_13608_),
    .ZN(_13620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22578_ (.A1(_11989_),
    .A2(_13620_),
    .ZN(_13621_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22579_ (.I(\u0.w[0][16] ),
    .ZN(_13622_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22580_ (.I(_13618_),
    .ZN(_13623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22581_ (.A1(_13621_),
    .A2(_13622_),
    .A3(_13623_),
    .ZN(_13624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22582_ (.A1(_13624_),
    .A2(_13619_),
    .ZN(_15810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22583_ (.A1(\sa20_sr[2] ),
    .A2(\sa30_sr[2] ),
    .ZN(_13625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22584_ (.I(_13625_),
    .ZN(_13626_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22585_ (.A1(\sa20_sr[2] ),
    .A2(\sa30_sr[2] ),
    .ZN(_13627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22586_ (.A1(_13626_),
    .A2(_13627_),
    .B(\sa00_sr[2] ),
    .ZN(_13628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22587_ (.A1(_10417_),
    .A2(_10423_),
    .ZN(_13629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22588_ (.A1(_13629_),
    .A2(_10450_),
    .A3(_13625_),
    .ZN(_13630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22589_ (.A1(_13628_),
    .A2(_13630_),
    .ZN(_13631_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _22590_ (.A1(net614),
    .A2(\sa10_sr[1] ),
    .ZN(_13632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22591_ (.I(_13632_),
    .ZN(_13633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22592_ (.A1(_13631_),
    .A2(_13633_),
    .ZN(_13634_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22593_ (.A1(_13628_),
    .A2(_13630_),
    .A3(_13632_),
    .ZN(_13635_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22594_ (.A1(net811),
    .A2(_13635_),
    .A3(_13634_),
    .ZN(_13636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22595_ (.A1(_10431_),
    .A2(\text_in_r[114] ),
    .ZN(_13637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22596_ (.A1(_13637_),
    .A2(_13636_),
    .ZN(_13638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22597_ (.A1(_13638_),
    .A2(\u0.w[0][18] ),
    .ZN(_13639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22598_ (.I(\u0.w[0][18] ),
    .ZN(_13640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22599_ (.A1(_13636_),
    .A2(_13640_),
    .A3(_13637_),
    .ZN(_13641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22600_ (.A1(_13641_),
    .A2(_13639_),
    .ZN(_13642_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22601_ (.I(_13642_),
    .Z(_15826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _22602_ (.A1(_13616_),
    .A2(_13618_),
    .B(_13622_),
    .ZN(_13643_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22603_ (.A1(_13623_),
    .A2(\u0.w[0][16] ),
    .A3(_13621_),
    .ZN(_13644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22604_ (.A1(_13643_),
    .A2(_13644_),
    .ZN(_15801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22605_ (.A1(_13638_),
    .A2(_13640_),
    .ZN(_13645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22606_ (.A1(_13636_),
    .A2(\u0.w[0][18] ),
    .A3(_13637_),
    .ZN(_13646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22607_ (.A1(_13646_),
    .A2(_13645_),
    .ZN(_13647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22608_ (.I(_13647_),
    .Z(_15819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22609_ (.I(\sa30_sr[4] ),
    .ZN(_13648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22610_ (.A1(_10512_),
    .A2(_13648_),
    .ZN(_13649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22611_ (.A1(\sa20_sr[4] ),
    .A2(\sa30_sr[4] ),
    .ZN(_13650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22612_ (.A1(_13649_),
    .A2(_13650_),
    .ZN(_13651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22613_ (.A1(_10458_),
    .A2(_13580_),
    .ZN(_13652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22614_ (.A1(\sa20_sr[3] ),
    .A2(net47),
    .ZN(_13653_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22615_ (.A1(_13651_),
    .A2(_13652_),
    .A3(_13653_),
    .ZN(_13654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22616_ (.A1(_13652_),
    .A2(_13653_),
    .ZN(_13655_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22617_ (.A1(_13655_),
    .A2(_13650_),
    .A3(_13649_),
    .ZN(_13656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22618_ (.A1(_13654_),
    .A2(_13656_),
    .Z(_13657_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22619_ (.A1(\sa00_sr[4] ),
    .A2(_10473_),
    .Z(_13658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22620_ (.A1(_13657_),
    .A2(_13658_),
    .ZN(_13659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22621_ (.A1(_13654_),
    .A2(_13656_),
    .ZN(_13660_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22622_ (.A1(\sa00_sr[4] ),
    .A2(_10469_),
    .Z(_13661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22623_ (.A1(_13660_),
    .A2(_13661_),
    .ZN(_13662_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22624_ (.A1(_13659_),
    .A2(_13662_),
    .A3(_10523_),
    .ZN(_13663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22625_ (.A1(_10526_),
    .A2(\text_in_r[116] ),
    .ZN(_13664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22626_ (.A1(_13663_),
    .A2(_13664_),
    .ZN(_13665_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22627_ (.I(\u0.w[0][20] ),
    .ZN(_13666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22628_ (.A1(_13665_),
    .A2(_13666_),
    .ZN(_13667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22629_ (.A1(_13663_),
    .A2(\u0.w[0][20] ),
    .A3(_13664_),
    .ZN(_13668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22630_ (.A1(_13667_),
    .A2(_13668_),
    .ZN(_13669_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22631_ (.I(_13669_),
    .Z(_13670_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22632_ (.I(_13670_),
    .Z(_13671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22633_ (.I(_15803_),
    .ZN(_13672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22634_ (.A1(_15826_),
    .A2(_13672_),
    .Z(_13673_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22635_ (.I(_15811_),
    .ZN(_13674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22636_ (.A1(_15819_),
    .A2(_13674_),
    .ZN(_13675_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22637_ (.I(_13675_),
    .ZN(_13676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22638_ (.A1(_10417_),
    .A2(_13580_),
    .ZN(_13677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22639_ (.A1(\sa20_sr[2] ),
    .A2(_10634_),
    .ZN(_13678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22640_ (.A1(_13677_),
    .A2(_13678_),
    .ZN(_13679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22641_ (.A1(_10449_),
    .A2(_13679_),
    .ZN(_13680_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22642_ (.A1(\sa20_sr[2] ),
    .A2(_10634_),
    .Z(_13681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22643_ (.A1(_13681_),
    .A2(_10462_),
    .ZN(_13682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22644_ (.A1(_13680_),
    .A2(_13682_),
    .ZN(_13683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22645_ (.I(_13683_),
    .ZN(_13684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22646_ (.A1(net682),
    .A2(_10425_),
    .ZN(_13685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22647_ (.A1(net46),
    .A2(\sa10_sr[2] ),
    .ZN(_13686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22648_ (.A1(_13685_),
    .A2(_13686_),
    .ZN(_13687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22649_ (.A1(_13687_),
    .A2(\sa00_sr[3] ),
    .ZN(_13688_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22650_ (.I(\sa00_sr[3] ),
    .ZN(_13689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22651_ (.A1(_13685_),
    .A2(_13689_),
    .A3(_13686_),
    .ZN(_13690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22652_ (.A1(_13688_),
    .A2(_13690_),
    .ZN(_13691_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22653_ (.I(_13691_),
    .ZN(_13692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22654_ (.A1(_13684_),
    .A2(_13692_),
    .ZN(_13693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22655_ (.A1(_13683_),
    .A2(_13691_),
    .ZN(_13694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22656_ (.A1(_13693_),
    .A2(_11989_),
    .A3(_13694_),
    .ZN(_13695_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22657_ (.A1(_10586_),
    .A2(\text_in_r[115] ),
    .ZN(_13696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22658_ (.A1(_13695_),
    .A2(_13696_),
    .ZN(_13697_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22659_ (.I(\u0.w[0][19] ),
    .ZN(_13698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22660_ (.A1(_13697_),
    .A2(_13698_),
    .ZN(_13699_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22661_ (.A1(_13695_),
    .A2(\u0.w[0][19] ),
    .A3(_13696_),
    .ZN(_13700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22662_ (.A1(_13699_),
    .A2(_13700_),
    .ZN(_13701_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22663_ (.I(_13701_),
    .Z(_13702_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22664_ (.I(_13702_),
    .Z(_13703_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22665_ (.A1(_13673_),
    .A2(_13676_),
    .B(_13703_),
    .ZN(_13704_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22666_ (.I(_15804_),
    .ZN(_13705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22667_ (.A1(_13705_),
    .A2(net674),
    .ZN(_13706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22668_ (.A1(_13697_),
    .A2(\u0.w[0][19] ),
    .ZN(_13707_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22669_ (.A1(_13695_),
    .A2(_13698_),
    .A3(_13696_),
    .ZN(_13708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22670_ (.A1(_13707_),
    .A2(_13708_),
    .ZN(_13709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22671_ (.A1(_13709_),
    .A2(_13706_),
    .Z(_13710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22672_ (.A1(net28),
    .A2(net666),
    .A3(_15826_),
    .ZN(_13711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22673_ (.A1(_13710_),
    .A2(_13711_),
    .ZN(_13712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22674_ (.A1(_13704_),
    .A2(_13712_),
    .ZN(_13713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22675_ (.A1(net686),
    .A2(net660),
    .ZN(_13714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22676_ (.I(_13709_),
    .Z(_13715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22677_ (.A1(_13714_),
    .A2(_13715_),
    .Z(_13716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22678_ (.A1(\u0.w[0][17] ),
    .A2(_13599_),
    .ZN(_13717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22679_ (.A1(_13598_),
    .A2(_13600_),
    .A3(net673),
    .ZN(_13718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22680_ (.A1(_13718_),
    .A2(_13717_),
    .ZN(_15802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22681_ (.A1(net19),
    .A2(net83),
    .ZN(_13719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22682_ (.A1(_13716_),
    .A2(_13719_),
    .ZN(_13720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22683_ (.A1(net657),
    .A2(net671),
    .ZN(_13721_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22684_ (.I(_13701_),
    .Z(_13722_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _22685_ (.I(_13642_),
    .Z(_13723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22686_ (.A1(net665),
    .A2(_13723_),
    .ZN(_13724_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22687_ (.A1(_13721_),
    .A2(_13722_),
    .A3(_13724_),
    .ZN(_13725_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22688_ (.I(_13670_),
    .Z(_13726_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22689_ (.A1(_13720_),
    .A2(_13725_),
    .A3(_13726_),
    .ZN(_13727_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22690_ (.I(\sa00_sr[5] ),
    .ZN(_13728_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22691_ (.A1(_13728_),
    .A2(_10545_),
    .Z(_13729_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _22692_ (.A1(\sa10_sr[4] ),
    .A2(\sa20_sr[4] ),
    .ZN(_13730_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22693_ (.I(_13730_),
    .ZN(_13731_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22694_ (.A1(_13729_),
    .A2(_13731_),
    .Z(_13732_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22695_ (.A1(_13729_),
    .A2(_13731_),
    .ZN(_13733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22696_ (.A1(_10411_),
    .A2(\text_in_r[117] ),
    .ZN(_13734_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _22697_ (.A1(_13732_),
    .A2(_10526_),
    .A3(_13733_),
    .B(_13734_),
    .ZN(_13735_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22698_ (.A1(_13735_),
    .A2(\u0.w[0][21] ),
    .Z(_13736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22699_ (.A1(_13735_),
    .A2(\u0.w[0][21] ),
    .ZN(_13737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22700_ (.A1(_13736_),
    .A2(_13737_),
    .ZN(_13738_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22701_ (.I(_13738_),
    .ZN(_13739_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22702_ (.I(_13739_),
    .Z(_13740_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22703_ (.A1(_13671_),
    .A2(_13713_),
    .B(_13727_),
    .C(_13740_),
    .ZN(_13741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22704_ (.I(\sa00_sr[6] ),
    .ZN(_13742_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22705_ (.A1(_13742_),
    .A2(_10582_),
    .Z(_13743_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22706_ (.A1(\sa10_sr[5] ),
    .A2(\sa20_sr[5] ),
    .A3(_13743_),
    .Z(_13744_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22707_ (.A1(_10483_),
    .A2(\text_in_r[118] ),
    .Z(_13745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22708_ (.A1(_13744_),
    .A2(_11348_),
    .B(_13745_),
    .ZN(_13746_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22709_ (.A1(\u0.w[0][22] ),
    .A2(_13746_),
    .Z(_13747_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22710_ (.I(_13747_),
    .Z(_13748_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22711_ (.I(_13748_),
    .Z(_13749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22712_ (.A1(net872),
    .A2(_13705_),
    .ZN(_13750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22713_ (.A1(_13750_),
    .A2(_13702_),
    .ZN(_13751_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22714_ (.A1(_13751_),
    .A2(_13670_),
    .Z(_13752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22715_ (.A1(net672),
    .A2(net19),
    .ZN(_13753_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22716_ (.I(_13753_),
    .ZN(_13754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22717_ (.A1(_13754_),
    .A2(_13715_),
    .ZN(_13755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22718_ (.I(_13706_),
    .ZN(_13756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22719_ (.I(_13709_),
    .Z(_13757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22720_ (.A1(_13757_),
    .A2(_13756_),
    .ZN(_13758_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22721_ (.A1(_13752_),
    .A2(_13755_),
    .A3(_13758_),
    .Z(_13759_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22722_ (.A1(_15826_),
    .A2(_13674_),
    .Z(_13760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22723_ (.A1(net686),
    .A2(_13672_),
    .ZN(_13761_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22724_ (.I(_13761_),
    .ZN(_13762_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22725_ (.I(_13715_),
    .Z(_13763_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22726_ (.A1(_13760_),
    .A2(_13762_),
    .B(_13763_),
    .ZN(_13764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22727_ (.A1(_13701_),
    .A2(_13706_),
    .ZN(_13765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _22728_ (.I(_13765_),
    .ZN(_13766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22729_ (.A1(_15826_),
    .A2(_15803_),
    .ZN(_13767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22730_ (.A1(_13766_),
    .A2(_13767_),
    .ZN(_13768_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22731_ (.I(_13669_),
    .Z(_13769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22732_ (.A1(_13768_),
    .A2(_13764_),
    .B(_13769_),
    .ZN(_13770_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22733_ (.I(_13738_),
    .Z(_13771_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22734_ (.I(_13771_),
    .Z(_13772_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22735_ (.A1(_13770_),
    .A2(_13759_),
    .B(_13772_),
    .ZN(_13773_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22736_ (.A1(_13741_),
    .A2(_13773_),
    .A3(_13749_),
    .ZN(_13774_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _22737_ (.I(_13714_),
    .ZN(_13775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22738_ (.A1(net28),
    .A2(_13775_),
    .ZN(_13776_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22739_ (.I(_13701_),
    .Z(_13777_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22740_ (.I(_13777_),
    .Z(_13778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22741_ (.A1(net872),
    .A2(net670),
    .ZN(_13779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22742_ (.A1(_13776_),
    .A2(_13778_),
    .A3(_13779_),
    .ZN(_13780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22743_ (.I(_15805_),
    .ZN(_13781_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22744_ (.A1(net672),
    .A2(_13781_),
    .ZN(_13782_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22745_ (.A1(_13715_),
    .A2(_13782_),
    .B(_13670_),
    .ZN(_13783_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22746_ (.A1(_13780_),
    .A2(_13755_),
    .A3(_13783_),
    .ZN(_13784_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22747_ (.I(_15817_),
    .ZN(_13785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22748_ (.A1(net675),
    .A2(_13785_),
    .ZN(_13786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22749_ (.A1(_13786_),
    .A2(_13777_),
    .Z(_13787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22750_ (.A1(_13665_),
    .A2(\u0.w[0][20] ),
    .ZN(_13788_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22751_ (.A1(_13663_),
    .A2(_13666_),
    .A3(_13664_),
    .ZN(_13789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22752_ (.A1(_13788_),
    .A2(_13789_),
    .ZN(_13790_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22753_ (.I(_13790_),
    .Z(_13791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22754_ (.A1(_13787_),
    .A2(_13779_),
    .B(_13791_),
    .ZN(_13792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22755_ (.A1(net19),
    .A2(_13647_),
    .ZN(_13793_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22756_ (.I(_13793_),
    .Z(_13794_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22757_ (.A1(_13794_),
    .A2(_13757_),
    .Z(_13795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22758_ (.A1(net872),
    .A2(net671),
    .A3(net656),
    .ZN(_13796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22759_ (.A1(_13795_),
    .A2(net1132),
    .ZN(_13797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22760_ (.A1(_13792_),
    .A2(_13797_),
    .ZN(_13798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22761_ (.A1(_13784_),
    .A2(_13772_),
    .A3(_13798_),
    .ZN(_13799_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22762_ (.A1(net661),
    .A2(net686),
    .ZN(_13800_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22763_ (.A1(_13777_),
    .A2(_13800_),
    .ZN(_13801_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22764_ (.A1(_13801_),
    .A2(_13769_),
    .ZN(_13802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22765_ (.I(_15808_),
    .ZN(_13803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22766_ (.A1(_15819_),
    .A2(_13803_),
    .ZN(_13804_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22767_ (.A1(_13804_),
    .A2(_13777_),
    .Z(_13805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22768_ (.A1(_13805_),
    .A2(_13796_),
    .ZN(_13806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22769_ (.A1(_13802_),
    .A2(_13806_),
    .B(_13771_),
    .ZN(_13807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22770_ (.A1(net83),
    .A2(_15819_),
    .ZN(_13808_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22771_ (.A1(_13808_),
    .A2(_13715_),
    .Z(_13809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22772_ (.A1(_13809_),
    .A2(_13796_),
    .ZN(_13810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22773_ (.A1(_13785_),
    .A2(net872),
    .ZN(_13811_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22774_ (.A1(_13811_),
    .A2(_13701_),
    .Z(_13812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22775_ (.A1(_13812_),
    .A2(net659),
    .ZN(_13813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22776_ (.A1(_13810_),
    .A2(_13813_),
    .A3(_13726_),
    .ZN(_13814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22777_ (.A1(_13807_),
    .A2(_13814_),
    .B(_13748_),
    .ZN(_13815_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22778_ (.A1(net76),
    .A2(\sa10_sr[6] ),
    .A3(\sa20_sr[6] ),
    .Z(_13816_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22779_ (.A1(net47),
    .A2(net68),
    .A3(_13816_),
    .Z(_13817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22780_ (.A1(_10639_),
    .A2(\text_in_r[119] ),
    .Z(_13818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22781_ (.A1(_13817_),
    .A2(_12965_),
    .B(_13818_),
    .ZN(_13819_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _22782_ (.A1(\u0.w[0][23] ),
    .A2(_13819_),
    .Z(_13820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22783_ (.I(_13820_),
    .ZN(_13821_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22784_ (.I(_13821_),
    .Z(_13822_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22785_ (.A1(_13799_),
    .A2(_13815_),
    .B(_13822_),
    .ZN(_13823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22786_ (.A1(_13774_),
    .A2(_13823_),
    .ZN(_13824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22787_ (.A1(_13721_),
    .A2(_15819_),
    .A3(_13715_),
    .ZN(_13825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22788_ (.A1(_13723_),
    .A2(_15808_),
    .ZN(_13826_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _22789_ (.A1(_13826_),
    .A2(_13777_),
    .Z(_13827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22790_ (.A1(_13825_),
    .A2(_13827_),
    .Z(_13828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22791_ (.A1(_13724_),
    .A2(_13761_),
    .Z(_13829_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22792_ (.I(_13709_),
    .Z(_13830_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22793_ (.A1(_13829_),
    .A2(_13830_),
    .Z(_13831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22794_ (.A1(_13723_),
    .A2(_15805_),
    .ZN(_13832_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22795_ (.A1(_13832_),
    .A2(_13777_),
    .Z(_13833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22796_ (.A1(_13833_),
    .A2(_13790_),
    .Z(_13834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22797_ (.A1(_13828_),
    .A2(_13831_),
    .A3(_13834_),
    .ZN(_13835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22798_ (.A1(net668),
    .A2(net672),
    .ZN(_13836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22799_ (.I(_13836_),
    .ZN(_13837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _22800_ (.A1(_13837_),
    .A2(_13830_),
    .B(_13790_),
    .ZN(_13838_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22801_ (.I(_13702_),
    .Z(_13839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22802_ (.A1(_13839_),
    .A2(_15824_),
    .ZN(_13840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22803_ (.A1(_13838_),
    .A2(_13840_),
    .B(_13740_),
    .ZN(_13841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22804_ (.A1(_13835_),
    .A2(_13841_),
    .ZN(_13842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22805_ (.A1(net657),
    .A2(net686),
    .ZN(_13843_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22806_ (.I(_13843_),
    .ZN(_13844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22807_ (.A1(_13844_),
    .A2(net693),
    .ZN(_13845_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22808_ (.I(_15813_),
    .ZN(_13846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22809_ (.A1(_13723_),
    .A2(_13846_),
    .ZN(_13847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22810_ (.A1(_13847_),
    .A2(_13777_),
    .Z(_13848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22811_ (.A1(_13845_),
    .A2(_13848_),
    .ZN(_13849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22812_ (.A1(_13849_),
    .A2(_13783_),
    .ZN(_13850_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22813_ (.A1(_13723_),
    .A2(_15811_),
    .ZN(_13851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22814_ (.A1(_13851_),
    .A2(_13715_),
    .ZN(_13852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22815_ (.I(_13852_),
    .ZN(_13853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22816_ (.A1(net871),
    .A2(_13853_),
    .ZN(_13854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22817_ (.A1(_13782_),
    .A2(_13777_),
    .ZN(_13855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22818_ (.A1(_13670_),
    .A2(_13855_),
    .ZN(_13856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22819_ (.I(_13856_),
    .ZN(_13857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22820_ (.A1(_13854_),
    .A2(_13857_),
    .ZN(_13858_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22821_ (.A1(_13850_),
    .A2(_13858_),
    .A3(_13740_),
    .ZN(_13859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22822_ (.A1(_13842_),
    .A2(_13859_),
    .A3(_13749_),
    .ZN(_13860_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22823_ (.A1(_15826_),
    .A2(_13846_),
    .ZN(_13861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22824_ (.A1(_13861_),
    .A2(_13715_),
    .ZN(_13862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22825_ (.A1(_13862_),
    .A2(_13670_),
    .Z(_13863_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22826_ (.A1(_13863_),
    .A2(_13765_),
    .A3(_13827_),
    .ZN(_13864_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22827_ (.I(_13790_),
    .Z(_13865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22828_ (.A1(_13827_),
    .A2(_13865_),
    .Z(_13866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22829_ (.A1(_13780_),
    .A2(_13866_),
    .ZN(_13867_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22830_ (.I(_13771_),
    .Z(_13868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22831_ (.A1(_13864_),
    .A2(_13867_),
    .A3(_13868_),
    .ZN(_13869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22832_ (.A1(_13843_),
    .A2(_13709_),
    .ZN(_13870_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22833_ (.I(_13870_),
    .ZN(_13871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22834_ (.A1(_13871_),
    .A2(net680),
    .ZN(_13872_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22835_ (.I(_13865_),
    .Z(_13873_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22836_ (.I(_13702_),
    .Z(_13874_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22837_ (.A1(_13775_),
    .A2(_13760_),
    .B(_13874_),
    .ZN(_13875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22838_ (.A1(_13872_),
    .A2(_13873_),
    .A3(_13875_),
    .ZN(_13876_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22839_ (.A1(_13805_),
    .A2(_13791_),
    .ZN(_13877_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22840_ (.A1(_13673_),
    .A2(_13782_),
    .B(_13763_),
    .ZN(_13878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22841_ (.A1(_13877_),
    .A2(_13878_),
    .B(_13771_),
    .ZN(_13879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22842_ (.A1(_13876_),
    .A2(_13879_),
    .ZN(_13880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22843_ (.I(_13748_),
    .ZN(_13881_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22844_ (.I(_13881_),
    .Z(_13882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22845_ (.A1(_13869_),
    .A2(_13880_),
    .A3(_13882_),
    .ZN(_13883_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22846_ (.A1(_13860_),
    .A2(_13883_),
    .A3(_13822_),
    .ZN(_13884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22847_ (.A1(_13824_),
    .A2(_13884_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22848_ (.A1(net28),
    .A2(net694),
    .B(_13779_),
    .C(_13874_),
    .ZN(_13885_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22849_ (.I(_13865_),
    .Z(_13886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22850_ (.A1(_13836_),
    .A2(_13757_),
    .Z(_13887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22851_ (.A1(_13887_),
    .A2(_13808_),
    .ZN(_13888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22852_ (.A1(_13885_),
    .A2(_13886_),
    .A3(_13888_),
    .ZN(_13889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22853_ (.A1(_13829_),
    .A2(_13763_),
    .ZN(_13890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22854_ (.A1(_13766_),
    .A2(_13826_),
    .ZN(_13891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22855_ (.A1(_13890_),
    .A2(_13891_),
    .ZN(_13892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22856_ (.A1(_13892_),
    .A2(_13671_),
    .ZN(_13893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22857_ (.A1(_13889_),
    .A2(_13893_),
    .A3(_13772_),
    .ZN(_13894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22858_ (.A1(_13793_),
    .A2(_13808_),
    .ZN(_13895_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22859_ (.I(_13715_),
    .Z(_13896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22860_ (.A1(_13895_),
    .A2(_13896_),
    .ZN(_13897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22861_ (.A1(_13812_),
    .A2(_13794_),
    .ZN(_13898_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22862_ (.I(_13670_),
    .Z(_13899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22863_ (.A1(_13897_),
    .A2(_13898_),
    .A3(_13899_),
    .ZN(_13900_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22864_ (.I(_13739_),
    .Z(_13901_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22865_ (.I(_13901_),
    .Z(_13902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22866_ (.A1(net669),
    .A2(_15819_),
    .ZN(_13903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22867_ (.A1(_13711_),
    .A2(_13874_),
    .A3(_13903_),
    .ZN(_13904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22868_ (.A1(_15819_),
    .A2(_15808_),
    .ZN(_13905_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22869_ (.I(_13905_),
    .ZN(_13906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _22870_ (.I(_13669_),
    .Z(_13907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22871_ (.A1(_13906_),
    .A2(_13896_),
    .B(_13907_),
    .ZN(_13908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22872_ (.A1(_13904_),
    .A2(_13908_),
    .ZN(_13909_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22873_ (.A1(_13900_),
    .A2(_13902_),
    .A3(_13909_),
    .ZN(_13910_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22874_ (.A1(_13894_),
    .A2(_13910_),
    .A3(_13882_),
    .ZN(_13911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22875_ (.A1(_13766_),
    .A2(_13779_),
    .ZN(_13912_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22876_ (.A1(_13804_),
    .A2(_13709_),
    .Z(_13913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22877_ (.A1(_13913_),
    .A2(_13724_),
    .ZN(_13914_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22878_ (.A1(_13912_),
    .A2(_13914_),
    .A3(_13671_),
    .ZN(_13915_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22879_ (.A1(_13777_),
    .A2(_15826_),
    .Z(_13916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22880_ (.A1(_13916_),
    .A2(_13721_),
    .B(_13769_),
    .ZN(_13917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22881_ (.A1(_13871_),
    .A2(_13719_),
    .ZN(_13918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22882_ (.A1(_13917_),
    .A2(_13918_),
    .ZN(_13919_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22883_ (.A1(_13915_),
    .A2(_13919_),
    .A3(_13902_),
    .ZN(_13920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22884_ (.A1(_13827_),
    .A2(_13794_),
    .Z(_13921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22885_ (.A1(net658),
    .A2(_15826_),
    .ZN(_13922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22886_ (.A1(_13922_),
    .A2(_13778_),
    .B(_13865_),
    .ZN(_13923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22887_ (.A1(_13921_),
    .A2(_13923_),
    .B(_13740_),
    .ZN(_13924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22888_ (.A1(_13787_),
    .A2(_13750_),
    .ZN(_13925_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22889_ (.A1(_13925_),
    .A2(_13791_),
    .Z(_13926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22890_ (.A1(_13926_),
    .A2(_13828_),
    .ZN(_13927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22891_ (.A1(_13924_),
    .A2(_13927_),
    .ZN(_13928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22892_ (.A1(_13920_),
    .A2(_13928_),
    .A3(_13749_),
    .ZN(_13929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22893_ (.A1(_13911_),
    .A2(_13929_),
    .A3(_13822_),
    .ZN(_13930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22894_ (.A1(_13776_),
    .A2(net1132),
    .A3(_13703_),
    .ZN(_13931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22895_ (.A1(_13809_),
    .A2(_13767_),
    .ZN(_13932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22896_ (.A1(_13931_),
    .A2(_13740_),
    .A3(_13932_),
    .ZN(_13933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22897_ (.A1(_13716_),
    .A2(_13922_),
    .ZN(_13934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22898_ (.A1(_13805_),
    .A2(net867),
    .ZN(_13935_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22899_ (.I(_13738_),
    .Z(_13936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22900_ (.A1(_13934_),
    .A2(_13935_),
    .A3(_13936_),
    .ZN(_13937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22901_ (.A1(_13933_),
    .A2(_13937_),
    .B(_13886_),
    .ZN(_13938_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22902_ (.A1(_13901_),
    .A2(_15827_),
    .A3(_13763_),
    .Z(_13939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22903_ (.A1(_13776_),
    .A2(_13853_),
    .ZN(_13940_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22904_ (.A1(_13939_),
    .A2(_13886_),
    .A3(_13940_),
    .Z(_13941_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22905_ (.A1(_13938_),
    .A2(_13941_),
    .B(_13749_),
    .ZN(_13942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22906_ (.A1(_13776_),
    .A2(_13801_),
    .ZN(_13943_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22907_ (.A1(_13765_),
    .A2(_13865_),
    .Z(_13944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22908_ (.A1(_13943_),
    .A2(_13944_),
    .B(_13901_),
    .ZN(_13945_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22909_ (.A1(_13786_),
    .A2(_13715_),
    .Z(_13946_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22910_ (.A1(_15826_),
    .A2(_13781_),
    .ZN(_13947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22911_ (.A1(_13946_),
    .A2(_13947_),
    .B(_13791_),
    .ZN(_13948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22912_ (.A1(_13948_),
    .A2(_13904_),
    .ZN(_13949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22913_ (.A1(_13945_),
    .A2(_13949_),
    .B(_13748_),
    .ZN(_13950_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22914_ (.A1(_13724_),
    .A2(_13702_),
    .Z(_13951_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22915_ (.A1(_13951_),
    .A2(_13670_),
    .Z(_13952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22916_ (.A1(_13837_),
    .A2(_13722_),
    .ZN(_13953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22917_ (.A1(_13782_),
    .A2(_13757_),
    .ZN(_13954_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22918_ (.A1(_13953_),
    .A2(_13954_),
    .Z(_13955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22919_ (.A1(_13762_),
    .A2(_13703_),
    .ZN(_13956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22920_ (.A1(_13952_),
    .A2(_13955_),
    .A3(_13956_),
    .ZN(_13957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22921_ (.A1(_13716_),
    .A2(_13767_),
    .ZN(_13958_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _22922_ (.I(_13790_),
    .Z(_13959_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22923_ (.A1(_13958_),
    .A2(_13935_),
    .A3(_13959_),
    .ZN(_13960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22924_ (.A1(_13957_),
    .A2(_13740_),
    .A3(_13960_),
    .ZN(_13961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22925_ (.A1(_13950_),
    .A2(_13961_),
    .B(_13821_),
    .ZN(_13962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22926_ (.A1(_13942_),
    .A2(_13962_),
    .ZN(_13963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22927_ (.A1(_13930_),
    .A2(_13963_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22928_ (.A1(_13808_),
    .A2(_13847_),
    .A3(_13757_),
    .ZN(_13964_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22929_ (.A1(_13706_),
    .A2(_13836_),
    .A3(_13722_),
    .ZN(_13965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22930_ (.A1(_13964_),
    .A2(_13965_),
    .ZN(_13966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22931_ (.A1(_13966_),
    .A2(_13791_),
    .ZN(_13967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22932_ (.A1(_15819_),
    .A2(_15813_),
    .ZN(_13968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22933_ (.A1(_13753_),
    .A2(_13778_),
    .A3(_13968_),
    .ZN(_13969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22934_ (.A1(net872),
    .A2(_15817_),
    .ZN(_13970_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22935_ (.A1(net684),
    .A2(_13970_),
    .A3(_13830_),
    .ZN(_13971_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22936_ (.A1(_13969_),
    .A2(_13769_),
    .A3(_13971_),
    .ZN(_13972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22937_ (.A1(_13967_),
    .A2(_13972_),
    .ZN(_13973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22938_ (.A1(_13973_),
    .A2(_13902_),
    .B(_13748_),
    .ZN(_13974_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22939_ (.A1(_13794_),
    .A2(_13722_),
    .Z(_13975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22940_ (.A1(_15826_),
    .A2(_13803_),
    .ZN(_13976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22941_ (.A1(_13975_),
    .A2(_13976_),
    .ZN(_13977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22942_ (.A1(_13977_),
    .A2(_13866_),
    .A3(_13862_),
    .ZN(_13978_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22943_ (.A1(_13714_),
    .A2(_13826_),
    .A3(_13777_),
    .Z(_13979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22944_ (.A1(_13970_),
    .A2(_13830_),
    .ZN(_13980_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22945_ (.I(_13980_),
    .ZN(_13981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22946_ (.A1(_13979_),
    .A2(_13981_),
    .B(_13863_),
    .ZN(_13982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22947_ (.A1(_13978_),
    .A2(_13982_),
    .A3(_13772_),
    .ZN(_13983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22948_ (.A1(_13974_),
    .A2(_13983_),
    .B(_13822_),
    .ZN(_13984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22949_ (.A1(_13872_),
    .A2(_13791_),
    .ZN(_13985_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22950_ (.A1(_13979_),
    .A2(_13794_),
    .Z(_13986_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22951_ (.A1(_13985_),
    .A2(_13986_),
    .ZN(_13987_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22952_ (.A1(_13721_),
    .A2(_13843_),
    .A3(_13778_),
    .ZN(_13988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22953_ (.A1(_13970_),
    .A2(_13905_),
    .ZN(_13989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22954_ (.A1(_13989_),
    .A2(_13757_),
    .ZN(_13990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22955_ (.A1(_13988_),
    .A2(_13990_),
    .B(_13959_),
    .ZN(_13991_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22956_ (.A1(_13987_),
    .A2(_13991_),
    .B(_13772_),
    .ZN(_13992_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22957_ (.A1(_13753_),
    .A2(_13830_),
    .A3(_13903_),
    .ZN(_13993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22958_ (.I(_13993_),
    .ZN(_13994_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22959_ (.A1(_13714_),
    .A2(_13832_),
    .A3(_13778_),
    .Z(_13995_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22960_ (.A1(_13994_),
    .A2(_13995_),
    .B(_13899_),
    .ZN(_13996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22961_ (.A1(_13711_),
    .A2(_13703_),
    .A3(_13786_),
    .ZN(_13997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22962_ (.A1(_13796_),
    .A2(_13763_),
    .ZN(_13998_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22963_ (.A1(_13997_),
    .A2(_13873_),
    .A3(_13998_),
    .ZN(_13999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22964_ (.A1(_13996_),
    .A2(_13999_),
    .A3(_13902_),
    .ZN(_14000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22965_ (.A1(_13992_),
    .A2(_13749_),
    .A3(_14000_),
    .ZN(_14001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22966_ (.A1(_13984_),
    .A2(_14001_),
    .ZN(_14002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22967_ (.A1(net680),
    .A2(_13722_),
    .ZN(_14003_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22968_ (.A1(_13870_),
    .A2(_13673_),
    .B1(_13676_),
    .B2(_14003_),
    .ZN(_14004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22969_ (.A1(_14004_),
    .A2(_13671_),
    .ZN(_14005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22970_ (.A1(_13719_),
    .A2(_13702_),
    .Z(_14006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22971_ (.A1(_14006_),
    .A2(_13843_),
    .ZN(_14007_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22972_ (.A1(_13778_),
    .A2(_15827_),
    .Z(_14008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22973_ (.A1(_14007_),
    .A2(_13873_),
    .A3(_14008_),
    .ZN(_14009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22974_ (.A1(_14005_),
    .A2(_13772_),
    .A3(_14009_),
    .ZN(_14010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22975_ (.I(_13751_),
    .ZN(_14011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22976_ (.A1(_13845_),
    .A2(_14011_),
    .ZN(_14012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22977_ (.A1(_15824_),
    .A2(_13763_),
    .B(_13907_),
    .ZN(_14013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22978_ (.A1(_14012_),
    .A2(_14013_),
    .B(_13936_),
    .ZN(_14014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22979_ (.A1(_13922_),
    .A2(_13714_),
    .ZN(_14015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22980_ (.A1(_14015_),
    .A2(_13874_),
    .ZN(_14016_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22981_ (.A1(_13872_),
    .A2(_14016_),
    .A3(_13726_),
    .ZN(_14017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22982_ (.A1(_14014_),
    .A2(_14017_),
    .B(_13748_),
    .ZN(_14018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22983_ (.A1(_14010_),
    .A2(_14018_),
    .ZN(_14019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22984_ (.A1(_13753_),
    .A2(_13779_),
    .ZN(_14020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22985_ (.I(_13782_),
    .ZN(_14021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22986_ (.A1(_14021_),
    .A2(_13905_),
    .ZN(_14022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22987_ (.A1(_14020_),
    .A2(_14022_),
    .B(_13703_),
    .ZN(_14023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22988_ (.A1(_14023_),
    .A2(_13671_),
    .A3(_13940_),
    .ZN(_14024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22989_ (.A1(_13762_),
    .A2(_13757_),
    .ZN(_14025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22990_ (.A1(_14025_),
    .A2(_13865_),
    .Z(_14026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22991_ (.A1(_13766_),
    .A2(_13976_),
    .ZN(_14027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22992_ (.A1(_14027_),
    .A2(_14026_),
    .B(_13936_),
    .ZN(_14028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22993_ (.A1(_14024_),
    .A2(_14028_),
    .ZN(_14029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22994_ (.A1(_13896_),
    .A2(_15831_),
    .ZN(_14030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22995_ (.A1(_13988_),
    .A2(_13726_),
    .A3(_14030_),
    .ZN(_14031_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22996_ (.A1(_13830_),
    .A2(_15822_),
    .Z(_14032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22997_ (.A1(_13998_),
    .A2(_13959_),
    .A3(_14032_),
    .ZN(_14033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22998_ (.A1(_14031_),
    .A2(_14033_),
    .A3(_13868_),
    .ZN(_14034_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22999_ (.A1(_13749_),
    .A2(_14034_),
    .A3(_14029_),
    .ZN(_14035_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23000_ (.A1(_14035_),
    .A2(_14019_),
    .A3(_13822_),
    .ZN(_14036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23001_ (.A1(_14036_),
    .A2(_14002_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23002_ (.A1(_13847_),
    .A2(_13709_),
    .Z(_14037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23003_ (.A1(_14037_),
    .A2(_13903_),
    .ZN(_14038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23004_ (.A1(_13898_),
    .A2(_14038_),
    .A3(_13907_),
    .ZN(_14039_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23005_ (.A1(_13719_),
    .A2(_13724_),
    .A3(_13790_),
    .Z(_14040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23006_ (.A1(_13778_),
    .A2(_15819_),
    .ZN(_14041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23007_ (.A1(_14040_),
    .A2(_14041_),
    .ZN(_14042_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23008_ (.A1(_14039_),
    .A2(_13771_),
    .A3(_14042_),
    .Z(_14043_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23009_ (.A1(_14043_),
    .A2(_13749_),
    .ZN(_14044_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23010_ (.A1(_13895_),
    .A2(_13722_),
    .A3(_13837_),
    .Z(_14045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23011_ (.A1(_13753_),
    .A2(_13702_),
    .Z(_14046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23012_ (.A1(_13724_),
    .A2(_13675_),
    .Z(_14047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23013_ (.A1(_14046_),
    .A2(_14047_),
    .ZN(_14048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23014_ (.A1(_14045_),
    .A2(_14048_),
    .A3(_13959_),
    .ZN(_14049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _23015_ (.I(_13710_),
    .ZN(_14050_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23016_ (.A1(_14050_),
    .A2(_13760_),
    .B(_13725_),
    .C(_13769_),
    .ZN(_14051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23017_ (.A1(_14049_),
    .A2(_14051_),
    .ZN(_14052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23018_ (.A1(_14052_),
    .A2(_13902_),
    .ZN(_14053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23019_ (.A1(_14044_),
    .A2(_14053_),
    .ZN(_14054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23020_ (.A1(_13761_),
    .A2(_13750_),
    .ZN(_14055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23021_ (.A1(_14055_),
    .A2(_13874_),
    .ZN(_14056_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23022_ (.A1(_13839_),
    .A2(_14047_),
    .B(_14056_),
    .C(_13726_),
    .ZN(_14057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23023_ (.A1(_13787_),
    .A2(_13976_),
    .ZN(_14058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23024_ (.A1(_14058_),
    .A2(_13993_),
    .A3(_13873_),
    .ZN(_14059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23025_ (.A1(_14057_),
    .A2(_14059_),
    .A3(_13902_),
    .ZN(_14060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23026_ (.A1(_14015_),
    .A2(_13896_),
    .ZN(_14061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23027_ (.A1(_14061_),
    .A2(_13752_),
    .B(_13740_),
    .ZN(_14062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23028_ (.A1(_13716_),
    .A2(_13721_),
    .ZN(_14063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23029_ (.A1(_13766_),
    .A2(_13753_),
    .ZN(_14064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23030_ (.A1(_14063_),
    .A2(_14064_),
    .A3(_13959_),
    .ZN(_14065_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23031_ (.A1(_14065_),
    .A2(_14062_),
    .B(_13881_),
    .ZN(_14066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23032_ (.A1(_14066_),
    .A2(_14060_),
    .B(_13820_),
    .ZN(_14067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23033_ (.A1(_14054_),
    .A2(_14067_),
    .ZN(_14068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23034_ (.A1(_13861_),
    .A2(_13722_),
    .ZN(_14069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23035_ (.A1(_13901_),
    .A2(_14069_),
    .Z(_14070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23036_ (.A1(_14070_),
    .A2(_13964_),
    .B(_13726_),
    .ZN(_14071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23037_ (.A1(_13803_),
    .A2(_13781_),
    .Z(_14072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23038_ (.A1(_14072_),
    .A2(_15819_),
    .ZN(_14073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23039_ (.A1(_13702_),
    .A2(_14073_),
    .Z(_14074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23040_ (.A1(_14074_),
    .A2(_13811_),
    .ZN(_14075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23041_ (.A1(_13801_),
    .A2(_13706_),
    .ZN(_14076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23042_ (.A1(_14075_),
    .A2(_14076_),
    .A3(_13936_),
    .ZN(_14077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23043_ (.A1(_14071_),
    .A2(_14077_),
    .B(_13882_),
    .ZN(_14078_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _23044_ (.A1(_13844_),
    .A2(_13852_),
    .B1(_13830_),
    .B2(_13750_),
    .ZN(_14079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23045_ (.A1(_14079_),
    .A2(_13771_),
    .ZN(_14080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23046_ (.I(_13758_),
    .ZN(_14081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _23047_ (.A1(_14081_),
    .A2(_13901_),
    .B1(_13703_),
    .B2(net1133),
    .ZN(_14082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23048_ (.A1(_14080_),
    .A2(_14082_),
    .ZN(_14083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23049_ (.A1(_14083_),
    .A2(_13671_),
    .ZN(_14084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23050_ (.A1(_14078_),
    .A2(_14084_),
    .ZN(_14085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23051_ (.I(_13811_),
    .ZN(_14086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23052_ (.A1(_13800_),
    .A2(_13861_),
    .B(_13702_),
    .ZN(_14087_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23053_ (.A1(_14050_),
    .A2(_14086_),
    .B(_14087_),
    .C(_13769_),
    .ZN(_14088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23054_ (.A1(_13831_),
    .A2(_13918_),
    .A3(_13873_),
    .ZN(_14089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23055_ (.A1(_14088_),
    .A2(_14089_),
    .A3(_13902_),
    .ZN(_14090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23056_ (.A1(_13847_),
    .A2(_14074_),
    .ZN(_14091_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23057_ (.A1(_13940_),
    .A2(_13959_),
    .A3(_14091_),
    .ZN(_14092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23058_ (.I(_13971_),
    .ZN(_14093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23059_ (.A1(_14093_),
    .A2(_13726_),
    .B(_13901_),
    .ZN(_14094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23060_ (.A1(_14092_),
    .A2(_14094_),
    .B(_13748_),
    .ZN(_14095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23061_ (.A1(_14095_),
    .A2(_14090_),
    .ZN(_14096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23062_ (.A1(_14096_),
    .A2(_14085_),
    .A3(_13820_),
    .ZN(_14097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23063_ (.A1(_14097_),
    .A2(_14068_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _23064_ (.A1(_13671_),
    .A2(_13935_),
    .A3(_13755_),
    .A4(_14025_),
    .ZN(_14098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23065_ (.A1(_13716_),
    .A2(_13811_),
    .B(_13916_),
    .ZN(_14099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23066_ (.A1(_14099_),
    .A2(_13886_),
    .ZN(_14100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23067_ (.A1(_14098_),
    .A2(_14100_),
    .A3(_13772_),
    .ZN(_14101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23068_ (.A1(_13913_),
    .A2(_13836_),
    .ZN(_14102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23069_ (.A1(_13780_),
    .A2(_13886_),
    .A3(_14102_),
    .ZN(_14103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23070_ (.A1(_13947_),
    .A2(_13757_),
    .ZN(_14104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23071_ (.A1(_14104_),
    .A2(_13907_),
    .Z(_14105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23072_ (.A1(_13711_),
    .A2(_13839_),
    .ZN(_14106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23073_ (.A1(_14105_),
    .A2(_14106_),
    .B(_13936_),
    .ZN(_14107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23074_ (.A1(_14103_),
    .A2(_14107_),
    .ZN(_14108_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23075_ (.A1(_14101_),
    .A2(_13882_),
    .A3(_14108_),
    .ZN(_14109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _23076_ (.I(_15815_),
    .ZN(_14110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23077_ (.A1(_13830_),
    .A2(_14110_),
    .ZN(_14111_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _23078_ (.A1(_14003_),
    .A2(_14111_),
    .A3(_13865_),
    .Z(_14112_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23079_ (.A1(_13868_),
    .A2(_14112_),
    .ZN(_14113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23080_ (.A1(_13848_),
    .A2(_13794_),
    .ZN(_14114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23081_ (.A1(_14114_),
    .A2(_13825_),
    .A3(_13899_),
    .ZN(_14115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23082_ (.A1(_14113_),
    .A2(_14115_),
    .B(_13882_),
    .ZN(_14116_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23083_ (.A1(_13721_),
    .A2(net867),
    .A3(_13896_),
    .ZN(_14117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23084_ (.A1(_13848_),
    .A2(net685),
    .ZN(_14118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23085_ (.A1(_14117_),
    .A2(_14118_),
    .A3(_13899_),
    .ZN(_14119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23086_ (.A1(_13878_),
    .A2(_13725_),
    .A3(_13873_),
    .ZN(_14120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23087_ (.A1(_14119_),
    .A2(_14120_),
    .A3(_13868_),
    .ZN(_14121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23088_ (.A1(_14121_),
    .A2(_14116_),
    .B(_13822_),
    .ZN(_14122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23089_ (.A1(_14109_),
    .A2(_14122_),
    .ZN(_14123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23090_ (.A1(_13827_),
    .A2(_13907_),
    .Z(_14124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23091_ (.A1(_13968_),
    .A2(_13953_),
    .Z(_14125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23092_ (.A1(_14125_),
    .A2(_14124_),
    .B(_13936_),
    .ZN(_14126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23093_ (.A1(_13946_),
    .A2(_13750_),
    .ZN(_14127_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23094_ (.A1(_13849_),
    .A2(_13873_),
    .A3(_14127_),
    .ZN(_14128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23095_ (.A1(_14128_),
    .A2(_14126_),
    .B(_13882_),
    .ZN(_14129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23096_ (.A1(_13845_),
    .A2(_13839_),
    .A3(_13753_),
    .ZN(_14130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23097_ (.A1(_13990_),
    .A2(_13907_),
    .Z(_14131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23098_ (.A1(_14130_),
    .A2(_14131_),
    .B(_13740_),
    .ZN(_14132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23099_ (.A1(_13922_),
    .A2(_13761_),
    .ZN(_14133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23100_ (.A1(_14133_),
    .A2(_13839_),
    .ZN(_14134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23101_ (.A1(_13828_),
    .A2(_13886_),
    .A3(_14134_),
    .ZN(_14135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23102_ (.A1(_14132_),
    .A2(_14135_),
    .ZN(_14136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23103_ (.A1(_14136_),
    .A2(_14129_),
    .ZN(_14137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23104_ (.A1(_13975_),
    .A2(_13767_),
    .ZN(_14138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23105_ (.A1(net28),
    .A2(net662),
    .ZN(_14139_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23106_ (.A1(_14139_),
    .A2(_13794_),
    .A3(_13757_),
    .ZN(_14140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23107_ (.A1(_14138_),
    .A2(_13671_),
    .A3(_14140_),
    .ZN(_14141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23108_ (.A1(_14007_),
    .A2(_13873_),
    .A3(_13934_),
    .ZN(_14142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23109_ (.A1(_14141_),
    .A2(_14142_),
    .A3(_13772_),
    .ZN(_14143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23110_ (.A1(_13922_),
    .A2(_13722_),
    .A3(_13808_),
    .ZN(_14144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23111_ (.A1(_13932_),
    .A2(_14144_),
    .A3(_13959_),
    .ZN(_14145_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23112_ (.A1(_14021_),
    .A2(_13670_),
    .Z(_14146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23113_ (.I(_13848_),
    .ZN(_14147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23114_ (.A1(_14146_),
    .A2(_14147_),
    .B(_13771_),
    .ZN(_14148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23115_ (.A1(_14145_),
    .A2(_14148_),
    .B(_13748_),
    .ZN(_14149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23116_ (.A1(_14143_),
    .A2(_14149_),
    .ZN(_14150_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23117_ (.A1(_13822_),
    .A2(_14150_),
    .A3(_14137_),
    .ZN(_14151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23118_ (.A1(_14123_),
    .A2(_14151_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23119_ (.A1(_13702_),
    .A2(_15808_),
    .Z(_14152_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23120_ (.A1(_13856_),
    .A2(_14152_),
    .ZN(_14153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23121_ (.A1(_13845_),
    .A2(_14037_),
    .ZN(_14154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23122_ (.A1(_14153_),
    .A2(_14154_),
    .ZN(_14155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23123_ (.A1(_13989_),
    .A2(_13722_),
    .ZN(_14156_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23124_ (.A1(_13783_),
    .A2(_14156_),
    .A3(_13755_),
    .ZN(_14157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23125_ (.A1(_14155_),
    .A2(_14157_),
    .A3(_13901_),
    .ZN(_14158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23126_ (.A1(_14087_),
    .A2(_14050_),
    .A3(_13791_),
    .ZN(_14159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23127_ (.A1(_13913_),
    .A2(_13790_),
    .ZN(_14160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23128_ (.A1(_13916_),
    .A2(_13721_),
    .ZN(_14161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23129_ (.A1(_14160_),
    .A2(_14161_),
    .ZN(_14162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23130_ (.A1(_14159_),
    .A2(_14162_),
    .A3(_13771_),
    .ZN(_14163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23131_ (.A1(_14163_),
    .A2(_14158_),
    .ZN(_14164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23132_ (.A1(_14164_),
    .A2(_13882_),
    .ZN(_14165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23133_ (.A1(_13722_),
    .A2(net28),
    .ZN(_14166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23134_ (.A1(_14140_),
    .A2(_14166_),
    .ZN(_14167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23135_ (.A1(_14167_),
    .A2(_13791_),
    .ZN(_14168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23136_ (.A1(_13801_),
    .A2(_14139_),
    .B(_13865_),
    .ZN(_14169_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23137_ (.A1(net684),
    .A2(net19),
    .B(_13851_),
    .ZN(_14170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23138_ (.A1(_14170_),
    .A2(_13778_),
    .ZN(_14171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23139_ (.A1(_14169_),
    .A2(_14171_),
    .ZN(_14172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23140_ (.A1(_14168_),
    .A2(_14172_),
    .A3(_13740_),
    .ZN(_14173_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23141_ (.A1(_13844_),
    .A2(_14104_),
    .ZN(_14174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23142_ (.I(_13953_),
    .ZN(_14175_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23143_ (.A1(_14174_),
    .A2(_14175_),
    .B(_13769_),
    .ZN(_14176_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23144_ (.A1(_13673_),
    .A2(_13765_),
    .B(_13980_),
    .C(_13791_),
    .ZN(_14177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23145_ (.A1(_14176_),
    .A2(_14177_),
    .A3(_13868_),
    .ZN(_14178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23146_ (.A1(_14173_),
    .A2(_14178_),
    .A3(_13749_),
    .ZN(_14179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23147_ (.A1(_14179_),
    .A2(_14165_),
    .ZN(_14180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23148_ (.A1(_14180_),
    .A2(_13822_),
    .ZN(_14181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23149_ (.A1(_13776_),
    .A2(_13763_),
    .ZN(_14182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23150_ (.A1(_13760_),
    .A2(_13703_),
    .ZN(_14183_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23151_ (.A1(_14182_),
    .A2(_14086_),
    .B(_13726_),
    .C(_14183_),
    .ZN(_14184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23152_ (.A1(_13775_),
    .A2(_13830_),
    .ZN(_14185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23153_ (.A1(_13780_),
    .A2(_13866_),
    .A3(_14185_),
    .ZN(_14186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23154_ (.A1(_14184_),
    .A2(_14186_),
    .A3(_13772_),
    .ZN(_14187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23155_ (.A1(net667),
    .A2(_13874_),
    .B(_13907_),
    .ZN(_14188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23156_ (.A1(_13720_),
    .A2(_14188_),
    .B(_13936_),
    .ZN(_14189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23157_ (.A1(_13766_),
    .A2(_13796_),
    .ZN(_14190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23158_ (.A1(_14037_),
    .A2(_13794_),
    .ZN(_14191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23159_ (.A1(_14190_),
    .A2(_14191_),
    .A3(_13726_),
    .ZN(_14192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23160_ (.A1(_14189_),
    .A2(_14192_),
    .B(_13748_),
    .ZN(_14193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23161_ (.A1(_14187_),
    .A2(_14193_),
    .ZN(_14194_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23162_ (.I(_13812_),
    .ZN(_14195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23163_ (.A1(_14124_),
    .A2(_14195_),
    .B(_13936_),
    .ZN(_14196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23164_ (.I(_13776_),
    .ZN(_14197_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23165_ (.A1(_14074_),
    .A2(_13769_),
    .ZN(_14198_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23166_ (.A1(_14197_),
    .A2(_13998_),
    .B(_14198_),
    .ZN(_14199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23167_ (.A1(_14196_),
    .A2(_14199_),
    .ZN(_14200_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _23168_ (.I(_13903_),
    .ZN(_14201_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23169_ (.A1(_14201_),
    .A2(_14086_),
    .A3(_13778_),
    .Z(_14202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23170_ (.A1(_13766_),
    .A2(_13851_),
    .ZN(_14203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23171_ (.A1(_14202_),
    .A2(_13899_),
    .A3(_14203_),
    .ZN(_14204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23172_ (.A1(_13674_),
    .A2(_13874_),
    .B(_13907_),
    .ZN(_14205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23173_ (.A1(_14182_),
    .A2(_14205_),
    .B(_13901_),
    .ZN(_14206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23174_ (.A1(_14204_),
    .A2(_14206_),
    .ZN(_14207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23175_ (.A1(_14200_),
    .A2(_14207_),
    .A3(_13749_),
    .ZN(_14208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23176_ (.A1(_14194_),
    .A2(_14208_),
    .A3(_13820_),
    .ZN(_14209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23177_ (.A1(_14181_),
    .A2(_14209_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23178_ (.A1(_14006_),
    .A2(_13946_),
    .B(_13724_),
    .ZN(_14210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23179_ (.A1(_14210_),
    .A2(_13671_),
    .ZN(_14211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23180_ (.A1(_13709_),
    .A2(net19),
    .ZN(_14212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23181_ (.A1(_14040_),
    .A2(_14212_),
    .B(_13936_),
    .ZN(_14213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23182_ (.A1(_14211_),
    .A2(_14213_),
    .ZN(_14214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23183_ (.A1(_14201_),
    .A2(_13763_),
    .ZN(_14215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23184_ (.A1(_14087_),
    .A2(_13959_),
    .A3(_14215_),
    .ZN(_14216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23185_ (.A1(_13810_),
    .A2(_13923_),
    .ZN(_14217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23186_ (.A1(_14216_),
    .A2(_14217_),
    .A3(_13868_),
    .ZN(_14218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23187_ (.A1(_14218_),
    .A2(_14214_),
    .B(_13749_),
    .ZN(_14219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23188_ (.A1(_13979_),
    .A2(_13873_),
    .A3(_13794_),
    .ZN(_14220_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23189_ (.A1(_14114_),
    .A2(_13726_),
    .A3(_13852_),
    .ZN(_14221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23190_ (.A1(_14220_),
    .A2(_14221_),
    .A3(_13868_),
    .ZN(_14222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23191_ (.A1(_13812_),
    .A2(_13903_),
    .ZN(_14223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23192_ (.A1(_13952_),
    .A2(_14223_),
    .ZN(_14224_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23193_ (.I(_15821_),
    .ZN(_14225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23194_ (.A1(_14225_),
    .A2(_13874_),
    .B(_13907_),
    .ZN(_14226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23195_ (.A1(_14191_),
    .A2(_14226_),
    .ZN(_14227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23196_ (.A1(_14224_),
    .A2(_13740_),
    .A3(_14227_),
    .ZN(_14228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23197_ (.A1(_14222_),
    .A2(_14228_),
    .B(_13882_),
    .ZN(_14229_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23198_ (.A1(_14219_),
    .A2(_14229_),
    .B(_13820_),
    .ZN(_14230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23199_ (.A1(_13916_),
    .A2(_14139_),
    .ZN(_14231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23200_ (.A1(_13786_),
    .A2(_13847_),
    .A3(_13757_),
    .ZN(_14232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23201_ (.A1(_14231_),
    .A2(_13855_),
    .A3(_14232_),
    .ZN(_14233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23202_ (.A1(_14233_),
    .A2(_13959_),
    .ZN(_14234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23203_ (.A1(_13968_),
    .A2(_13832_),
    .Z(_14235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23204_ (.A1(_14235_),
    .A2(_13778_),
    .A3(_13826_),
    .ZN(_14236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23205_ (.A1(_14236_),
    .A2(_13838_),
    .A3(_14185_),
    .ZN(_14237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23206_ (.A1(_14234_),
    .A2(_14237_),
    .ZN(_14238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23207_ (.A1(_14238_),
    .A2(_13772_),
    .ZN(_14239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23208_ (.A1(_14046_),
    .A2(_13721_),
    .ZN(_14240_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23209_ (.A1(_15820_),
    .A2(_15829_),
    .Z(_14241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23210_ (.A1(_13763_),
    .A2(_14241_),
    .B(_13907_),
    .ZN(_14242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23211_ (.A1(_14240_),
    .A2(_14242_),
    .B(_13771_),
    .ZN(_14243_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23212_ (.A1(_13896_),
    .A2(_14235_),
    .B(_14025_),
    .C(_13769_),
    .ZN(_14244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23213_ (.A1(_14243_),
    .A2(_14244_),
    .B(_13748_),
    .ZN(_14245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23214_ (.A1(_14239_),
    .A2(_14245_),
    .ZN(_14246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23215_ (.A1(_13916_),
    .A2(net694),
    .B(_13769_),
    .ZN(_14247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23216_ (.A1(_13887_),
    .A2(_14073_),
    .ZN(_14248_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23217_ (.A1(_14247_),
    .A2(_13725_),
    .A3(_14248_),
    .ZN(_14249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23218_ (.A1(_13721_),
    .A2(_13922_),
    .A3(_13874_),
    .ZN(_14250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23219_ (.A1(_13760_),
    .A2(_13763_),
    .B(_13865_),
    .ZN(_14251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23220_ (.A1(_14250_),
    .A2(_14251_),
    .B(_13901_),
    .ZN(_14252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23221_ (.A1(_14249_),
    .A2(_14252_),
    .B(_13881_),
    .ZN(_14253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23222_ (.A1(_13975_),
    .A2(_13796_),
    .ZN(_14254_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23223_ (.A1(_14104_),
    .A2(_14201_),
    .Z(_14255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23224_ (.A1(_14255_),
    .A2(_13873_),
    .A3(_14254_),
    .ZN(_14256_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23225_ (.A1(_13796_),
    .A2(_13896_),
    .A3(net659),
    .ZN(_14257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23226_ (.A1(_14257_),
    .A2(_13899_),
    .A3(_14032_),
    .ZN(_14258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23227_ (.A1(_14256_),
    .A2(_14258_),
    .A3(_13902_),
    .ZN(_14259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23228_ (.A1(_14259_),
    .A2(_14253_),
    .ZN(_14260_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23229_ (.A1(_14260_),
    .A2(_14246_),
    .A3(_13822_),
    .ZN(_14261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23230_ (.A1(_14230_),
    .A2(_14261_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23231_ (.A1(net663),
    .A2(_13839_),
    .B(_14144_),
    .ZN(_14262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23232_ (.A1(_14262_),
    .A2(_13671_),
    .ZN(_14263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23233_ (.A1(_13795_),
    .A2(_13711_),
    .ZN(_14264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23234_ (.A1(_14264_),
    .A2(_14007_),
    .A3(_13886_),
    .ZN(_14265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23235_ (.A1(_14263_),
    .A2(_14265_),
    .A3(_13902_),
    .ZN(_14266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23236_ (.A1(_13845_),
    .A2(_13839_),
    .ZN(_14267_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23237_ (.A1(_13711_),
    .A2(_13896_),
    .A3(_13903_),
    .ZN(_14268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23238_ (.A1(_14267_),
    .A2(_14268_),
    .A3(_13899_),
    .ZN(_14269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23239_ (.A1(_13758_),
    .A2(_13865_),
    .Z(_14270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23240_ (.A1(_13895_),
    .A2(_13703_),
    .ZN(_14271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23241_ (.A1(_14270_),
    .A2(_14271_),
    .B(_13901_),
    .ZN(_14272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23242_ (.A1(_14272_),
    .A2(_14269_),
    .B(_13881_),
    .ZN(_14273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23243_ (.A1(_14266_),
    .A2(_14273_),
    .B(_13822_),
    .ZN(_14274_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23244_ (.A1(_14020_),
    .A2(_13762_),
    .Z(_14275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23245_ (.A1(_14275_),
    .A2(_13839_),
    .ZN(_14276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23246_ (.A1(_13845_),
    .A2(net870),
    .B(_13791_),
    .ZN(_14277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23247_ (.A1(_14276_),
    .A2(_14277_),
    .ZN(_14278_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23248_ (.I(_13946_),
    .ZN(_14279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23249_ (.A1(_14114_),
    .A2(_13886_),
    .A3(_14279_),
    .ZN(_14280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23250_ (.A1(_14278_),
    .A2(_13902_),
    .A3(_14280_),
    .ZN(_14281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23251_ (.A1(_14016_),
    .A2(_13886_),
    .A3(_14232_),
    .ZN(_14282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23252_ (.A1(_13925_),
    .A2(_14076_),
    .A3(_13899_),
    .ZN(_14283_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23253_ (.A1(_14282_),
    .A2(_14283_),
    .A3(_13868_),
    .ZN(_14284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23254_ (.A1(_14281_),
    .A2(_13882_),
    .A3(_14284_),
    .ZN(_14285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23255_ (.A1(_14274_),
    .A2(_14285_),
    .ZN(_14286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23256_ (.A1(_13839_),
    .A2(_14110_),
    .ZN(_14287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23257_ (.A1(_14287_),
    .A2(_13834_),
    .B(_13771_),
    .ZN(_14288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23258_ (.A1(_14212_),
    .A2(_13670_),
    .Z(_14289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23259_ (.A1(_13935_),
    .A2(_14289_),
    .A3(_14185_),
    .ZN(_14290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23260_ (.A1(_14288_),
    .A2(_14290_),
    .B(_13881_),
    .ZN(_14291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23261_ (.A1(_14011_),
    .A2(_13903_),
    .ZN(_14292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23262_ (.A1(_13801_),
    .A2(_13794_),
    .ZN(_14293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23263_ (.A1(_14292_),
    .A2(_14293_),
    .A3(_13899_),
    .ZN(_14294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23264_ (.A1(_13750_),
    .A2(_13968_),
    .Z(_14295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23265_ (.A1(_13874_),
    .A2(_15829_),
    .ZN(_14296_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23266_ (.A1(_14295_),
    .A2(_13839_),
    .B(_13959_),
    .C(_14296_),
    .ZN(_14297_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23267_ (.A1(_14294_),
    .A2(_14297_),
    .A3(_13868_),
    .ZN(_14298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23268_ (.A1(_14298_),
    .A2(_14291_),
    .B(_13820_),
    .ZN(_14299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23269_ (.A1(_14275_),
    .A2(_13896_),
    .ZN(_14300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23270_ (.A1(_13903_),
    .A2(_13851_),
    .A3(_13703_),
    .ZN(_14301_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23271_ (.A1(_14300_),
    .A2(_13886_),
    .A3(_14301_),
    .ZN(_14302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23272_ (.A1(_13800_),
    .A2(_13830_),
    .ZN(_14303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23273_ (.A1(_14289_),
    .A2(_14303_),
    .Z(_14304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _23274_ (.A1(_14091_),
    .A2(_14304_),
    .B(_13936_),
    .ZN(_14305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23275_ (.A1(_14302_),
    .A2(_14305_),
    .ZN(_14306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23276_ (.A1(_13896_),
    .A2(_15808_),
    .ZN(_14307_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23277_ (.A1(_14240_),
    .A2(_13899_),
    .A3(_14307_),
    .ZN(_14308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23278_ (.A1(_13754_),
    .A2(_13703_),
    .ZN(_14309_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23279_ (.A1(_13834_),
    .A2(_13761_),
    .A3(_14309_),
    .ZN(_14310_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23280_ (.A1(_14308_),
    .A2(_14310_),
    .A3(_13868_),
    .ZN(_14311_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23281_ (.A1(_13882_),
    .A2(_14311_),
    .A3(_14306_),
    .ZN(_14312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23282_ (.A1(_14312_),
    .A2(_14299_),
    .ZN(_14313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23283_ (.A1(_14313_),
    .A2(_14286_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _23284_ (.I(\sa21_sr[7] ),
    .ZN(_14314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23285_ (.A1(_14314_),
    .A2(\sa21_sr[0] ),
    .ZN(_14315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23286_ (.A1(_11194_),
    .A2(_11436_),
    .ZN(_14316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23287_ (.A1(_14315_),
    .A2(_14316_),
    .ZN(_14317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23288_ (.A1(_14317_),
    .A2(_11161_),
    .Z(_14318_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23289_ (.A1(_11161_),
    .A2(_14317_),
    .ZN(_14319_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23290_ (.A1(_14318_),
    .A2(_14319_),
    .ZN(_14320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23291_ (.A1(_11174_),
    .A2(_11212_),
    .ZN(_14321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23292_ (.A1(\sa01_sr[1] ),
    .A2(_11170_),
    .ZN(_14322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23293_ (.A1(_14321_),
    .A2(_14322_),
    .Z(_14323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23294_ (.A1(_14320_),
    .A2(_14323_),
    .ZN(_14324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23295_ (.A1(_11194_),
    .A2(_14314_),
    .ZN(_14325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23296_ (.A1(\sa21_sr[0] ),
    .A2(_11436_),
    .ZN(_14326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23297_ (.A1(_14325_),
    .A2(_14326_),
    .ZN(_14327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23298_ (.A1(_11147_),
    .A2(_14327_),
    .ZN(_14328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23299_ (.A1(_11161_),
    .A2(_14317_),
    .ZN(_14329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23300_ (.A1(_14328_),
    .A2(_14329_),
    .ZN(_14330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23301_ (.A1(_14321_),
    .A2(_14322_),
    .ZN(_14331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23302_ (.A1(_14330_),
    .A2(_14331_),
    .ZN(_14332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _23303_ (.I(_10378_),
    .Z(_14333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23304_ (.A1(_14333_),
    .A2(_14332_),
    .A3(_14324_),
    .ZN(_14334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23305_ (.A1(_11203_),
    .A2(\text_in_r[81] ),
    .ZN(_14335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23306_ (.A1(_14335_),
    .A2(_14334_),
    .ZN(_14336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23307_ (.A1(_14336_),
    .A2(_07874_),
    .ZN(_14337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23308_ (.A1(net512),
    .A2(net1031),
    .A3(_14335_),
    .ZN(_14338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23309_ (.A1(_14337_),
    .A2(_14338_),
    .ZN(_15839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23310_ (.A1(_11165_),
    .A2(net516),
    .ZN(_14339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23311_ (.A1(_11190_),
    .A2(_11168_),
    .ZN(_14340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23312_ (.A1(_14339_),
    .A2(_14340_),
    .ZN(_14341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23313_ (.A1(_14341_),
    .A2(net812),
    .ZN(_14342_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23314_ (.A1(_14339_),
    .A2(_14340_),
    .A3(_11149_),
    .ZN(_14343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23315_ (.A1(_14342_),
    .A2(_14343_),
    .A3(net551),
    .ZN(_14344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23316_ (.A1(\sa01_sr[0] ),
    .A2(_11168_),
    .ZN(_14345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23317_ (.I(_14345_),
    .ZN(_14346_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23318_ (.A1(net798),
    .A2(net43),
    .ZN(_14347_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23319_ (.A1(_14346_),
    .A2(_14347_),
    .B(net517),
    .ZN(_14348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23320_ (.A1(_11149_),
    .A2(_11165_),
    .ZN(_14349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23321_ (.A1(_14349_),
    .A2(_11190_),
    .A3(_14345_),
    .ZN(_14350_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23322_ (.A1(_14327_),
    .A2(_14348_),
    .A3(_14350_),
    .ZN(_14351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _23323_ (.A1(_14344_),
    .A2(net521),
    .B(_10410_),
    .ZN(_14352_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23324_ (.I(\text_in_r[80] ),
    .ZN(_14353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23325_ (.A1(_14353_),
    .A2(_10431_),
    .Z(_14354_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23326_ (.A1(_14352_),
    .A2(_14354_),
    .B(\u0.w[1][16] ),
    .ZN(_14355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23327_ (.A1(_14351_),
    .A2(_14344_),
    .ZN(_14356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23328_ (.A1(_11989_),
    .A2(_14356_),
    .ZN(_14357_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23329_ (.I(_14354_),
    .ZN(_14358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23330_ (.A1(_14357_),
    .A2(_07869_),
    .A3(_14358_),
    .ZN(_14359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23331_ (.A1(_14355_),
    .A2(_14359_),
    .ZN(_15842_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23332_ (.A1(_11218_),
    .A2(\sa30_sub[2] ),
    .Z(_14360_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23333_ (.A1(_11218_),
    .A2(\sa30_sub[2] ),
    .ZN(_14361_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23334_ (.A1(_14360_),
    .A2(_14361_),
    .B(\sa01_sr[2] ),
    .ZN(_14362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23335_ (.A1(_11216_),
    .A2(_11221_),
    .ZN(_14363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23336_ (.A1(_11218_),
    .A2(\sa30_sub[2] ),
    .ZN(_14364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23337_ (.A1(_14363_),
    .A2(_11250_),
    .A3(_14364_),
    .ZN(_14365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23338_ (.A1(_14362_),
    .A2(_14365_),
    .ZN(_14366_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23339_ (.A1(net808),
    .A2(\sa21_sr[1] ),
    .ZN(_14367_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23340_ (.I(_14367_),
    .ZN(_14368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23341_ (.A1(_14366_),
    .A2(_14368_),
    .ZN(_14369_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23342_ (.A1(_14362_),
    .A2(_14365_),
    .A3(_14367_),
    .ZN(_14370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _23343_ (.A1(_14369_),
    .A2(_14370_),
    .B(_10482_),
    .ZN(_14371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23344_ (.I(\text_in_r[82] ),
    .ZN(_14372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23345_ (.A1(_14372_),
    .A2(_11202_),
    .Z(_14373_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23346_ (.A1(_14371_),
    .A2(_14373_),
    .B(_07879_),
    .ZN(_14374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23347_ (.A1(_14369_),
    .A2(_14370_),
    .ZN(_14375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23348_ (.A1(_14375_),
    .A2(_14333_),
    .ZN(_14376_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23349_ (.I(_14373_),
    .ZN(_14377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23350_ (.A1(_14376_),
    .A2(\u0.w[1][18] ),
    .A3(_14377_),
    .ZN(_14378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23351_ (.A1(_14374_),
    .A2(_14378_),
    .ZN(_14379_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23352_ (.I(_14379_),
    .Z(_15858_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23353_ (.A1(_14354_),
    .A2(_14352_),
    .B(_07869_),
    .ZN(_14380_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23354_ (.A1(_14358_),
    .A2(\u0.w[1][16] ),
    .A3(_14357_),
    .ZN(_14381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23355_ (.A1(_14380_),
    .A2(_14381_),
    .ZN(_15833_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23356_ (.A1(_14371_),
    .A2(_14373_),
    .B(\u0.w[1][18] ),
    .ZN(_14382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23357_ (.A1(_14376_),
    .A2(_07879_),
    .A3(_14377_),
    .ZN(_14383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23358_ (.A1(_14383_),
    .A2(_14382_),
    .ZN(_14384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _23359_ (.I(_14384_),
    .Z(_15851_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _23360_ (.I(_14379_),
    .Z(_14385_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _23361_ (.I(_15836_),
    .ZN(_14386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23362_ (.A1(_14385_),
    .A2(_14386_),
    .ZN(_14387_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23363_ (.I(_14387_),
    .ZN(_14388_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23364_ (.A1(_11218_),
    .A2(_11436_),
    .Z(_14389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23365_ (.A1(_14389_),
    .A2(_11262_),
    .ZN(_14390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23366_ (.A1(_11216_),
    .A2(_14314_),
    .ZN(_14391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23367_ (.A1(_11218_),
    .A2(net26),
    .ZN(_14392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23368_ (.A1(_14391_),
    .A2(_14392_),
    .ZN(_14393_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23369_ (.A1(_11249_),
    .A2(_14393_),
    .ZN(_14394_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23370_ (.A1(_14390_),
    .A2(_14394_),
    .ZN(_14395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23371_ (.A1(_11165_),
    .A2(_11223_),
    .ZN(_14396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23372_ (.A1(net523),
    .A2(\sa11_sr[2] ),
    .ZN(_14397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23373_ (.A1(_14396_),
    .A2(_14397_),
    .ZN(_14398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23374_ (.A1(_14398_),
    .A2(\sa01_sr[3] ),
    .ZN(_14399_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23375_ (.I(\sa01_sr[3] ),
    .ZN(_14400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23376_ (.A1(_14396_),
    .A2(_14400_),
    .A3(_14397_),
    .ZN(_14401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23377_ (.A1(_14399_),
    .A2(_14401_),
    .ZN(_14402_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23378_ (.I(_14402_),
    .ZN(_14403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23379_ (.A1(_14395_),
    .A2(_14403_),
    .ZN(_14404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23380_ (.A1(_11249_),
    .A2(_14393_),
    .ZN(_14405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23381_ (.A1(_14389_),
    .A2(_11262_),
    .ZN(_14406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23382_ (.A1(_14405_),
    .A2(_14406_),
    .ZN(_14407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23383_ (.A1(_14407_),
    .A2(_14402_),
    .ZN(_14408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23384_ (.A1(_14404_),
    .A2(_14408_),
    .A3(_14333_),
    .ZN(_14409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23385_ (.A1(_11203_),
    .A2(\text_in_r[83] ),
    .ZN(_14410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23386_ (.A1(_14409_),
    .A2(_14410_),
    .ZN(_14411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23387_ (.A1(_14411_),
    .A2(_07884_),
    .ZN(_14412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23388_ (.A1(_14409_),
    .A2(\u0.w[1][19] ),
    .A3(_14410_),
    .ZN(_14413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23389_ (.A1(_14412_),
    .A2(_14413_),
    .ZN(_14414_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23390_ (.I(_14414_),
    .Z(_14415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23391_ (.A1(_14388_),
    .A2(_14415_),
    .ZN(_14416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23392_ (.A1(_11258_),
    .A2(_14314_),
    .ZN(_14417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23393_ (.A1(\sa21_sr[3] ),
    .A2(_11436_),
    .ZN(_14418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23394_ (.A1(_14417_),
    .A2(_14418_),
    .ZN(_14419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23395_ (.A1(_11305_),
    .A2(_14419_),
    .ZN(_14420_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23396_ (.I(_14419_),
    .ZN(_14421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23397_ (.A1(_14421_),
    .A2(_11304_),
    .ZN(_14422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23398_ (.A1(_14420_),
    .A2(_14422_),
    .ZN(_14423_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23399_ (.A1(_11273_),
    .A2(\sa01_sr[4] ),
    .Z(_14424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23400_ (.A1(_11273_),
    .A2(\sa01_sr[4] ),
    .ZN(_14425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23401_ (.A1(_14424_),
    .A2(_14425_),
    .ZN(_14426_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23402_ (.A1(_14423_),
    .A2(_14426_),
    .Z(_14427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23403_ (.A1(_14423_),
    .A2(_14426_),
    .ZN(_14428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23404_ (.A1(_14427_),
    .A2(_11989_),
    .A3(_14428_),
    .ZN(_14429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23405_ (.A1(_10586_),
    .A2(\text_in_r[84] ),
    .ZN(_14430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23406_ (.A1(_14429_),
    .A2(_14430_),
    .ZN(_14431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23407_ (.A1(_14431_),
    .A2(\u0.w[1][20] ),
    .ZN(_14432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23408_ (.A1(_14429_),
    .A2(_07888_),
    .A3(_14430_),
    .ZN(_14433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23409_ (.A1(_14432_),
    .A2(_14433_),
    .ZN(_14434_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _23410_ (.I(_14434_),
    .ZN(_14435_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23411_ (.I(_14435_),
    .Z(_14436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23412_ (.A1(_14416_),
    .A2(_14436_),
    .Z(_14437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23413_ (.A1(_14374_),
    .A2(_14386_),
    .A3(_14378_),
    .ZN(_14438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23414_ (.A1(_14411_),
    .A2(\u0.w[1][19] ),
    .ZN(_14439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23415_ (.A1(_14409_),
    .A2(_07884_),
    .A3(_14410_),
    .ZN(_14440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23416_ (.A1(_14439_),
    .A2(_14440_),
    .ZN(_14441_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23417_ (.I(_14441_),
    .Z(_14442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23418_ (.A1(_14438_),
    .A2(_14442_),
    .Z(_14443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23419_ (.A1(_14336_),
    .A2(net1031),
    .ZN(_14444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23420_ (.A1(_14334_),
    .A2(_07874_),
    .A3(_14335_),
    .ZN(_14445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23421_ (.A1(_14444_),
    .A2(_14445_),
    .ZN(_15834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23422_ (.A1(net504),
    .A2(_14385_),
    .ZN(_14446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23423_ (.A1(_14443_),
    .A2(_14446_),
    .ZN(_14447_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23424_ (.A1(\sa01_sr[5] ),
    .A2(_11339_),
    .ZN(_14448_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23425_ (.A1(\sa11_sr[4] ),
    .A2(\sa21_sr[4] ),
    .ZN(_14449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23426_ (.I(_14449_),
    .ZN(_14450_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23427_ (.A1(_14448_),
    .A2(_14450_),
    .Z(_14451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23428_ (.A1(_14448_),
    .A2(_14450_),
    .ZN(_14452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23429_ (.A1(_14451_),
    .A2(_14452_),
    .A3(_10403_),
    .ZN(_14453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23430_ (.A1(_12115_),
    .A2(\text_in_r[85] ),
    .ZN(_14454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23431_ (.A1(_14453_),
    .A2(_14454_),
    .ZN(_14455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23432_ (.A1(_14455_),
    .A2(\u0.w[1][21] ),
    .ZN(_14456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23433_ (.A1(_14453_),
    .A2(_07893_),
    .A3(_14454_),
    .ZN(_14457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23434_ (.A1(_14456_),
    .A2(_14457_),
    .ZN(_14458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23435_ (.I(_14458_),
    .ZN(_14459_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23436_ (.I(_14459_),
    .Z(_14460_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23437_ (.A1(_14437_),
    .A2(_14447_),
    .B(_14460_),
    .ZN(_14461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23438_ (.I(_15835_),
    .ZN(_14462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23439_ (.A1(_14384_),
    .A2(_14462_),
    .ZN(_14463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23440_ (.I(_14463_),
    .ZN(_14464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23441_ (.A1(_14464_),
    .A2(_14442_),
    .ZN(_14465_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23442_ (.I(_14434_),
    .Z(_14466_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23443_ (.A1(_14465_),
    .A2(_14466_),
    .Z(_14467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23444_ (.A1(net950),
    .A2(_14438_),
    .ZN(_14468_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _23445_ (.I(_14468_),
    .ZN(_14469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23446_ (.A1(_15858_),
    .A2(_15835_),
    .ZN(_14470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23447_ (.A1(_14469_),
    .A2(_14470_),
    .ZN(_14471_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23448_ (.I(_15843_),
    .ZN(_14472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23449_ (.A1(_15858_),
    .A2(_14472_),
    .Z(_14473_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23450_ (.I(_14442_),
    .Z(_14474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23451_ (.A1(_14473_),
    .A2(_14474_),
    .ZN(_14475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23452_ (.A1(_14467_),
    .A2(_14471_),
    .A3(_14475_),
    .ZN(_14476_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23453_ (.A1(\sa11_sr[5] ),
    .A2(\sa21_sr[5] ),
    .ZN(_14477_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23454_ (.I(\sa01_sr[6] ),
    .ZN(_14478_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23455_ (.A1(_14478_),
    .A2(_11382_),
    .Z(_14479_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23456_ (.A1(_14477_),
    .A2(_14479_),
    .ZN(_14480_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23457_ (.A1(_11203_),
    .A2(\text_in_r[86] ),
    .Z(_14481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23458_ (.A1(_14480_),
    .A2(_10523_),
    .B(_14481_),
    .ZN(_14482_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23459_ (.A1(\u0.w[1][22] ),
    .A2(_14482_),
    .Z(_14483_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23460_ (.I(_14483_),
    .Z(_14484_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _23461_ (.I(_14484_),
    .ZN(_14485_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23462_ (.I(_14485_),
    .Z(_14486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23463_ (.A1(_14461_),
    .A2(_14476_),
    .B(_14486_),
    .ZN(_14487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23464_ (.A1(_14384_),
    .A2(_15842_),
    .ZN(_14488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23465_ (.A1(_14488_),
    .A2(_14441_),
    .ZN(_14489_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _23466_ (.I(_14489_),
    .ZN(_14490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23467_ (.A1(net2),
    .A2(net522),
    .ZN(_14491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23468_ (.A1(_14490_),
    .A2(_14491_),
    .ZN(_14492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23469_ (.A1(net552),
    .A2(_15833_),
    .ZN(_14493_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23470_ (.I(_14414_),
    .Z(_14494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23471_ (.A1(_14385_),
    .A2(_15842_),
    .ZN(_14495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23472_ (.A1(_14493_),
    .A2(_14494_),
    .A3(_14495_),
    .ZN(_14496_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23473_ (.I(_14436_),
    .Z(_14497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23474_ (.A1(_14492_),
    .A2(_14496_),
    .A3(_14497_),
    .ZN(_14498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23475_ (.A1(net14),
    .A2(_15842_),
    .A3(_15858_),
    .ZN(_14499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23476_ (.A1(_14499_),
    .A2(_14443_),
    .ZN(_14500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23477_ (.A1(_15858_),
    .A2(_14462_),
    .ZN(_14501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23478_ (.A1(_15851_),
    .A2(_14472_),
    .ZN(_14502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23479_ (.A1(_14501_),
    .A2(_14502_),
    .ZN(_14503_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23480_ (.I(_14415_),
    .Z(_14504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23481_ (.A1(_14503_),
    .A2(_14504_),
    .ZN(_14505_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23482_ (.I(_14466_),
    .Z(_14506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23483_ (.A1(_14500_),
    .A2(_14505_),
    .A3(_14506_),
    .ZN(_14507_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23484_ (.I(_14459_),
    .Z(_14508_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23485_ (.I(_14508_),
    .Z(_14509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23486_ (.A1(_14498_),
    .A2(_14507_),
    .A3(_14509_),
    .ZN(_14510_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23487_ (.A1(net35),
    .A2(\sa11_sr[6] ),
    .Z(_14511_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23488_ (.A1(\sa21_sr[6] ),
    .A2(_14511_),
    .Z(_14512_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _23489_ (.A1(net26),
    .A2(net819),
    .A3(_14512_),
    .Z(_14513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _23490_ (.I0(_14513_),
    .I1(\text_in_r[87] ),
    .S(_10639_),
    .Z(_14514_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23491_ (.A1(_07904_),
    .A2(_14514_),
    .Z(_14515_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23492_ (.I(_14515_),
    .Z(_14516_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _23493_ (.I(_14516_),
    .ZN(_14517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23494_ (.A1(_14487_),
    .A2(_14510_),
    .B(_14517_),
    .ZN(_14518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23495_ (.A1(_14384_),
    .A2(net503),
    .ZN(_14519_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23496_ (.I(_14519_),
    .ZN(_14520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23497_ (.A1(_14385_),
    .A2(net513),
    .ZN(_14521_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23498_ (.I(_14441_),
    .Z(_14522_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23499_ (.A1(_14521_),
    .A2(net2),
    .B(_14522_),
    .ZN(_14523_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23500_ (.I(_15849_),
    .ZN(_14524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23501_ (.A1(_14384_),
    .A2(_14524_),
    .ZN(_14525_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23502_ (.I(net951),
    .Z(_14526_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23503_ (.A1(_14521_),
    .A2(_14525_),
    .A3(_14526_),
    .ZN(_14527_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23504_ (.I(_14435_),
    .Z(_14528_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23505_ (.A1(_14520_),
    .A2(_14523_),
    .B(_14527_),
    .C(_14528_),
    .ZN(_14529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23506_ (.I(_14488_),
    .ZN(_14530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23507_ (.A1(_14530_),
    .A2(net14),
    .ZN(_14531_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23508_ (.I(net949),
    .Z(_14532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23509_ (.A1(_14531_),
    .A2(_14532_),
    .A3(_14521_),
    .ZN(_14533_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23510_ (.I(_14446_),
    .ZN(_14534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _23511_ (.I(_15837_),
    .ZN(_14535_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23512_ (.A1(_14385_),
    .A2(_14535_),
    .ZN(_14536_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23513_ (.I(_14522_),
    .Z(_14537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23514_ (.A1(_14534_),
    .A2(_14536_),
    .B(_14537_),
    .ZN(_14538_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23515_ (.A1(_14533_),
    .A2(_14538_),
    .A3(_14506_),
    .ZN(_14539_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23516_ (.I(_14458_),
    .Z(_14540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23517_ (.A1(_14529_),
    .A2(_14539_),
    .A3(_14540_),
    .ZN(_14541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23518_ (.A1(_14521_),
    .A2(net2),
    .ZN(_14542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _23519_ (.I(_15840_),
    .ZN(_14543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23520_ (.A1(_14384_),
    .A2(_14543_),
    .ZN(_14544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23521_ (.A1(_14544_),
    .A2(_14415_),
    .ZN(_14545_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23522_ (.A1(_14542_),
    .A2(_14545_),
    .ZN(_14546_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23523_ (.I(_14435_),
    .Z(_14547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23524_ (.A1(_14521_),
    .A2(_14522_),
    .ZN(_14548_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _23525_ (.I(_14548_),
    .ZN(_14549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23526_ (.A1(_14546_),
    .A2(_14547_),
    .A3(_14549_),
    .Z(_14550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23527_ (.A1(_14524_),
    .A2(_14385_),
    .ZN(_14551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23528_ (.A1(_14551_),
    .A2(net951),
    .ZN(_14552_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23529_ (.I(_14552_),
    .ZN(_14553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23530_ (.A1(_14553_),
    .A2(_14438_),
    .ZN(_14554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23531_ (.A1(_14384_),
    .A2(_15833_),
    .ZN(_14555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23532_ (.A1(_14493_),
    .A2(_14537_),
    .A3(_14555_),
    .ZN(_14556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23533_ (.A1(_14554_),
    .A2(_14556_),
    .A3(_14528_),
    .ZN(_14557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23534_ (.A1(_14550_),
    .A2(_14509_),
    .A3(_14557_),
    .ZN(_14558_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23535_ (.A1(_14541_),
    .A2(_14558_),
    .A3(_14486_),
    .ZN(_14559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23536_ (.A1(_14518_),
    .A2(_14559_),
    .ZN(_14560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23537_ (.A1(net552),
    .A2(_14384_),
    .ZN(_14561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23538_ (.A1(_14561_),
    .A2(_14522_),
    .Z(_14562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23539_ (.A1(_14382_),
    .A2(net508),
    .A3(_14383_),
    .ZN(_14563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23540_ (.A1(_14562_),
    .A2(_14563_),
    .ZN(_14564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23541_ (.A1(_14385_),
    .A2(_15843_),
    .ZN(_14565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23542_ (.A1(_14565_),
    .A2(_14494_),
    .Z(_14566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23543_ (.A1(_14566_),
    .A2(_14555_),
    .ZN(_14567_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23544_ (.I(_14435_),
    .Z(_14568_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23545_ (.A1(_14564_),
    .A2(_14567_),
    .B(_14568_),
    .ZN(_14569_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23546_ (.I(_14536_),
    .ZN(_14570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23547_ (.A1(_14570_),
    .A2(_14501_),
    .ZN(_14571_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23548_ (.I(_14442_),
    .Z(_14572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23549_ (.A1(_14571_),
    .A2(_14572_),
    .ZN(_14573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23550_ (.I(_14434_),
    .Z(_14574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23551_ (.A1(_14573_),
    .A2(_14545_),
    .B(_14574_),
    .ZN(_14575_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23552_ (.A1(_14569_),
    .A2(_14575_),
    .B(_14486_),
    .ZN(_14576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23553_ (.A1(_14536_),
    .A2(_14415_),
    .ZN(_14577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23554_ (.A1(_14577_),
    .A2(_14436_),
    .Z(_14578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23555_ (.A1(_14565_),
    .A2(_14522_),
    .ZN(_14579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23556_ (.I(_14579_),
    .ZN(_14580_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23557_ (.A1(_14379_),
    .A2(_15842_),
    .ZN(_14581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23558_ (.A1(_14581_),
    .A2(net14),
    .ZN(_14582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23559_ (.A1(_14580_),
    .A2(_14582_),
    .ZN(_14583_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23560_ (.I(_14485_),
    .Z(_14584_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23561_ (.A1(_14578_),
    .A2(_14583_),
    .B(_14584_),
    .ZN(_14585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23562_ (.I(_15845_),
    .ZN(_14586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23563_ (.A1(_14385_),
    .A2(_14586_),
    .ZN(_14587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23564_ (.A1(_14587_),
    .A2(net951),
    .ZN(_14588_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _23565_ (.I(_14588_),
    .ZN(_14589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23566_ (.A1(_14589_),
    .A2(_14582_),
    .ZN(_14590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23567_ (.A1(_14536_),
    .A2(_14572_),
    .ZN(_14591_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23568_ (.A1(_14590_),
    .A2(_14574_),
    .A3(_14591_),
    .ZN(_14592_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23569_ (.I(_14458_),
    .Z(_14593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23570_ (.A1(_14585_),
    .A2(_14592_),
    .B(_14593_),
    .ZN(_14594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23571_ (.A1(_14576_),
    .A2(_14594_),
    .ZN(_14595_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23572_ (.A1(_15851_),
    .A2(_14543_),
    .ZN(_14596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23573_ (.A1(_14537_),
    .A2(_14596_),
    .B(_14436_),
    .ZN(_14597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23574_ (.A1(_14533_),
    .A2(_14597_),
    .ZN(_14598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23575_ (.A1(_15858_),
    .A2(net919),
    .ZN(_14599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23576_ (.A1(_14384_),
    .A2(_15845_),
    .ZN(_14600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23577_ (.A1(_14599_),
    .A2(_14600_),
    .ZN(_14601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23578_ (.A1(_14601_),
    .A2(_14537_),
    .ZN(_14602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23579_ (.A1(_14602_),
    .A2(_14468_),
    .A3(_14568_),
    .ZN(_14603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23580_ (.A1(_14598_),
    .A2(_14603_),
    .A3(_14584_),
    .ZN(_14604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23581_ (.A1(_14495_),
    .A2(_14463_),
    .ZN(_14605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23582_ (.A1(_14605_),
    .A2(_14526_),
    .B(_14436_),
    .ZN(_14606_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23583_ (.I(_14441_),
    .Z(_14607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23584_ (.A1(_14385_),
    .A2(_14543_),
    .ZN(_14608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23585_ (.A1(_14582_),
    .A2(_14607_),
    .A3(_14608_),
    .ZN(_14609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23586_ (.A1(_14385_),
    .A2(_15837_),
    .ZN(_14610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23587_ (.I(_14610_),
    .ZN(_14611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23588_ (.A1(_14611_),
    .A2(_14442_),
    .Z(_14612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23589_ (.I(_14612_),
    .ZN(_14613_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23590_ (.A1(_14606_),
    .A2(_14609_),
    .A3(_14613_),
    .ZN(_14614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23591_ (.A1(_14504_),
    .A2(_15856_),
    .ZN(_14615_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23592_ (.I(_14563_),
    .ZN(_14616_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23593_ (.I(_14522_),
    .Z(_14617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _23594_ (.A1(_14616_),
    .A2(_14617_),
    .B(_14434_),
    .ZN(_14618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23595_ (.A1(_14615_),
    .A2(_14618_),
    .B(_14485_),
    .ZN(_14619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23596_ (.A1(_14614_),
    .A2(_14619_),
    .ZN(_14620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23597_ (.A1(_14604_),
    .A2(_14620_),
    .A3(_14540_),
    .ZN(_14621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23598_ (.A1(_14595_),
    .A2(_14621_),
    .A3(_14517_),
    .ZN(_14622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23599_ (.A1(_14560_),
    .A2(_14622_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23600_ (.A1(_14552_),
    .A2(_14520_),
    .B(_14436_),
    .ZN(_14623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23601_ (.A1(_14519_),
    .A2(_14555_),
    .ZN(_14624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23602_ (.A1(_14624_),
    .A2(_14607_),
    .Z(_14625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23603_ (.A1(_14623_),
    .A2(_14625_),
    .ZN(_14626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23604_ (.A1(_14446_),
    .A2(_14521_),
    .A3(_14438_),
    .ZN(_14627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23605_ (.A1(_15851_),
    .A2(net919),
    .ZN(_14628_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23606_ (.A1(_14628_),
    .A2(_14532_),
    .B(_14434_),
    .ZN(_14629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23607_ (.A1(_14627_),
    .A2(_14504_),
    .B(_14629_),
    .ZN(_14630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23608_ (.A1(_14626_),
    .A2(_14630_),
    .B(_14460_),
    .ZN(_14631_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23609_ (.A1(_14495_),
    .A2(_14463_),
    .A3(_14617_),
    .ZN(_14632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23610_ (.A1(_14599_),
    .A2(net510),
    .A3(_14532_),
    .ZN(_14633_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23611_ (.I(_14434_),
    .Z(_14634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23612_ (.A1(_14632_),
    .A2(_14633_),
    .B(_14634_),
    .ZN(_14635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23613_ (.A1(_14563_),
    .A2(_14442_),
    .ZN(_14636_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23614_ (.A1(_14636_),
    .A2(_14581_),
    .B(_14466_),
    .ZN(_14637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23615_ (.A1(_15842_),
    .A2(net511),
    .ZN(_14638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23616_ (.A1(_14638_),
    .A2(_14555_),
    .B(_14607_),
    .ZN(_14639_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23617_ (.A1(_14637_),
    .A2(_14639_),
    .ZN(_14640_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23618_ (.A1(_14635_),
    .A2(_14640_),
    .B(_14593_),
    .ZN(_14641_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23619_ (.A1(_14631_),
    .A2(_14486_),
    .A3(_14641_),
    .ZN(_14642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23620_ (.A1(_15851_),
    .A2(_15849_),
    .ZN(_14643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23621_ (.A1(_14643_),
    .A2(_14563_),
    .ZN(_14644_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23622_ (.A1(_14644_),
    .A2(_14494_),
    .B(_14435_),
    .ZN(_14645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23623_ (.A1(_14645_),
    .A2(_14609_),
    .ZN(_14646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _23624_ (.A1(_14596_),
    .A2(_14442_),
    .B(_14434_),
    .ZN(_14647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23625_ (.A1(net14),
    .A2(_15858_),
    .ZN(_14648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23626_ (.A1(_14648_),
    .A2(net951),
    .ZN(_14649_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23627_ (.A1(_14647_),
    .A2(net509),
    .A3(_14649_),
    .ZN(_14650_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23628_ (.A1(_14646_),
    .A2(_14650_),
    .A3(_14458_),
    .ZN(_14651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23629_ (.A1(_14469_),
    .A2(_14521_),
    .ZN(_14652_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23630_ (.A1(_14495_),
    .A2(_14544_),
    .A3(_14607_),
    .ZN(_14653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23631_ (.I(_14435_),
    .Z(_14654_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23632_ (.A1(_14652_),
    .A2(_14653_),
    .A3(_14654_),
    .ZN(_14655_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23633_ (.A1(_14441_),
    .A2(_15851_),
    .ZN(_14656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23634_ (.A1(_14656_),
    .A2(_14493_),
    .B(_14435_),
    .ZN(_14657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23635_ (.A1(_14561_),
    .A2(_14491_),
    .A3(_14607_),
    .ZN(_14658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23636_ (.A1(_14657_),
    .A2(_14658_),
    .ZN(_14659_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23637_ (.A1(_14655_),
    .A2(_14659_),
    .A3(_14508_),
    .ZN(_14660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23638_ (.A1(_14660_),
    .A2(_14651_),
    .ZN(_14661_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23639_ (.I(_14484_),
    .Z(_14662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23640_ (.A1(_14661_),
    .A2(_14662_),
    .ZN(_14663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23641_ (.A1(_14663_),
    .A2(_14642_),
    .ZN(_14664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23642_ (.A1(_14664_),
    .A2(_14517_),
    .ZN(_14665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23643_ (.A1(_14495_),
    .A2(net952),
    .ZN(_14666_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23644_ (.A1(_14563_),
    .A2(_14607_),
    .ZN(_14667_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23645_ (.A1(_14666_),
    .A2(_14667_),
    .ZN(_14668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23646_ (.A1(_14536_),
    .A2(_14537_),
    .B(_14634_),
    .ZN(_14669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23647_ (.A1(_14464_),
    .A2(_14494_),
    .ZN(_14670_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23648_ (.A1(_14668_),
    .A2(_14669_),
    .A3(_14670_),
    .ZN(_14671_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23649_ (.A1(_14446_),
    .A2(_14532_),
    .A3(_14544_),
    .ZN(_14672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23650_ (.A1(_14488_),
    .A2(_14470_),
    .A3(_14537_),
    .ZN(_14673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23651_ (.A1(_14672_),
    .A2(_14673_),
    .A3(_14574_),
    .ZN(_14674_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23652_ (.A1(_14671_),
    .A2(_14674_),
    .A3(_14460_),
    .ZN(_14675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23653_ (.A1(_14531_),
    .A2(_14549_),
    .ZN(_14676_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23654_ (.A1(_14468_),
    .A2(_14466_),
    .Z(_14677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23655_ (.A1(_14676_),
    .A2(_14677_),
    .B(_14508_),
    .ZN(_14678_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23656_ (.A1(_14525_),
    .A2(_14442_),
    .Z(_14679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23657_ (.A1(_15858_),
    .A2(_14535_),
    .ZN(_14680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23658_ (.A1(_14679_),
    .A2(_14680_),
    .B(_14634_),
    .ZN(_14681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23659_ (.A1(_14627_),
    .A2(_14504_),
    .ZN(_14682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23660_ (.A1(_14681_),
    .A2(_14682_),
    .ZN(_14683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23661_ (.A1(_14678_),
    .A2(_14683_),
    .ZN(_14684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23662_ (.A1(_14675_),
    .A2(_14684_),
    .B(_14662_),
    .ZN(_14685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23663_ (.A1(_14490_),
    .A2(_14648_),
    .ZN(_14686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23664_ (.A1(_14686_),
    .A2(_14672_),
    .ZN(_14687_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23665_ (.A1(_14687_),
    .A2(_14593_),
    .B(_14506_),
    .ZN(_14688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23666_ (.A1(_14495_),
    .A2(net14),
    .ZN(_14689_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _23667_ (.I(_14415_),
    .Z(_14690_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23668_ (.A1(_14689_),
    .A2(_14581_),
    .B(_14690_),
    .ZN(_14691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23669_ (.A1(_14555_),
    .A2(_14470_),
    .A3(_14617_),
    .ZN(_14692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23670_ (.A1(_14691_),
    .A2(_14692_),
    .ZN(_14693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23671_ (.A1(_14693_),
    .A2(_14460_),
    .ZN(_14694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23672_ (.I(_15859_),
    .ZN(_14695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23673_ (.A1(_14415_),
    .A2(_14695_),
    .Z(_14696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23674_ (.A1(_14696_),
    .A2(_14458_),
    .B(_14654_),
    .ZN(_14697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23675_ (.A1(_14531_),
    .A2(_14580_),
    .ZN(_14698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23676_ (.A1(_14697_),
    .A2(_14698_),
    .ZN(_14699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23677_ (.A1(_14699_),
    .A2(_14484_),
    .ZN(_14700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23678_ (.A1(_14688_),
    .A2(_14694_),
    .B(_14700_),
    .ZN(_14701_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23679_ (.A1(_14685_),
    .A2(_14701_),
    .B(_14516_),
    .ZN(_14702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23680_ (.A1(_14665_),
    .A2(_14702_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23681_ (.A1(_14525_),
    .A2(net950),
    .Z(_14703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23682_ (.A1(_14703_),
    .A2(_14499_),
    .ZN(_14704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23683_ (.A1(_14704_),
    .A2(_14523_),
    .ZN(_14705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23684_ (.A1(_14705_),
    .A2(_14574_),
    .ZN(_14706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23685_ (.A1(_15851_),
    .A2(net507),
    .ZN(_14707_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23686_ (.A1(_14446_),
    .A2(_14607_),
    .A3(_14707_),
    .ZN(_14708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23687_ (.A1(_14488_),
    .A2(_14610_),
    .A3(_14532_),
    .ZN(_14709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23688_ (.A1(_14708_),
    .A2(_14709_),
    .A3(_14547_),
    .ZN(_14710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23689_ (.A1(_14706_),
    .A2(_14460_),
    .A3(_14710_),
    .ZN(_14711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23690_ (.A1(_14689_),
    .A2(_14494_),
    .ZN(_14712_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23691_ (.A1(_14544_),
    .A2(_14551_),
    .A3(_14607_),
    .ZN(_14713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23692_ (.A1(_14712_),
    .A2(_14713_),
    .ZN(_14714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23693_ (.A1(_14714_),
    .A2(_14547_),
    .B(_14508_),
    .ZN(_14715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23694_ (.A1(_14582_),
    .A2(_14608_),
    .ZN(_14716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23695_ (.A1(_14716_),
    .A2(_14532_),
    .ZN(_14717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23696_ (.A1(_14717_),
    .A2(_14564_),
    .A3(_14634_),
    .ZN(_14718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23697_ (.A1(_14715_),
    .A2(_14718_),
    .ZN(_14719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23698_ (.A1(_14711_),
    .A2(_14719_),
    .ZN(_14720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23699_ (.A1(_14720_),
    .A2(_14662_),
    .ZN(_14721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23700_ (.A1(_15858_),
    .A2(_15849_),
    .ZN(_14722_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23701_ (.I(_14722_),
    .ZN(_14723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23702_ (.A1(_14489_),
    .A2(_14723_),
    .B(_14654_),
    .ZN(_14724_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23703_ (.A1(_14446_),
    .A2(_14532_),
    .A3(_14600_),
    .Z(_14725_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23704_ (.A1(_14724_),
    .A2(_14725_),
    .ZN(_14726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23705_ (.A1(_14563_),
    .A2(_14415_),
    .Z(_14727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23706_ (.A1(_14727_),
    .A2(_14438_),
    .ZN(_14728_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23707_ (.A1(_14555_),
    .A2(_14587_),
    .A3(_14617_),
    .ZN(_14729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23708_ (.A1(_14728_),
    .A2(_14729_),
    .B(_14568_),
    .ZN(_14730_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23709_ (.A1(_14726_),
    .A2(_14730_),
    .B(_14509_),
    .ZN(_14731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23710_ (.A1(net509),
    .A2(_14690_),
    .A3(_14608_),
    .ZN(_14732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23711_ (.A1(_14732_),
    .A2(_14602_),
    .A3(_14574_),
    .ZN(_14733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23712_ (.A1(_14488_),
    .A2(_14532_),
    .ZN(_14734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23713_ (.A1(_14722_),
    .A2(_14607_),
    .ZN(_14735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23714_ (.A1(_14734_),
    .A2(_14596_),
    .B(_14735_),
    .ZN(_14736_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23715_ (.I(_14600_),
    .ZN(_14737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23716_ (.A1(_14737_),
    .A2(_14607_),
    .ZN(_14738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23717_ (.A1(_14738_),
    .A2(_14436_),
    .Z(_14739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23718_ (.A1(_14736_),
    .A2(_14739_),
    .ZN(_14740_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23719_ (.A1(_14733_),
    .A2(_14740_),
    .A3(_14593_),
    .ZN(_14741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23720_ (.A1(_14731_),
    .A2(_14741_),
    .A3(_14486_),
    .ZN(_14742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23721_ (.A1(_14721_),
    .A2(_14742_),
    .A3(_14516_),
    .ZN(_14743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23722_ (.A1(_14446_),
    .A2(_14415_),
    .Z(_14744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23723_ (.A1(_14744_),
    .A2(_14555_),
    .ZN(_14745_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _23724_ (.I(_14458_),
    .Z(_14746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23725_ (.A1(_14564_),
    .A2(_14745_),
    .B(_14746_),
    .ZN(_14747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23726_ (.A1(_14727_),
    .A2(_14502_),
    .B(_14508_),
    .ZN(_14748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23727_ (.A1(_14562_),
    .A2(_14501_),
    .ZN(_14749_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23728_ (.A1(_14748_),
    .A2(_14749_),
    .Z(_14750_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23729_ (.A1(_14747_),
    .A2(_14750_),
    .B(_14497_),
    .ZN(_14751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23730_ (.A1(_15856_),
    .A2(_14572_),
    .B(_14458_),
    .ZN(_14752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23731_ (.A1(_14387_),
    .A2(_14415_),
    .Z(_14753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23732_ (.A1(_14753_),
    .A2(_14582_),
    .ZN(_14754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23733_ (.A1(_14752_),
    .A2(_14754_),
    .B(_14568_),
    .ZN(_14755_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23734_ (.A1(_14561_),
    .A2(_14491_),
    .A3(_14494_),
    .ZN(_14756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23735_ (.A1(_14474_),
    .A2(_14695_),
    .ZN(_14757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23736_ (.A1(_14756_),
    .A2(_14593_),
    .A3(_14757_),
    .ZN(_14758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23737_ (.A1(_14755_),
    .A2(_14758_),
    .B(_14662_),
    .ZN(_14759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23738_ (.A1(_14751_),
    .A2(_14759_),
    .ZN(_14760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23739_ (.A1(_14656_),
    .A2(_14638_),
    .ZN(_14761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23740_ (.A1(_14761_),
    .A2(_14654_),
    .Z(_14762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23741_ (.A1(_14494_),
    .A2(_15851_),
    .ZN(_14763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23742_ (.A1(_14535_),
    .A2(_14543_),
    .Z(_14764_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23743_ (.A1(_14763_),
    .A2(_14764_),
    .Z(_14765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23744_ (.A1(_14762_),
    .A2(_14698_),
    .A3(_14765_),
    .ZN(_14766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23745_ (.A1(_14469_),
    .A2(_14608_),
    .ZN(_14767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23746_ (.A1(_14467_),
    .A2(_14767_),
    .B(_14746_),
    .ZN(_14768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23747_ (.A1(_14768_),
    .A2(_14766_),
    .ZN(_14769_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23748_ (.A1(_14522_),
    .A2(_15854_),
    .Z(_14770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23749_ (.A1(_14523_),
    .A2(_14770_),
    .ZN(_14771_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23750_ (.A1(_14771_),
    .A2(_14547_),
    .Z(_14772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23751_ (.A1(_15863_),
    .A2(_14537_),
    .B(_14466_),
    .ZN(_14773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23752_ (.A1(_14773_),
    .A2(_14712_),
    .B(_14508_),
    .ZN(_14774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23753_ (.A1(_14772_),
    .A2(_14774_),
    .ZN(_14775_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23754_ (.A1(_14769_),
    .A2(_14662_),
    .A3(_14775_),
    .ZN(_14776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23755_ (.A1(_14776_),
    .A2(_14760_),
    .A3(_14517_),
    .ZN(_14777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23756_ (.A1(_14743_),
    .A2(_14777_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23757_ (.A1(_14624_),
    .A2(_14636_),
    .Z(_14778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23758_ (.A1(_14495_),
    .A2(_14502_),
    .Z(_14779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23759_ (.A1(_14744_),
    .A2(_14779_),
    .ZN(_14780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23760_ (.A1(_14778_),
    .A2(_14780_),
    .A3(_14574_),
    .ZN(_14781_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _23761_ (.I(_14438_),
    .ZN(_14782_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23762_ (.A1(_14473_),
    .A2(_14494_),
    .A3(_14782_),
    .Z(_14783_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23763_ (.A1(_14783_),
    .A2(_14568_),
    .A3(_14496_),
    .ZN(_14784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23764_ (.A1(_14781_),
    .A2(_14784_),
    .ZN(_14785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23765_ (.A1(_14785_),
    .A2(_14509_),
    .ZN(_14786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23766_ (.A1(_14493_),
    .A2(_14488_),
    .ZN(_14787_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23767_ (.A1(_14787_),
    .A2(_14466_),
    .Z(_14788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23768_ (.A1(_14788_),
    .A2(_14763_),
    .B(_14460_),
    .ZN(_14789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23769_ (.A1(_14587_),
    .A2(_14522_),
    .Z(_14790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23770_ (.A1(_14790_),
    .A2(_14707_),
    .Z(_14791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23771_ (.A1(_14623_),
    .A2(_14791_),
    .Z(_14792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23772_ (.A1(_14789_),
    .A2(_14792_),
    .B(_14662_),
    .ZN(_14793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23773_ (.A1(_14786_),
    .A2(_14793_),
    .ZN(_14794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23774_ (.A1(_14779_),
    .A2(_14617_),
    .ZN(_14795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23775_ (.A1(_14387_),
    .A2(_14463_),
    .A3(_14532_),
    .ZN(_14796_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23776_ (.A1(_14795_),
    .A2(_14508_),
    .A3(_14796_),
    .ZN(_14797_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23777_ (.A1(_14686_),
    .A2(_14458_),
    .A3(_14416_),
    .ZN(_14798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23778_ (.A1(_14797_),
    .A2(_14798_),
    .ZN(_14799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23779_ (.A1(_14799_),
    .A2(_14497_),
    .ZN(_14800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23780_ (.A1(_14490_),
    .A2(_14493_),
    .ZN(_14801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23781_ (.A1(_14469_),
    .A2(_14446_),
    .ZN(_14802_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23782_ (.A1(_14801_),
    .A2(_14802_),
    .A3(_14593_),
    .ZN(_14803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23783_ (.A1(_14703_),
    .A2(_14608_),
    .ZN(_14804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23784_ (.A1(_14804_),
    .A2(_14708_),
    .A3(_14460_),
    .ZN(_14805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23785_ (.A1(_14506_),
    .A2(_14805_),
    .A3(_14803_),
    .ZN(_14806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23786_ (.A1(_14800_),
    .A2(_14806_),
    .A3(_14662_),
    .ZN(_14807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23787_ (.A1(_14794_),
    .A2(_14807_),
    .A3(_14517_),
    .ZN(_14808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23788_ (.A1(_14737_),
    .A2(_14690_),
    .B(_14458_),
    .ZN(_14809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23789_ (.A1(_14809_),
    .A2(_14729_),
    .B(_14568_),
    .ZN(_14810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23790_ (.A1(_14549_),
    .A2(_14438_),
    .ZN(_14811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23791_ (.A1(_15851_),
    .A2(_14764_),
    .ZN(_14812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23792_ (.A1(_14812_),
    .A2(_14415_),
    .Z(_14813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23793_ (.A1(_14813_),
    .A2(net514),
    .ZN(_14814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23794_ (.A1(_14811_),
    .A2(_14814_),
    .A3(_14746_),
    .ZN(_14815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23795_ (.A1(_14810_),
    .A2(_14815_),
    .B(_14584_),
    .ZN(_14816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23796_ (.A1(_14782_),
    .A2(_14442_),
    .ZN(_14817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23797_ (.I(_14817_),
    .ZN(_14818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _23798_ (.A1(_14818_),
    .A2(_14508_),
    .B1(_14690_),
    .B2(_14536_),
    .ZN(_14819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23799_ (.I(_14561_),
    .ZN(_14820_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23800_ (.A1(_14820_),
    .A2(_14579_),
    .B(_14416_),
    .ZN(_14821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23801_ (.A1(_14821_),
    .A2(_14458_),
    .ZN(_14822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23802_ (.A1(_14819_),
    .A2(_14822_),
    .ZN(_14823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23803_ (.A1(_14823_),
    .A2(_14497_),
    .ZN(_14824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23804_ (.A1(_14816_),
    .A2(_14824_),
    .B(_14517_),
    .ZN(_14825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23805_ (.A1(_14813_),
    .A2(_14587_),
    .ZN(_14826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23806_ (.A1(_14698_),
    .A2(_14826_),
    .B(_14568_),
    .ZN(_14827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23807_ (.I(_14724_),
    .ZN(_14828_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23808_ (.A1(_14827_),
    .A2(_14828_),
    .B(_14540_),
    .ZN(_14829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23809_ (.A1(_14606_),
    .A2(_14658_),
    .ZN(_14830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23810_ (.A1(_14443_),
    .A2(net514),
    .ZN(_14831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23811_ (.A1(_14521_),
    .A2(_14600_),
    .ZN(_14832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23812_ (.A1(_14832_),
    .A2(_14526_),
    .ZN(_14833_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23813_ (.A1(_14831_),
    .A2(_14833_),
    .A3(_14528_),
    .ZN(_14834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23814_ (.A1(_14830_),
    .A2(_14834_),
    .A3(_14509_),
    .ZN(_14835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23815_ (.A1(_14829_),
    .A2(_14835_),
    .A3(_14486_),
    .ZN(_14836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23816_ (.A1(_14825_),
    .A2(_14836_),
    .ZN(_14837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23817_ (.A1(_14808_),
    .A2(_14837_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23818_ (.A1(_14533_),
    .A2(_14506_),
    .ZN(_14838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23819_ (.A1(_14544_),
    .A2(_14537_),
    .ZN(_14839_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23820_ (.A1(_14839_),
    .A2(_14616_),
    .ZN(_14840_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23821_ (.A1(_14680_),
    .A2(_14442_),
    .ZN(_14841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23822_ (.A1(_14841_),
    .A2(_14436_),
    .Z(_14842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23823_ (.A1(_14499_),
    .A2(_14690_),
    .ZN(_14843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23824_ (.A1(_14842_),
    .A2(_14843_),
    .B(_14746_),
    .ZN(_14844_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23825_ (.A1(_14838_),
    .A2(_14840_),
    .B(_14844_),
    .ZN(_14845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23826_ (.A1(_14490_),
    .A2(net514),
    .ZN(_14846_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23827_ (.A1(_14656_),
    .A2(_14547_),
    .ZN(_14847_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23828_ (.A1(_14846_),
    .A2(_14847_),
    .B(_14460_),
    .ZN(_14848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23829_ (.A1(_14446_),
    .A2(_14463_),
    .ZN(_14849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23830_ (.A1(_14849_),
    .A2(_14474_),
    .ZN(_14850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23831_ (.A1(_14850_),
    .A2(_14672_),
    .A3(_14497_),
    .ZN(_14851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23832_ (.A1(_14848_),
    .A2(_14851_),
    .ZN(_14852_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23833_ (.A1(_14845_),
    .A2(_14852_),
    .A3(_14486_),
    .ZN(_14853_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23834_ (.I(_15847_),
    .ZN(_14854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23835_ (.A1(_14854_),
    .A2(_14572_),
    .B(_14654_),
    .ZN(_14855_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23836_ (.I(_14727_),
    .ZN(_14856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23837_ (.A1(_14855_),
    .A2(_14856_),
    .B(_14746_),
    .ZN(_14857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23838_ (.A1(_14589_),
    .A2(net509),
    .ZN(_14858_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23839_ (.A1(_14493_),
    .A2(_15851_),
    .A3(_14617_),
    .ZN(_14859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23840_ (.A1(_14858_),
    .A2(_14859_),
    .A3(_14528_),
    .ZN(_14860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23841_ (.A1(_14857_),
    .A2(_14860_),
    .B(_14584_),
    .ZN(_14861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23842_ (.A1(_14519_),
    .A2(_14638_),
    .ZN(_14862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23843_ (.A1(_14862_),
    .A2(_14617_),
    .ZN(_14863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23844_ (.A1(_14589_),
    .A2(_14488_),
    .ZN(_14864_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23845_ (.A1(_14863_),
    .A2(_14864_),
    .A3(_14497_),
    .ZN(_14865_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23846_ (.A1(_14573_),
    .A2(_14506_),
    .A3(_14496_),
    .ZN(_14866_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23847_ (.A1(_14865_),
    .A2(_14866_),
    .A3(_14540_),
    .ZN(_14867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23848_ (.A1(_14861_),
    .A2(_14867_),
    .ZN(_14868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23849_ (.A1(_14853_),
    .A2(_14516_),
    .A3(_14868_),
    .ZN(_14869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23850_ (.A1(_14756_),
    .A2(_14634_),
    .Z(_14870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23851_ (.A1(_14870_),
    .A2(_14686_),
    .ZN(_14871_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23852_ (.A1(_14862_),
    .A2(_14532_),
    .Z(_14872_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23853_ (.A1(net509),
    .A2(_14504_),
    .A3(_14470_),
    .ZN(_14873_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23854_ (.A1(_14872_),
    .A2(_14873_),
    .A3(_14497_),
    .ZN(_14874_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23855_ (.A1(_14871_),
    .A2(_14874_),
    .A3(_14540_),
    .ZN(_14875_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23856_ (.A1(_14649_),
    .A2(_14581_),
    .Z(_14876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23857_ (.A1(_14876_),
    .A2(_14506_),
    .A3(_14692_),
    .ZN(_14877_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23858_ (.A1(_14570_),
    .A2(_14436_),
    .Z(_14878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23859_ (.A1(_14878_),
    .A2(_14588_),
    .B(_14746_),
    .ZN(_14879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23860_ (.A1(_14877_),
    .A2(_14879_),
    .B(_14484_),
    .ZN(_14880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23861_ (.A1(_14875_),
    .A2(_14880_),
    .ZN(_14881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23862_ (.A1(_14582_),
    .A2(_14526_),
    .ZN(_14882_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23863_ (.A1(_14882_),
    .A2(_14534_),
    .B(_14713_),
    .C(_14568_),
    .ZN(_14883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23864_ (.A1(_14670_),
    .A2(_14466_),
    .Z(_14884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23865_ (.A1(_14656_),
    .A2(net14),
    .ZN(_14885_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23866_ (.A1(_14884_),
    .A2(_14609_),
    .A3(_14885_),
    .ZN(_14886_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23867_ (.A1(_14883_),
    .A2(_14886_),
    .A3(_14540_),
    .ZN(_14887_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23868_ (.A1(_14667_),
    .A2(_14737_),
    .ZN(_14888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23869_ (.A1(_14647_),
    .A2(_14888_),
    .B(_14746_),
    .ZN(_14889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23870_ (.A1(_14644_),
    .A2(_14572_),
    .ZN(_14890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23871_ (.A1(_14590_),
    .A2(_14574_),
    .A3(_14890_),
    .ZN(_14891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23872_ (.A1(_14889_),
    .A2(_14891_),
    .B(_14584_),
    .ZN(_14892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23873_ (.A1(_14887_),
    .A2(_14892_),
    .ZN(_14893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23874_ (.A1(_14881_),
    .A2(_14893_),
    .A3(_14517_),
    .ZN(_14894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23875_ (.A1(_14869_),
    .A2(_14894_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23876_ (.A1(_14531_),
    .A2(_14565_),
    .ZN(_14895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23877_ (.A1(_14895_),
    .A2(_14526_),
    .ZN(_14896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23878_ (.A1(_14549_),
    .A2(_14638_),
    .ZN(_14897_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23879_ (.A1(_14896_),
    .A2(_14568_),
    .A3(_14897_),
    .Z(_14898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23880_ (.A1(_14526_),
    .A2(net2),
    .ZN(_14899_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23881_ (.A1(_14863_),
    .A2(_14634_),
    .A3(_14899_),
    .Z(_14900_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23882_ (.A1(_14898_),
    .A2(_14900_),
    .B(_14509_),
    .ZN(_14901_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23883_ (.A1(_14841_),
    .A2(_14820_),
    .ZN(_14902_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23884_ (.A1(_14902_),
    .A2(_14667_),
    .B(_14547_),
    .ZN(_14903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23885_ (.A1(_14469_),
    .A2(_14501_),
    .ZN(_14904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23886_ (.A1(_14904_),
    .A2(_14634_),
    .A3(_14735_),
    .ZN(_14905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23887_ (.A1(_14905_),
    .A2(_14903_),
    .ZN(_14906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23888_ (.A1(_14906_),
    .A2(_14540_),
    .B(_14486_),
    .ZN(_14907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23889_ (.A1(_14907_),
    .A2(_14901_),
    .ZN(_14908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23890_ (.A1(_14553_),
    .A2(_14544_),
    .ZN(_14909_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23891_ (.A1(_14538_),
    .A2(_14506_),
    .A3(_14909_),
    .ZN(_14910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23892_ (.A1(_14790_),
    .A2(_14582_),
    .ZN(_14911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23893_ (.A1(_14504_),
    .A2(net920),
    .ZN(_14912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23894_ (.A1(_14578_),
    .A2(_14911_),
    .A3(_14912_),
    .ZN(_14913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23895_ (.A1(_14910_),
    .A2(_14913_),
    .A3(_14509_),
    .ZN(_14914_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23896_ (.A1(_14443_),
    .A2(_14547_),
    .ZN(_14915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23897_ (.A1(_14915_),
    .A2(_14833_),
    .B(_14508_),
    .ZN(_14916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23898_ (.A1(_14656_),
    .A2(_14493_),
    .ZN(_14917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23899_ (.A1(_14917_),
    .A2(_14528_),
    .A3(_14839_),
    .ZN(_14918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23900_ (.A1(_14916_),
    .A2(_14918_),
    .B(_14484_),
    .ZN(_14919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23901_ (.A1(_14914_),
    .A2(_14919_),
    .B(_14516_),
    .ZN(_14920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23902_ (.A1(_14908_),
    .A2(_14920_),
    .ZN(_14921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23903_ (.A1(_14530_),
    .A2(_14617_),
    .ZN(_14922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23904_ (.I(_14922_),
    .ZN(_14923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23905_ (.A1(_14531_),
    .A2(_14572_),
    .A3(net515),
    .ZN(_14924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23906_ (.A1(_14473_),
    .A2(_14526_),
    .B(_14634_),
    .ZN(_14925_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23907_ (.A1(_14924_),
    .A2(_14925_),
    .B(_14460_),
    .ZN(_14926_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23908_ (.A1(_14598_),
    .A2(_14923_),
    .B(_14926_),
    .ZN(_14927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23909_ (.A1(_15842_),
    .A2(_14690_),
    .B(_14654_),
    .ZN(_14928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23910_ (.A1(_14928_),
    .A2(_14492_),
    .B(_14746_),
    .ZN(_14929_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23911_ (.A1(_14542_),
    .A2(_14468_),
    .Z(_14930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23912_ (.A1(_14790_),
    .A2(_14519_),
    .ZN(_14931_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23913_ (.A1(_14930_),
    .A2(_14931_),
    .A3(_14528_),
    .ZN(_14932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23914_ (.A1(_14929_),
    .A2(_14932_),
    .B(_14484_),
    .ZN(_14933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23915_ (.A1(_14927_),
    .A2(_14933_),
    .ZN(_14934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23916_ (.A1(_14469_),
    .A2(_14565_),
    .ZN(_14935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23917_ (.A1(net515),
    .A2(_14707_),
    .A3(_14537_),
    .ZN(_14936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23918_ (.A1(_14935_),
    .A2(_14936_),
    .A3(_14528_),
    .ZN(_14937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23919_ (.A1(_14472_),
    .A2(_14690_),
    .B(_14654_),
    .ZN(_14938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23920_ (.A1(_14531_),
    .A2(_14474_),
    .ZN(_14939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23921_ (.A1(_14938_),
    .A2(_14939_),
    .ZN(_14940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23922_ (.A1(_14937_),
    .A2(_14940_),
    .A3(_14593_),
    .ZN(_14941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23923_ (.A1(_14647_),
    .A2(_14552_),
    .B(_14746_),
    .ZN(_14942_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23924_ (.A1(_14689_),
    .A2(_14581_),
    .B(_14572_),
    .ZN(_14943_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23925_ (.A1(_14813_),
    .A2(_14654_),
    .ZN(_14944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23926_ (.A1(_14943_),
    .A2(_14944_),
    .ZN(_14945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23927_ (.A1(_14942_),
    .A2(_14945_),
    .ZN(_14946_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23928_ (.A1(_14941_),
    .A2(_14662_),
    .A3(_14946_),
    .ZN(_14947_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23929_ (.A1(_14934_),
    .A2(_14516_),
    .A3(_14947_),
    .ZN(_14948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23930_ (.A1(_14921_),
    .A2(_14948_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23931_ (.A1(_14790_),
    .A2(_14525_),
    .ZN(_14949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23932_ (.A1(_14949_),
    .A2(_14577_),
    .A3(_14761_),
    .ZN(_14950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23933_ (.A1(_14950_),
    .A2(_14574_),
    .ZN(_14951_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _23934_ (.A1(_14526_),
    .A2(_14599_),
    .A3(_14610_),
    .A4(_14600_),
    .ZN(_14952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23935_ (.A1(_14952_),
    .A2(_14618_),
    .A3(_14922_),
    .ZN(_14953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23936_ (.A1(_14951_),
    .A2(_14953_),
    .ZN(_14954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23937_ (.A1(_14954_),
    .A2(_14540_),
    .ZN(_14955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23938_ (.A1(_14862_),
    .A2(_14690_),
    .ZN(_14956_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23939_ (.A1(_15852_),
    .A2(_15861_),
    .Z(_14957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23940_ (.A1(_14572_),
    .A2(_14957_),
    .B(_14654_),
    .ZN(_14958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23941_ (.A1(_14956_),
    .A2(_14958_),
    .B(_14746_),
    .ZN(_14959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23942_ (.A1(_14610_),
    .A2(_14600_),
    .Z(_14960_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23943_ (.A1(_14474_),
    .A2(_14960_),
    .B(_14465_),
    .C(_14568_),
    .ZN(_14961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23944_ (.A1(_14959_),
    .A2(_14961_),
    .B(_14662_),
    .ZN(_14962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23945_ (.A1(_14955_),
    .A2(_14962_),
    .ZN(_14963_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23946_ (.A1(_14771_),
    .A2(_14547_),
    .A3(_14817_),
    .ZN(_14964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23947_ (.A1(_14519_),
    .A2(_14494_),
    .ZN(_14965_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23948_ (.A1(_14965_),
    .A2(_14542_),
    .B(_14841_),
    .ZN(_14966_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23949_ (.I(_14707_),
    .ZN(_14967_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23950_ (.A1(_14967_),
    .A2(_14617_),
    .B(_14435_),
    .ZN(_14968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23951_ (.A1(_14966_),
    .A2(_14968_),
    .ZN(_14969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23952_ (.A1(_14964_),
    .A2(_14969_),
    .ZN(_14970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23953_ (.A1(_14970_),
    .A2(_14509_),
    .ZN(_14971_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23954_ (.A1(_14582_),
    .A2(_14690_),
    .A3(_14495_),
    .ZN(_14972_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23955_ (.A1(_14812_),
    .A2(_14563_),
    .A3(_14572_),
    .ZN(_14973_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23956_ (.A1(_14972_),
    .A2(_14506_),
    .A3(_14973_),
    .ZN(_14974_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23957_ (.A1(_14530_),
    .A2(net2),
    .B(_14526_),
    .ZN(_14975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23958_ (.A1(_14473_),
    .A2(_14537_),
    .B(_14466_),
    .ZN(_14976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23959_ (.A1(_14975_),
    .A2(_14976_),
    .B(_14508_),
    .ZN(_14977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23960_ (.A1(_14974_),
    .A2(_14977_),
    .B(_14584_),
    .ZN(_14978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23961_ (.A1(_14971_),
    .A2(_14978_),
    .ZN(_14979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23962_ (.A1(_14963_),
    .A2(_14517_),
    .A3(_14979_),
    .ZN(_14980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23963_ (.A1(_14717_),
    .A2(_14634_),
    .ZN(_14981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23964_ (.A1(_14588_),
    .A2(_14520_),
    .B(_14579_),
    .ZN(_14982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23965_ (.A1(_14982_),
    .A2(_14547_),
    .ZN(_14983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23966_ (.A1(_14981_),
    .A2(_14983_),
    .ZN(_14984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23967_ (.A1(_14984_),
    .A2(_14540_),
    .ZN(_14985_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23968_ (.A1(_14617_),
    .A2(_15853_),
    .Z(_14986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23969_ (.A1(_14931_),
    .A2(_14574_),
    .A3(_14986_),
    .ZN(_14987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23970_ (.I(_14666_),
    .ZN(_14988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23971_ (.A1(_14988_),
    .A2(_14436_),
    .Z(_14989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23972_ (.A1(_14553_),
    .A2(_14707_),
    .ZN(_14990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23973_ (.A1(_14989_),
    .A2(_14990_),
    .ZN(_14991_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23974_ (.A1(_14987_),
    .A2(_14991_),
    .A3(_14509_),
    .ZN(_14992_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23975_ (.A1(_14985_),
    .A2(_14992_),
    .A3(_14662_),
    .ZN(_14993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23976_ (.A1(_14787_),
    .A2(_14504_),
    .ZN(_14994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23977_ (.A1(_14521_),
    .A2(_14643_),
    .ZN(_14995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23978_ (.A1(_14995_),
    .A2(_14474_),
    .ZN(_14996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23979_ (.A1(_14994_),
    .A2(_14996_),
    .A3(_14528_),
    .ZN(_14997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23980_ (.A1(_14522_),
    .A2(net2),
    .ZN(_14998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23981_ (.A1(_14788_),
    .A2(_14998_),
    .ZN(_14999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23982_ (.A1(_14997_),
    .A2(_14999_),
    .A3(_14509_),
    .ZN(_15000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23983_ (.A1(_14556_),
    .A2(_14528_),
    .A3(_14649_),
    .ZN(_15001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23984_ (.A1(_14968_),
    .A2(_14833_),
    .ZN(_15002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23985_ (.A1(_15001_),
    .A2(_15002_),
    .A3(_14593_),
    .ZN(_15003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23986_ (.A1(_15000_),
    .A2(_15003_),
    .A3(_14486_),
    .ZN(_15004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23987_ (.A1(_14993_),
    .A2(_15004_),
    .A3(_14516_),
    .ZN(_15005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23988_ (.A1(_14980_),
    .A2(_15005_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23989_ (.A1(_14522_),
    .A2(_15833_),
    .Z(_15006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23990_ (.I(_15006_),
    .ZN(_15007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23991_ (.A1(_14876_),
    .A2(_15007_),
    .ZN(_15008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23992_ (.A1(_15008_),
    .A2(_14497_),
    .B(_14584_),
    .ZN(_15009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23993_ (.A1(_14820_),
    .A2(_14474_),
    .ZN(_15010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23994_ (.A1(_14870_),
    .A2(_14872_),
    .A3(_15010_),
    .ZN(_15011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23995_ (.A1(_15009_),
    .A2(_15011_),
    .ZN(_15012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23996_ (.A1(_14446_),
    .A2(_14463_),
    .A3(_14521_),
    .ZN(_15013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23997_ (.A1(_15013_),
    .A2(_14504_),
    .ZN(_15014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23998_ (.A1(_15014_),
    .A2(_14989_),
    .A3(_14859_),
    .ZN(_15015_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23999_ (.A1(_14679_),
    .A2(_14547_),
    .ZN(_15016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24000_ (.A1(_15016_),
    .A2(_14858_),
    .B(_14484_),
    .ZN(_15017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24001_ (.A1(_15015_),
    .A2(_15017_),
    .B(_14593_),
    .ZN(_15018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24002_ (.A1(_15012_),
    .A2(_15018_),
    .ZN(_15019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24003_ (.A1(_14745_),
    .A2(_14949_),
    .B(_14528_),
    .ZN(_15020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24004_ (.A1(_14644_),
    .A2(_14504_),
    .ZN(_15021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24005_ (.A1(_14811_),
    .A2(_15021_),
    .B(_14574_),
    .ZN(_15022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24006_ (.A1(_15020_),
    .A2(_15022_),
    .B(_14486_),
    .ZN(_15023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24007_ (.A1(_14627_),
    .A2(_14474_),
    .ZN(_15024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24008_ (.A1(_15024_),
    .A2(_14497_),
    .A3(_14882_),
    .ZN(_15025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24009_ (.A1(_14817_),
    .A2(_14466_),
    .Z(_15026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24010_ (.A1(_14624_),
    .A2(_14690_),
    .ZN(_15027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24011_ (.A1(_15026_),
    .A2(_15027_),
    .B(_14584_),
    .ZN(_15028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24012_ (.A1(_15025_),
    .A2(_15028_),
    .B(_14460_),
    .ZN(_15029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24013_ (.A1(_15023_),
    .A2(_15029_),
    .ZN(_15030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24014_ (.A1(_15019_),
    .A2(_14516_),
    .A3(_15030_),
    .ZN(_15031_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24015_ (.A1(_14854_),
    .A2(_14526_),
    .B(_14654_),
    .ZN(_15032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24016_ (.A1(_15032_),
    .A2(_14613_),
    .B(_14584_),
    .ZN(_15033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24017_ (.A1(_14998_),
    .A2(_14435_),
    .Z(_15034_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24018_ (.A1(_14672_),
    .A2(_15034_),
    .A3(_14922_),
    .ZN(_15035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24019_ (.A1(_15033_),
    .A2(_15035_),
    .B(_14593_),
    .ZN(_15036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24020_ (.A1(_15006_),
    .A2(_15858_),
    .ZN(_15037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24021_ (.A1(_15034_),
    .A2(_15037_),
    .Z(_15038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24022_ (.A1(_15038_),
    .A2(_14826_),
    .B(_14484_),
    .ZN(_15039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24023_ (.A1(_15013_),
    .A2(_14474_),
    .ZN(_15040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24024_ (.A1(_14566_),
    .A2(_14707_),
    .ZN(_15041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24025_ (.A1(_15040_),
    .A2(_14506_),
    .A3(_15041_),
    .ZN(_15042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24026_ (.A1(_15039_),
    .A2(_15042_),
    .ZN(_15043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24027_ (.A1(_15036_),
    .A2(_15043_),
    .B(_14516_),
    .ZN(_15044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24028_ (.A1(_14494_),
    .A2(_15861_),
    .ZN(_15045_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24029_ (.A1(_14738_),
    .A2(_14466_),
    .A3(_15045_),
    .Z(_15046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24030_ (.A1(_14388_),
    .A2(_14474_),
    .ZN(_15047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24031_ (.A1(_15046_),
    .A2(_15047_),
    .B(_14584_),
    .ZN(_15048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _24032_ (.A1(net509),
    .A2(_14549_),
    .B1(_14753_),
    .B2(_14707_),
    .ZN(_15049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24033_ (.A1(_15049_),
    .A2(_14497_),
    .ZN(_15050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24034_ (.A1(_15048_),
    .A2(_15050_),
    .ZN(_15051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24035_ (.A1(_15840_),
    .A2(_14572_),
    .B(_14634_),
    .ZN(_15052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24036_ (.A1(_14956_),
    .A2(_15052_),
    .B(_14484_),
    .ZN(_15053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24037_ (.A1(_14849_),
    .A2(_14504_),
    .ZN(_15054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24038_ (.A1(_14467_),
    .A2(_14613_),
    .A3(_15054_),
    .ZN(_15055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24039_ (.A1(_15053_),
    .A2(_15055_),
    .ZN(_15056_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24040_ (.A1(_15051_),
    .A2(_14540_),
    .A3(_15056_),
    .ZN(_15057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24041_ (.A1(_15044_),
    .A2(_15057_),
    .ZN(_15058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24042_ (.A1(_15031_),
    .A2(_15058_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _24043_ (.I(\sa20_sub[7] ),
    .ZN(_15059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24044_ (.A1(_12006_),
    .A2(_15059_),
    .ZN(_15060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24045_ (.A1(\sa20_sub[0] ),
    .A2(_12250_),
    .ZN(_15061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24046_ (.A1(_15060_),
    .A2(_15061_),
    .ZN(_15062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24047_ (.A1(_11964_),
    .A2(_15062_),
    .ZN(_15063_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24048_ (.A1(\sa20_sub[0] ),
    .A2(_12250_),
    .Z(_15064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24049_ (.A1(_15064_),
    .A2(net1175),
    .ZN(_15065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24050_ (.A1(_15065_),
    .A2(_15063_),
    .ZN(_15066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24051_ (.I(_15066_),
    .ZN(_15067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24052_ (.A1(_11977_),
    .A2(_12021_),
    .ZN(_15068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24053_ (.A1(_11984_),
    .A2(\sa02_sr[1] ),
    .ZN(_15069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24054_ (.A1(_15068_),
    .A2(_15069_),
    .ZN(_15070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24055_ (.I(_15070_),
    .ZN(_15071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24056_ (.A1(_15067_),
    .A2(_15071_),
    .ZN(_15072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24057_ (.A1(_15066_),
    .A2(_15070_),
    .ZN(_15073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24058_ (.A1(_15072_),
    .A2(_10402_),
    .A3(_15073_),
    .ZN(_15074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24059_ (.A1(_11203_),
    .A2(\text_in_r[49] ),
    .ZN(_15075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24060_ (.A1(_15074_),
    .A2(_15075_),
    .ZN(_15076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24061_ (.I(\u0.w[2][17] ),
    .ZN(_15077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24062_ (.A1(_15076_),
    .A2(_15077_),
    .ZN(_15078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24063_ (.A1(_15074_),
    .A2(\u0.w[2][17] ),
    .A3(_15075_),
    .ZN(_15079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24064_ (.A1(_15078_),
    .A2(_15079_),
    .ZN(_15871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24065_ (.A1(_11966_),
    .A2(_11980_),
    .ZN(_15080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24066_ (.A1(net1177),
    .A2(\sa12_sr[7] ),
    .ZN(_15081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24067_ (.A1(_15080_),
    .A2(_15081_),
    .ZN(_15082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24068_ (.A1(_15082_),
    .A2(net787),
    .ZN(_15083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24069_ (.A1(_15080_),
    .A2(_12002_),
    .A3(_15081_),
    .ZN(_15084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24070_ (.A1(_15083_),
    .A2(_15084_),
    .ZN(_15085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24071_ (.A1(_15085_),
    .A2(net633),
    .ZN(_15086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24072_ (.A1(_15083_),
    .A2(_15084_),
    .A3(_15062_),
    .ZN(_15087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24073_ (.A1(_15086_),
    .A2(_15087_),
    .B(_12193_),
    .ZN(_15088_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24074_ (.I(\text_in_r[48] ),
    .ZN(_15089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24075_ (.A1(_15089_),
    .A2(_10482_),
    .Z(_15090_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24076_ (.A1(_15088_),
    .A2(_15090_),
    .B(\u0.w[2][16] ),
    .ZN(_15091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24077_ (.A1(_15086_),
    .A2(_15087_),
    .ZN(_15092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24078_ (.A1(_15092_),
    .A2(_11279_),
    .ZN(_15093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24079_ (.I(\u0.w[2][16] ),
    .ZN(_15094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24080_ (.I(_15090_),
    .ZN(_15095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24081_ (.A1(_15093_),
    .A2(_15094_),
    .A3(_15095_),
    .ZN(_15096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24082_ (.A1(_15096_),
    .A2(_15091_),
    .ZN(_15874_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24083_ (.A1(_12027_),
    .A2(\sa31_sub[2] ),
    .Z(_15097_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24084_ (.A1(_12027_),
    .A2(\sa31_sub[2] ),
    .ZN(_15098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24085_ (.A1(_15097_),
    .A2(_15098_),
    .B(\sa02_sr[2] ),
    .ZN(_15099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24086_ (.A1(_12025_),
    .A2(_12030_),
    .ZN(_15100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24087_ (.A1(_12027_),
    .A2(\sa31_sub[2] ),
    .ZN(_15101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24088_ (.A1(_15100_),
    .A2(_12057_),
    .A3(_15101_),
    .ZN(_15102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24089_ (.A1(_15099_),
    .A2(_15102_),
    .ZN(_15103_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24090_ (.A1(\sa12_sr[1] ),
    .A2(\sa20_sub[1] ),
    .ZN(_15104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24091_ (.I(_15104_),
    .ZN(_15105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24092_ (.A1(_15103_),
    .A2(_15105_),
    .ZN(_15106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24093_ (.A1(_15099_),
    .A2(_15102_),
    .A3(_15104_),
    .ZN(_15107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24094_ (.A1(_15106_),
    .A2(_15107_),
    .B(_10381_),
    .ZN(_15108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24095_ (.I(\text_in_r[50] ),
    .ZN(_15109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24096_ (.A1(_15109_),
    .A2(net596),
    .Z(_15110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24097_ (.I(\u0.w[2][18] ),
    .ZN(_15111_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24098_ (.A1(_15108_),
    .A2(_15110_),
    .B(_15111_),
    .ZN(_15112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24099_ (.A1(_15106_),
    .A2(_15107_),
    .ZN(_15113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24100_ (.A1(_15113_),
    .A2(_10402_),
    .ZN(_15114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24101_ (.I(_15110_),
    .ZN(_15115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24102_ (.A1(_15114_),
    .A2(\u0.w[2][18] ),
    .A3(_15115_),
    .ZN(_15116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24103_ (.A1(_15112_),
    .A2(_15116_),
    .ZN(_15117_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24104_ (.I(_15117_),
    .Z(_15890_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24105_ (.A1(_15088_),
    .A2(_15090_),
    .B(_15094_),
    .ZN(_15118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24106_ (.A1(_15093_),
    .A2(\u0.w[2][16] ),
    .A3(_15095_),
    .ZN(_15119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24107_ (.A1(_15118_),
    .A2(_15119_),
    .ZN(_15865_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _24108_ (.A1(_15108_),
    .A2(_15110_),
    .B(\u0.w[2][18] ),
    .ZN(_15120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24109_ (.A1(_15114_),
    .A2(_15111_),
    .A3(_15115_),
    .ZN(_15121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24110_ (.A1(_15120_),
    .A2(_15121_),
    .ZN(_15122_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24111_ (.I(_15122_),
    .Z(_15883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24112_ (.A1(_15890_),
    .A2(_15872_),
    .ZN(_15123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24113_ (.A1(_15112_),
    .A2(_15116_),
    .A3(_15877_),
    .ZN(_15124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24114_ (.A1(_11980_),
    .A2(_12032_),
    .ZN(_15125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24115_ (.A1(net72),
    .A2(\sa12_sr[2] ),
    .ZN(_15126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24116_ (.A1(_15125_),
    .A2(_15126_),
    .ZN(_15127_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24117_ (.A1(\sa02_sr[3] ),
    .A2(_15127_),
    .Z(_15128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24118_ (.A1(_12025_),
    .A2(_15059_),
    .ZN(_15129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24119_ (.A1(_12027_),
    .A2(_12250_),
    .ZN(_15130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24120_ (.A1(_15129_),
    .A2(_15130_),
    .ZN(_15131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24121_ (.A1(_12056_),
    .A2(_15131_),
    .ZN(_15132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24122_ (.A1(_15059_),
    .A2(_12027_),
    .ZN(_15133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24123_ (.A1(_12025_),
    .A2(net49),
    .ZN(_15134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24124_ (.A1(_15133_),
    .A2(_15134_),
    .ZN(_15135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24125_ (.A1(_12069_),
    .A2(_15135_),
    .ZN(_15136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24126_ (.A1(_15132_),
    .A2(_15136_),
    .ZN(_15137_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24127_ (.I(_15137_),
    .ZN(_15138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24128_ (.A1(_15128_),
    .A2(_15138_),
    .ZN(_15139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24129_ (.A1(_15127_),
    .A2(\sa02_sr[3] ),
    .Z(_15140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24130_ (.A1(_15127_),
    .A2(\sa02_sr[3] ),
    .ZN(_15141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24131_ (.A1(_15140_),
    .A2(_15141_),
    .ZN(_15142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24132_ (.A1(_15142_),
    .A2(_15137_),
    .ZN(_15143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24133_ (.A1(_15139_),
    .A2(_10522_),
    .A3(_15143_),
    .ZN(_15144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24134_ (.A1(_10525_),
    .A2(\text_in_r[51] ),
    .ZN(_15145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24135_ (.A1(_15144_),
    .A2(_15145_),
    .ZN(_15146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24136_ (.I(\u0.w[2][19] ),
    .ZN(_15147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24137_ (.A1(_15146_),
    .A2(_15147_),
    .ZN(_15148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24138_ (.A1(_15144_),
    .A2(\u0.w[2][19] ),
    .A3(_15145_),
    .ZN(_15149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24139_ (.A1(_15148_),
    .A2(_15149_),
    .ZN(_15150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24140_ (.I(_15150_),
    .Z(_15151_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24141_ (.I(_15151_),
    .Z(_15152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24142_ (.A1(_15123_),
    .A2(_15124_),
    .B(_15152_),
    .ZN(_15153_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24143_ (.A1(\sa20_sub[4] ),
    .A2(\sa31_sub[4] ),
    .Z(_15154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24144_ (.I(_15154_),
    .ZN(_15155_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24145_ (.A1(\sa20_sub[3] ),
    .A2(_12250_),
    .Z(_15156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24146_ (.A1(_15155_),
    .A2(_15156_),
    .ZN(_15157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24147_ (.I(_15156_),
    .ZN(_15158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24148_ (.A1(_15158_),
    .A2(_15154_),
    .ZN(_15159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24149_ (.A1(_15157_),
    .A2(_15159_),
    .Z(_15160_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24150_ (.A1(\sa02_sr[4] ),
    .A2(_12080_),
    .Z(_15161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24151_ (.A1(_15160_),
    .A2(_15161_),
    .ZN(_15162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24152_ (.A1(_15157_),
    .A2(_15159_),
    .ZN(_15163_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24153_ (.A1(\sa02_sr[4] ),
    .A2(_12076_),
    .Z(_15164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24154_ (.A1(_15163_),
    .A2(_15164_),
    .ZN(_15165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24155_ (.A1(_15162_),
    .A2(_15165_),
    .A3(_13010_),
    .ZN(_15166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24156_ (.A1(_11385_),
    .A2(\text_in_r[52] ),
    .ZN(_15167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24157_ (.A1(_15166_),
    .A2(_15167_),
    .ZN(_15168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24158_ (.A1(_15168_),
    .A2(\u0.w[2][20] ),
    .ZN(_15169_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24159_ (.I(\u0.w[2][20] ),
    .ZN(_15170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24160_ (.A1(_15166_),
    .A2(_15170_),
    .A3(_15167_),
    .ZN(_15171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24161_ (.A1(_15169_),
    .A2(_15171_),
    .ZN(_15172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24162_ (.I(_15172_),
    .Z(_15173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24163_ (.I(_15868_),
    .ZN(_15174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24164_ (.A1(_15122_),
    .A2(_15174_),
    .ZN(_15175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24165_ (.A1(_15150_),
    .A2(_15175_),
    .ZN(_15176_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24166_ (.I(_15176_),
    .ZN(_15177_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _24167_ (.A1(_15153_),
    .A2(_15173_),
    .A3(_15177_),
    .Z(_15178_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24168_ (.A1(\sa12_sr[4] ),
    .A2(\sa20_sub[4] ),
    .ZN(_15179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24169_ (.I(\sa02_sr[5] ),
    .ZN(_15180_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24170_ (.A1(_15180_),
    .A2(_12151_),
    .Z(_15181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24171_ (.A1(_15179_),
    .A2(_15181_),
    .Z(_15182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24172_ (.A1(_15182_),
    .A2(_10585_),
    .ZN(_15183_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24173_ (.A1(_11348_),
    .A2(\text_in_r[53] ),
    .Z(_15184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24174_ (.A1(_15183_),
    .A2(_15184_),
    .ZN(_15185_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24175_ (.I(\u0.w[2][21] ),
    .ZN(_15186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24176_ (.A1(_15185_),
    .A2(_15186_),
    .ZN(_15187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24177_ (.A1(_15183_),
    .A2(\u0.w[2][21] ),
    .A3(_15184_),
    .ZN(_15188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24178_ (.A1(_15187_),
    .A2(_15188_),
    .ZN(_15189_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24179_ (.I(_15189_),
    .Z(_15190_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24180_ (.I(_15190_),
    .Z(_15191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24181_ (.I(_15872_),
    .ZN(_15192_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24182_ (.A1(_15883_),
    .A2(_15192_),
    .ZN(_15193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24183_ (.A1(_15146_),
    .A2(\u0.w[2][19] ),
    .ZN(_15194_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24184_ (.A1(_15144_),
    .A2(_15147_),
    .A3(_15145_),
    .ZN(_15195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24185_ (.A1(_15194_),
    .A2(_15195_),
    .ZN(_15196_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24186_ (.I(_15196_),
    .Z(_15197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24187_ (.A1(_15193_),
    .A2(_15197_),
    .ZN(_15198_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24188_ (.I(_15172_),
    .Z(_15199_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24189_ (.A1(_15198_),
    .A2(_15199_),
    .Z(_15200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24190_ (.A1(net1258),
    .A2(_15117_),
    .ZN(_15201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24191_ (.A1(_15201_),
    .A2(_15151_),
    .Z(_15202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24192_ (.A1(_15883_),
    .A2(net1217),
    .A3(net834),
    .ZN(_15203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24193_ (.A1(_15202_),
    .A2(_15203_),
    .ZN(_15204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24194_ (.A1(_15200_),
    .A2(_15204_),
    .ZN(_15205_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24195_ (.A1(_15178_),
    .A2(_15191_),
    .A3(_15205_),
    .ZN(_15206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24196_ (.A1(_15122_),
    .A2(_15192_),
    .ZN(_15207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24197_ (.A1(_15207_),
    .A2(_15151_),
    .Z(_15208_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24198_ (.A1(_15208_),
    .A2(_15173_),
    .ZN(_15209_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24199_ (.I(_15867_),
    .ZN(_15210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24200_ (.A1(_15890_),
    .A2(_15210_),
    .Z(_15211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _24201_ (.I(_15122_),
    .Z(_15212_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24202_ (.A1(_15212_),
    .A2(_15869_),
    .Z(_15213_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24203_ (.I(_15196_),
    .Z(_15214_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24204_ (.I(_15214_),
    .Z(_15215_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24205_ (.A1(_15211_),
    .A2(_15213_),
    .B(_15215_),
    .ZN(_15216_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24206_ (.I(_15190_),
    .Z(_15217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24207_ (.A1(_15209_),
    .A2(_15216_),
    .B(_15217_),
    .ZN(_15218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24208_ (.A1(net1217),
    .A2(_15212_),
    .ZN(_15219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24209_ (.I(_15219_),
    .ZN(_15220_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _24210_ (.A1(_15212_),
    .A2(_15875_),
    .ZN(_15221_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24211_ (.I(_15150_),
    .Z(_15222_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24212_ (.I(_15222_),
    .Z(_15223_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24213_ (.A1(_15220_),
    .A2(_15221_),
    .B(_15223_),
    .ZN(_15224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24214_ (.A1(_15212_),
    .A2(net835),
    .ZN(_15225_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24215_ (.I(_15196_),
    .Z(_15226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24216_ (.A1(_15120_),
    .A2(_15868_),
    .A3(_15121_),
    .ZN(_15227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24217_ (.A1(_15225_),
    .A2(_15226_),
    .A3(_15227_),
    .ZN(_15228_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24218_ (.I(_15199_),
    .Z(_15229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24219_ (.A1(_15224_),
    .A2(_15228_),
    .A3(_15229_),
    .ZN(_15230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24220_ (.A1(_15218_),
    .A2(_15230_),
    .ZN(_15231_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24221_ (.A1(\sa12_sr[5] ),
    .A2(\sa20_sub[5] ),
    .ZN(_15232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24222_ (.I(\sa02_sr[6] ),
    .ZN(_15233_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24223_ (.A1(_15233_),
    .A2(_12190_),
    .Z(_15234_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24224_ (.A1(_15232_),
    .A2(_15234_),
    .ZN(_15235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24225_ (.A1(_11385_),
    .A2(\text_in_r[54] ),
    .Z(_15236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24226_ (.A1(_15235_),
    .A2(_10585_),
    .B(_15236_),
    .ZN(_15237_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24227_ (.A1(\u0.w[2][22] ),
    .A2(_15237_),
    .Z(_15238_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24228_ (.I(_15238_),
    .ZN(_15239_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24229_ (.I(_15239_),
    .Z(_15240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24230_ (.A1(_15206_),
    .A2(_15231_),
    .A3(_15240_),
    .ZN(_15241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24231_ (.A1(net8),
    .A2(_15883_),
    .A3(net1048),
    .ZN(_15242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24232_ (.A1(_15120_),
    .A2(_15192_),
    .A3(_15121_),
    .ZN(_15243_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24233_ (.A1(_15242_),
    .A2(_15226_),
    .A3(_15243_),
    .ZN(_15244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24234_ (.A1(net1217),
    .A2(_15117_),
    .ZN(_15245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24235_ (.A1(_15212_),
    .A2(_15210_),
    .ZN(_15246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24236_ (.A1(_15245_),
    .A2(_15246_),
    .ZN(_15247_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24237_ (.I(_15151_),
    .Z(_15248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24238_ (.A1(_15168_),
    .A2(_15170_),
    .ZN(_15249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24239_ (.A1(_15166_),
    .A2(\u0.w[2][20] ),
    .A3(_15167_),
    .ZN(_15250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24240_ (.A1(_15249_),
    .A2(_15250_),
    .ZN(_15251_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24241_ (.I(_15251_),
    .Z(_15252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24242_ (.A1(_15247_),
    .A2(_15248_),
    .B(_15252_),
    .ZN(_15253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24243_ (.A1(_15890_),
    .A2(_15869_),
    .Z(_15254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24244_ (.A1(_15254_),
    .A2(_15197_),
    .ZN(_15255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24245_ (.A1(_15244_),
    .A2(_15253_),
    .A3(_15255_),
    .ZN(_15256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24246_ (.I(_15227_),
    .ZN(_15257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24247_ (.A1(_15226_),
    .A2(_15257_),
    .B(_15172_),
    .ZN(_15258_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24248_ (.I(_15222_),
    .Z(_15259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24249_ (.A1(_15259_),
    .A2(_15888_),
    .ZN(_15260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24250_ (.I(_15189_),
    .ZN(_15261_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24251_ (.I(_15261_),
    .Z(_15262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24252_ (.A1(_15258_),
    .A2(_15260_),
    .B(_15262_),
    .ZN(_15263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24253_ (.A1(_15256_),
    .A2(_15263_),
    .ZN(_15264_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24254_ (.I(_15877_),
    .ZN(_15265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24255_ (.A1(_15120_),
    .A2(_15265_),
    .A3(_15121_),
    .ZN(_15266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24256_ (.A1(_15150_),
    .A2(_15266_),
    .ZN(_15267_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24257_ (.I(_15267_),
    .ZN(_15268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24258_ (.A1(_15242_),
    .A2(_15268_),
    .ZN(_15269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24259_ (.A1(_15213_),
    .A2(_15214_),
    .ZN(_15270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24260_ (.A1(_15269_),
    .A2(_15229_),
    .A3(_15270_),
    .ZN(_15271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24261_ (.A1(_15213_),
    .A2(_15222_),
    .ZN(_15272_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24262_ (.A1(_15272_),
    .A2(_15252_),
    .Z(_15273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24263_ (.A1(_15117_),
    .A2(_15875_),
    .ZN(_15274_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24264_ (.A1(_15274_),
    .A2(_15196_),
    .Z(_15275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24265_ (.A1(_15242_),
    .A2(_15275_),
    .ZN(_15276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24266_ (.A1(_15273_),
    .A2(_15276_),
    .ZN(_15277_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24267_ (.I(_15261_),
    .Z(_15278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24268_ (.A1(_15271_),
    .A2(_15277_),
    .A3(_15278_),
    .ZN(_15279_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24269_ (.I(_15238_),
    .Z(_15280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24270_ (.A1(_15264_),
    .A2(_15279_),
    .A3(_15280_),
    .ZN(_15281_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24271_ (.A1(net1173),
    .A2(\sa12_sr[6] ),
    .Z(_15282_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24272_ (.A1(\sa20_sub[6] ),
    .A2(_15282_),
    .Z(_15283_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _24273_ (.A1(net49),
    .A2(net642),
    .A3(_15283_),
    .Z(_15284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _24274_ (.I0(_15284_),
    .I1(\text_in_r[55] ),
    .S(_10587_),
    .Z(_15285_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24275_ (.A1(\u0.w[2][23] ),
    .A2(_15285_),
    .ZN(_15286_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24276_ (.I(_15286_),
    .Z(_15287_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24277_ (.I(_15287_),
    .ZN(_15288_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24278_ (.A1(_15241_),
    .A2(_15281_),
    .A3(_15288_),
    .ZN(_15289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24279_ (.A1(_15117_),
    .A2(_15174_),
    .ZN(_15290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24280_ (.A1(_15290_),
    .A2(_15151_),
    .Z(_15291_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24281_ (.A1(_15291_),
    .A2(_15199_),
    .ZN(_15292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24282_ (.A1(\u0.w[2][17] ),
    .A2(_15076_),
    .ZN(_15293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24283_ (.A1(_15074_),
    .A2(_15077_),
    .A3(_15075_),
    .ZN(_15294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24284_ (.A1(_15294_),
    .A2(_15293_),
    .ZN(_15866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24285_ (.A1(net546),
    .A2(_15117_),
    .ZN(_15295_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24286_ (.I(_15295_),
    .Z(_15296_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24287_ (.A1(_15296_),
    .A2(_15222_),
    .ZN(_15297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24288_ (.I(_15297_),
    .ZN(_15298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24289_ (.I(_15175_),
    .ZN(_15299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24290_ (.A1(_15299_),
    .A2(_15197_),
    .ZN(_15300_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24291_ (.A1(_15292_),
    .A2(_15298_),
    .A3(_15300_),
    .Z(_15301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24292_ (.A1(_15246_),
    .A2(_15151_),
    .Z(_15302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24293_ (.A1(_15221_),
    .A2(_15197_),
    .ZN(_15303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24294_ (.A1(_15302_),
    .A2(_15303_),
    .Z(_15304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24295_ (.A1(_15890_),
    .A2(_15867_),
    .ZN(_15305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24296_ (.A1(_15177_),
    .A2(_15305_),
    .ZN(_15306_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24297_ (.I(_15251_),
    .Z(_15307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24298_ (.A1(_15304_),
    .A2(_15306_),
    .B(_15307_),
    .ZN(_15308_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24299_ (.A1(_15301_),
    .A2(_15308_),
    .B(_15191_),
    .ZN(_15309_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24300_ (.I(_15875_),
    .ZN(_15310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24301_ (.A1(_15212_),
    .A2(_15310_),
    .ZN(_15311_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24302_ (.A1(_15867_),
    .A2(_15883_),
    .B(_15311_),
    .ZN(_15312_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24303_ (.I(_15251_),
    .Z(_15313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24304_ (.A1(_15312_),
    .A2(_15259_),
    .B(_15313_),
    .ZN(_15314_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24305_ (.A1(net8),
    .A2(net1220),
    .A3(_15890_),
    .ZN(_15315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24306_ (.A1(_15175_),
    .A2(_15197_),
    .Z(_15316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24307_ (.A1(_15315_),
    .A2(_15316_),
    .ZN(_15317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24308_ (.A1(_15314_),
    .A2(_15317_),
    .ZN(_15318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24309_ (.A1(_15219_),
    .A2(_15214_),
    .Z(_15319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24310_ (.A1(net10),
    .A2(net1048),
    .ZN(_15320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24311_ (.A1(_15319_),
    .A2(_15320_),
    .ZN(_15321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24312_ (.A1(net835),
    .A2(net1050),
    .ZN(_15322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24313_ (.A1(_15322_),
    .A2(_15152_),
    .A3(_15245_),
    .ZN(_15323_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24314_ (.I(_15251_),
    .Z(_15324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24315_ (.A1(_15321_),
    .A2(_15323_),
    .A3(_15324_),
    .ZN(_15325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24316_ (.A1(_15318_),
    .A2(_15278_),
    .A3(_15325_),
    .ZN(_15326_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24317_ (.A1(_15309_),
    .A2(_15326_),
    .A3(_15280_),
    .ZN(_15327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24318_ (.A1(_15201_),
    .A2(_15196_),
    .ZN(_15328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24319_ (.A1(_15328_),
    .A2(_15199_),
    .Z(_15329_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24320_ (.A1(net8),
    .A2(net1050),
    .A3(_15890_),
    .ZN(_15330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24321_ (.A1(_15330_),
    .A2(_15208_),
    .ZN(_15331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24322_ (.A1(_15329_),
    .A2(_15331_),
    .B(_15190_),
    .ZN(_15332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24323_ (.A1(_15122_),
    .A2(net1049),
    .ZN(_15333_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24324_ (.A1(_15333_),
    .A2(_15214_),
    .Z(_15334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24325_ (.A1(_15334_),
    .A2(_15330_),
    .ZN(_15335_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24326_ (.I(_15881_),
    .ZN(_15336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24327_ (.A1(_15117_),
    .A2(_15336_),
    .ZN(_15337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24328_ (.A1(_15177_),
    .A2(_15337_),
    .ZN(_15338_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24329_ (.A1(_15335_),
    .A2(_15338_),
    .A3(_15307_),
    .ZN(_15339_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24330_ (.I(_15238_),
    .Z(_15340_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24331_ (.A1(_15332_),
    .A2(_15339_),
    .B(_15340_),
    .ZN(_15341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24332_ (.A1(_15270_),
    .A2(_15172_),
    .ZN(_15342_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24333_ (.A1(_15342_),
    .A2(_15297_),
    .ZN(_15343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24334_ (.A1(_15343_),
    .A2(_15204_),
    .ZN(_15344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24335_ (.A1(_15212_),
    .A2(_15336_),
    .ZN(_15345_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24336_ (.A1(_15345_),
    .A2(_15222_),
    .Z(_15346_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24337_ (.I(_15172_),
    .Z(_15347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24338_ (.A1(_15346_),
    .A2(_15201_),
    .B(_15347_),
    .ZN(_15348_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24339_ (.I(_15214_),
    .Z(_15349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24340_ (.A1(net10),
    .A2(_15212_),
    .ZN(_15350_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24341_ (.A1(_15330_),
    .A2(_15349_),
    .A3(_15350_),
    .ZN(_15351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24342_ (.A1(_15348_),
    .A2(_15351_),
    .ZN(_15352_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24343_ (.I(_15190_),
    .Z(_15353_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24344_ (.A1(_15344_),
    .A2(_15352_),
    .A3(_15353_),
    .ZN(_15354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24345_ (.A1(_15341_),
    .A2(_15354_),
    .B(_15288_),
    .ZN(_15355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24346_ (.A1(_15327_),
    .A2(_15355_),
    .ZN(_15356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24347_ (.A1(_15289_),
    .A2(_15356_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24348_ (.A1(_15208_),
    .A2(_15296_),
    .ZN(_15357_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24349_ (.I(_15172_),
    .Z(_15358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24350_ (.A1(_15219_),
    .A2(_15305_),
    .A3(_15215_),
    .ZN(_15359_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24351_ (.A1(_15357_),
    .A2(_15358_),
    .A3(_15359_),
    .ZN(_15360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24352_ (.A1(_15213_),
    .A2(_15349_),
    .B(_15347_),
    .ZN(_15361_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24353_ (.A1(_15245_),
    .A2(_15152_),
    .Z(_15362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24354_ (.A1(_15246_),
    .A2(_15227_),
    .ZN(_15363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24355_ (.A1(_15363_),
    .A2(_15223_),
    .ZN(_15364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24356_ (.A1(_15361_),
    .A2(_15362_),
    .A3(_15364_),
    .ZN(_15365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24357_ (.A1(_15360_),
    .A2(_15365_),
    .A3(_15262_),
    .ZN(_15366_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _24358_ (.I(_15328_),
    .ZN(_15367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24359_ (.A1(_15367_),
    .A2(net548),
    .ZN(_15368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24360_ (.A1(_15199_),
    .A2(net1047),
    .Z(_15369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24361_ (.A1(_15369_),
    .A2(_15368_),
    .B(_15261_),
    .ZN(_15370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24362_ (.A1(_15345_),
    .A2(_15214_),
    .Z(_15371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24363_ (.I(_15869_),
    .ZN(_15372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24364_ (.A1(_15117_),
    .A2(_15372_),
    .ZN(_15373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24365_ (.A1(_15371_),
    .A2(_15373_),
    .B(_15347_),
    .ZN(_15374_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24366_ (.A1(_15212_),
    .A2(_15868_),
    .Z(_15375_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _24367_ (.I(_15375_),
    .ZN(_15376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24368_ (.A1(_15315_),
    .A2(_15248_),
    .A3(_15376_),
    .ZN(_15377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24369_ (.A1(_15374_),
    .A2(_15377_),
    .ZN(_15378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24370_ (.A1(_15370_),
    .A2(_15378_),
    .ZN(_15379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24371_ (.A1(_15379_),
    .A2(_15366_),
    .B(_15280_),
    .ZN(_15380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24372_ (.A1(_15334_),
    .A2(_15305_),
    .ZN(_15381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24373_ (.A1(_15151_),
    .A2(_15883_),
    .Z(_15382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24374_ (.A1(net8),
    .A2(net1217),
    .ZN(_15383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24375_ (.A1(_15382_),
    .A2(_15383_),
    .ZN(_15384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24376_ (.A1(_15381_),
    .A2(_15384_),
    .ZN(_15385_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _24377_ (.A1(_15196_),
    .A2(_15212_),
    .ZN(_15386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24378_ (.A1(_15386_),
    .A2(_15322_),
    .ZN(_15387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24379_ (.A1(_15387_),
    .A2(_15252_),
    .ZN(_15388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24380_ (.A1(net548),
    .A2(_15275_),
    .ZN(_15389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24381_ (.A1(_15389_),
    .A2(_15358_),
    .ZN(_15390_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24382_ (.A1(_15385_),
    .A2(_15388_),
    .B(_15390_),
    .ZN(_15391_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24383_ (.I(_15891_),
    .ZN(_15392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24384_ (.A1(_15259_),
    .A2(_15392_),
    .Z(_15393_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24385_ (.I(_15252_),
    .Z(_15394_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24386_ (.A1(_15393_),
    .A2(_15394_),
    .B(_15353_),
    .ZN(_15395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24387_ (.A1(_15190_),
    .A2(_15252_),
    .Z(_15396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24388_ (.A1(_15357_),
    .A2(_15396_),
    .ZN(_15397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24389_ (.A1(net836),
    .A2(_15890_),
    .ZN(_15398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24390_ (.A1(_15319_),
    .A2(_15398_),
    .ZN(_15399_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24391_ (.I(_15399_),
    .ZN(_15400_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24392_ (.A1(_15397_),
    .A2(_15400_),
    .B(_15340_),
    .ZN(_15401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24393_ (.A1(_15391_),
    .A2(_15395_),
    .B(_15401_),
    .ZN(_15402_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24394_ (.A1(_15380_),
    .A2(_15402_),
    .B(_15287_),
    .ZN(_15403_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24395_ (.I(_15197_),
    .Z(_15404_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24396_ (.A1(_15383_),
    .A2(_15883_),
    .A3(_15404_),
    .ZN(_15405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24397_ (.A1(_15337_),
    .A2(_15151_),
    .Z(_15406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24398_ (.A1(_15406_),
    .A2(_15350_),
    .ZN(_15407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24399_ (.A1(_15405_),
    .A2(_15407_),
    .A3(_15324_),
    .ZN(_15408_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24400_ (.A1(_15883_),
    .A2(_15872_),
    .Z(_15409_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24401_ (.I(_15251_),
    .Z(_15410_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24402_ (.A1(_15409_),
    .A2(_15349_),
    .B(_15410_),
    .ZN(_15411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24403_ (.A1(_15377_),
    .A2(_15411_),
    .ZN(_15412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24404_ (.A1(_15408_),
    .A2(_15412_),
    .A3(_15278_),
    .ZN(_15413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24405_ (.A1(net10),
    .A2(net1219),
    .ZN(_15414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24406_ (.A1(_15202_),
    .A2(_15414_),
    .ZN(_15415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24407_ (.A1(_15214_),
    .A2(_15227_),
    .Z(_15416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24408_ (.A1(_15416_),
    .A2(_15333_),
    .ZN(_15417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24409_ (.A1(_15415_),
    .A2(_15358_),
    .A3(_15417_),
    .ZN(_15418_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24410_ (.A1(_15299_),
    .A2(_15193_),
    .B(_15248_),
    .ZN(_15419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24411_ (.A1(_15247_),
    .A2(_15349_),
    .ZN(_15420_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24412_ (.A1(_15419_),
    .A2(_15420_),
    .A3(_15307_),
    .ZN(_15421_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24413_ (.A1(_15418_),
    .A2(_15421_),
    .A3(_15353_),
    .ZN(_15422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24414_ (.A1(_15413_),
    .A2(_15422_),
    .A3(_15240_),
    .ZN(_15423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24415_ (.A1(_15346_),
    .A2(_15290_),
    .B(_15410_),
    .ZN(_15424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24416_ (.A1(_15424_),
    .A2(_15244_),
    .ZN(_15425_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24417_ (.A1(_15198_),
    .A2(_15251_),
    .Z(_15426_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24418_ (.I(_15151_),
    .Z(_15427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24419_ (.A1(_15398_),
    .A2(_15427_),
    .ZN(_15428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24420_ (.A1(_15426_),
    .A2(_15350_),
    .A3(_15428_),
    .ZN(_15429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24421_ (.A1(_15425_),
    .A2(_15429_),
    .A3(_15353_),
    .ZN(_15430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24422_ (.A1(_15207_),
    .A2(_15196_),
    .Z(_15431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24423_ (.A1(_15431_),
    .A2(_15245_),
    .ZN(_15432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24424_ (.A1(_15201_),
    .A2(_15175_),
    .A3(_15248_),
    .ZN(_15433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24425_ (.A1(_15432_),
    .A2(_15433_),
    .A3(_15307_),
    .ZN(_15434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24426_ (.A1(_15386_),
    .A2(_15322_),
    .B(_15410_),
    .ZN(_15435_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24427_ (.A1(_15320_),
    .A2(_15225_),
    .A3(_15226_),
    .ZN(_15436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24428_ (.A1(_15435_),
    .A2(_15436_),
    .ZN(_15437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24429_ (.A1(_15434_),
    .A2(_15437_),
    .A3(_15262_),
    .ZN(_15438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24430_ (.A1(_15430_),
    .A2(_15280_),
    .A3(_15438_),
    .ZN(_15439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24431_ (.A1(_15423_),
    .A2(_15439_),
    .A3(_15288_),
    .ZN(_15440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24432_ (.A1(_15403_),
    .A2(_15440_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24433_ (.A1(_15296_),
    .A2(_15248_),
    .A3(_15124_),
    .ZN(_15441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24434_ (.A1(_15120_),
    .A2(_15121_),
    .A3(_15881_),
    .ZN(_15442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24435_ (.A1(_15219_),
    .A2(_15226_),
    .A3(_15442_),
    .ZN(_15443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24436_ (.A1(_15441_),
    .A2(_15313_),
    .A3(_15443_),
    .ZN(_15444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24437_ (.A1(_15333_),
    .A2(_15197_),
    .A3(_15266_),
    .ZN(_15445_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24438_ (.A1(net837),
    .A2(_15222_),
    .A3(_15227_),
    .ZN(_15446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24439_ (.A1(_15446_),
    .A2(_15445_),
    .ZN(_15447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24440_ (.A1(_15447_),
    .A2(_15173_),
    .ZN(_15448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24441_ (.A1(_15444_),
    .A2(_15448_),
    .A3(_15262_),
    .ZN(_15449_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24442_ (.A1(net8),
    .A2(_15890_),
    .ZN(_15450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24443_ (.A1(_15222_),
    .A2(_15243_),
    .ZN(_15451_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24444_ (.A1(_15450_),
    .A2(_15451_),
    .ZN(_15452_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24445_ (.A1(_15452_),
    .A2(_15153_),
    .B(_15173_),
    .ZN(_15453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24446_ (.A1(_15333_),
    .A2(_15152_),
    .A3(_15243_),
    .ZN(_15454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24447_ (.A1(_15442_),
    .A2(_15124_),
    .ZN(_15455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24448_ (.A1(_15455_),
    .A2(_15226_),
    .ZN(_15456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24449_ (.A1(_15454_),
    .A2(_15456_),
    .ZN(_15457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24450_ (.A1(_15457_),
    .A2(_15313_),
    .ZN(_15458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24451_ (.A1(_15453_),
    .A2(_15458_),
    .A3(_15353_),
    .ZN(_15459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24452_ (.A1(_15459_),
    .A2(_15449_),
    .ZN(_15460_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24453_ (.A1(_15240_),
    .A2(_15460_),
    .B(_15288_),
    .ZN(_15461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24454_ (.A1(_15322_),
    .A2(_15225_),
    .A3(_15152_),
    .ZN(_15462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24455_ (.A1(_15431_),
    .A2(_15337_),
    .ZN(_15463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24456_ (.A1(_15462_),
    .A2(_15463_),
    .ZN(_15464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24457_ (.A1(_15464_),
    .A2(_15307_),
    .ZN(_15465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24458_ (.A1(_15333_),
    .A2(_15243_),
    .ZN(_15466_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24459_ (.A1(_15466_),
    .A2(_15152_),
    .A3(_15350_),
    .ZN(_15467_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24460_ (.A1(_15467_),
    .A2(_15173_),
    .A3(_15228_),
    .ZN(_15468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24461_ (.A1(_15465_),
    .A2(_15468_),
    .ZN(_15469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24462_ (.A1(_15469_),
    .A2(_15191_),
    .ZN(_15470_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24463_ (.A1(_15315_),
    .A2(_15259_),
    .A3(_15345_),
    .ZN(_15471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24464_ (.A1(_15330_),
    .A2(_15215_),
    .ZN(_15472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24465_ (.A1(_15471_),
    .A2(_15229_),
    .A3(_15472_),
    .ZN(_15473_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24466_ (.A1(_15220_),
    .A2(_15254_),
    .B(_15427_),
    .ZN(_15474_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24467_ (.A1(_15398_),
    .A2(_15349_),
    .A3(net837),
    .ZN(_15475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24468_ (.A1(_15474_),
    .A2(_15475_),
    .A3(_15324_),
    .ZN(_15476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24469_ (.A1(_15473_),
    .A2(_15278_),
    .A3(_15476_),
    .ZN(_15477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24470_ (.A1(_15470_),
    .A2(_15477_),
    .A3(_15280_),
    .ZN(_15478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24471_ (.A1(_15461_),
    .A2(_15478_),
    .ZN(_15479_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24472_ (.A1(_15296_),
    .A2(_15201_),
    .ZN(_15480_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24473_ (.A1(_15372_),
    .A2(_15192_),
    .Z(_15481_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24474_ (.A1(_15890_),
    .A2(_15481_),
    .Z(_15482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24475_ (.I(_15482_),
    .ZN(_15483_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24476_ (.A1(_15480_),
    .A2(_15483_),
    .B(_15259_),
    .ZN(_15484_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24477_ (.A1(_15484_),
    .A2(_15394_),
    .A3(_15389_),
    .ZN(_15485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24478_ (.A1(_15302_),
    .A2(_15199_),
    .Z(_15486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24479_ (.A1(_15177_),
    .A2(_15243_),
    .ZN(_15487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24480_ (.A1(_15487_),
    .A2(_15486_),
    .B(_15217_),
    .ZN(_15488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24481_ (.A1(_15485_),
    .A2(_15488_),
    .ZN(_15489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24482_ (.A1(_15895_),
    .A2(_15349_),
    .B(_15347_),
    .ZN(_15490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24483_ (.A1(_15462_),
    .A2(_15490_),
    .B(_15262_),
    .ZN(_15491_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24484_ (.A1(_15226_),
    .A2(_15886_),
    .Z(_15492_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24485_ (.A1(_15472_),
    .A2(_15229_),
    .A3(_15492_),
    .ZN(_15493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24486_ (.A1(_15491_),
    .A2(_15493_),
    .ZN(_15494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24487_ (.A1(_15489_),
    .A2(_15494_),
    .A3(_15280_),
    .ZN(_15495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24488_ (.A1(_15225_),
    .A2(_15226_),
    .ZN(_15496_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24489_ (.A1(_15496_),
    .A2(_15211_),
    .ZN(_15497_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24490_ (.A1(_15311_),
    .A2(_15152_),
    .A3(_15227_),
    .Z(_15498_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24491_ (.A1(_15497_),
    .A2(_15498_),
    .B(_15324_),
    .ZN(_15499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24492_ (.A1(_15320_),
    .A2(_15225_),
    .A3(_15248_),
    .ZN(_15500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24493_ (.A1(_15404_),
    .A2(_15392_),
    .ZN(_15501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24494_ (.A1(_15500_),
    .A2(_15358_),
    .A3(_15501_),
    .ZN(_15502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24495_ (.A1(_15499_),
    .A2(_15191_),
    .A3(_15502_),
    .ZN(_15503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24496_ (.A1(net1051),
    .A2(_15291_),
    .ZN(_15504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24497_ (.A1(_15888_),
    .A2(_15215_),
    .B(_15252_),
    .ZN(_15505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24498_ (.A1(_15504_),
    .A2(_15505_),
    .B(_15190_),
    .ZN(_15506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24499_ (.A1(_15296_),
    .A2(_15248_),
    .A3(_15333_),
    .ZN(_15507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24500_ (.A1(_15228_),
    .A2(_15507_),
    .A3(_15307_),
    .ZN(_15508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24501_ (.A1(_15506_),
    .A2(_15508_),
    .B(_15340_),
    .ZN(_15509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24502_ (.A1(_15503_),
    .A2(_15509_),
    .ZN(_15510_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24503_ (.A1(_15495_),
    .A2(_15510_),
    .A3(_15288_),
    .ZN(_15511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24504_ (.A1(_15479_),
    .A2(_15511_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24505_ (.A1(_15382_),
    .A2(_15210_),
    .B(_15199_),
    .ZN(_15512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24506_ (.A1(_15245_),
    .A2(_15311_),
    .Z(_15513_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24507_ (.A1(_15513_),
    .A2(_15248_),
    .Z(_15514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24508_ (.I(_15290_),
    .ZN(_15515_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24509_ (.A1(_15515_),
    .A2(_15152_),
    .Z(_15516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24510_ (.I(_15516_),
    .ZN(_15517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24511_ (.A1(_15512_),
    .A2(_15514_),
    .A3(_15517_),
    .ZN(_15518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24512_ (.A1(_15296_),
    .A2(_15197_),
    .ZN(_15519_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24513_ (.A1(_15519_),
    .A2(_15375_),
    .Z(_15520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24514_ (.A1(_15346_),
    .A2(_15243_),
    .ZN(_15521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24515_ (.A1(_15520_),
    .A2(_15229_),
    .A3(_15521_),
    .ZN(_15522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24516_ (.A1(_15518_),
    .A2(_15522_),
    .A3(_15278_),
    .ZN(_15523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24517_ (.A1(_15296_),
    .A2(_15349_),
    .A3(_15333_),
    .ZN(_15524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24518_ (.A1(_15292_),
    .A2(_15524_),
    .B(_15261_),
    .ZN(_15525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24519_ (.A1(_15319_),
    .A2(_15322_),
    .ZN(_15526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24520_ (.A1(_15177_),
    .A2(_15296_),
    .ZN(_15527_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24521_ (.A1(_15526_),
    .A2(_15527_),
    .A3(_15358_),
    .ZN(_15528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24522_ (.A1(_15525_),
    .A2(_15528_),
    .B(_15240_),
    .ZN(_15529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24523_ (.A1(_15523_),
    .A2(_15529_),
    .B(_15287_),
    .ZN(_15530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24524_ (.A1(_15296_),
    .A2(_15151_),
    .Z(_15531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24525_ (.A1(_15531_),
    .A2(_15513_),
    .ZN(_15532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24526_ (.A1(_15416_),
    .A2(_15350_),
    .A3(_15333_),
    .ZN(_15533_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24527_ (.A1(_15532_),
    .A2(_15173_),
    .A3(_15533_),
    .Z(_15534_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _24528_ (.A1(_15299_),
    .A2(_15222_),
    .A3(_15221_),
    .Z(_15535_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24529_ (.A1(_15535_),
    .A2(_15313_),
    .A3(_15323_),
    .Z(_15536_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24530_ (.A1(_15534_),
    .A2(_15536_),
    .B(_15278_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24531_ (.A1(_15320_),
    .A2(_15245_),
    .A3(_15172_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24532_ (.I(_15382_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24533_ (.A1(_00550_),
    .A2(_00551_),
    .B(_15262_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24534_ (.A1(_15214_),
    .A2(_15266_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24535_ (.A1(_00553_),
    .A2(_15376_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24536_ (.A1(_15407_),
    .A2(_00554_),
    .A3(_15394_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24537_ (.A1(_00552_),
    .A2(_00555_),
    .B(_15340_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24538_ (.A1(_00549_),
    .A2(_00556_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24539_ (.A1(_15530_),
    .A2(_00557_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24540_ (.I(_15124_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24541_ (.A1(_15223_),
    .A2(_00559_),
    .B(_15190_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24542_ (.A1(_00560_),
    .A2(_15445_),
    .B(_15307_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24543_ (.A1(_15367_),
    .A2(_15175_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24544_ (.A1(_15883_),
    .A2(_15481_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24545_ (.A1(_00563_),
    .A2(_15222_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24546_ (.I(_15337_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24547_ (.A1(_00564_),
    .A2(_00565_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24548_ (.A1(_00562_),
    .A2(_00566_),
    .A3(_15217_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24549_ (.A1(_00561_),
    .A2(_00567_),
    .B(_15240_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24550_ (.A1(_15275_),
    .A2(_15225_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24551_ (.A1(_00569_),
    .A2(_15516_),
    .B(_15190_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24552_ (.I(_15300_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _24553_ (.A1(_00571_),
    .A2(_15261_),
    .B1(_15223_),
    .B2(_15213_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24554_ (.A1(_00570_),
    .A2(_00572_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24555_ (.A1(_00573_),
    .A2(_15394_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24556_ (.A1(_00568_),
    .A2(_00574_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24557_ (.A1(_15268_),
    .A2(_00563_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24558_ (.A1(_15389_),
    .A2(_00576_),
    .A3(_15358_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24559_ (.I(_15443_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24560_ (.A1(_00578_),
    .A2(_15307_),
    .B(_15261_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24561_ (.A1(_00577_),
    .A2(_00579_),
    .B(_15340_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24562_ (.I(_15201_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24563_ (.A1(_00581_),
    .A2(_00559_),
    .B(_15152_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24564_ (.A1(_15316_),
    .A2(_15337_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24565_ (.A1(_00582_),
    .A2(_00583_),
    .A3(_15324_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24566_ (.A1(_15253_),
    .A2(_15436_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24567_ (.A1(_00584_),
    .A2(_00585_),
    .A3(_15278_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24568_ (.A1(_00580_),
    .A2(_00586_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24569_ (.A1(_00575_),
    .A2(_00587_),
    .A3(_15287_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24570_ (.A1(_00558_),
    .A2(_00588_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24571_ (.A1(_15268_),
    .A2(_15350_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24572_ (.A1(_15450_),
    .A2(_15404_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24573_ (.A1(_15220_),
    .A2(_15226_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _24574_ (.A1(_15394_),
    .A2(_00589_),
    .A3(_00590_),
    .A4(_00591_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24575_ (.I(_15879_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24576_ (.A1(_00593_),
    .A2(_15404_),
    .B(_15410_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24577_ (.A1(_15259_),
    .A2(_15227_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24578_ (.A1(_00594_),
    .A2(_00595_),
    .B(_15217_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24579_ (.A1(_00592_),
    .A2(_00596_),
    .B(_15240_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24580_ (.A1(_15322_),
    .A2(_15295_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24581_ (.A1(_00598_),
    .A2(_15152_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24582_ (.A1(_15268_),
    .A2(_15219_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24583_ (.A1(_00599_),
    .A2(_00600_),
    .A3(_15394_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24584_ (.A1(_15216_),
    .A2(_15323_),
    .A3(_15229_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24585_ (.A1(_00601_),
    .A2(_00602_),
    .A3(_15191_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24586_ (.A1(_00597_),
    .A2(_00603_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24587_ (.A1(_15302_),
    .A2(_15252_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24588_ (.A1(_00605_),
    .A2(_15298_),
    .A3(_15357_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24589_ (.A1(_15319_),
    .A2(_15337_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24590_ (.A1(_15386_),
    .A2(_15313_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24591_ (.A1(_00607_),
    .A2(_00608_),
    .B(_15262_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24592_ (.A1(_00606_),
    .A2(_00609_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24593_ (.A1(_15373_),
    .A2(_15214_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24594_ (.A1(_00611_),
    .A2(_15347_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24595_ (.A1(_15315_),
    .A2(_15223_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24596_ (.A1(_00612_),
    .A2(_00613_),
    .B(_15217_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24597_ (.A1(_15431_),
    .A2(_15227_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24598_ (.A1(_15204_),
    .A2(_00615_),
    .A3(_15358_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24599_ (.A1(_00614_),
    .A2(_00616_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24600_ (.A1(_00610_),
    .A2(_00617_),
    .A3(_15240_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24601_ (.A1(_00604_),
    .A2(_15287_),
    .A3(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24602_ (.A1(_15531_),
    .A2(net1051),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24603_ (.A1(_00620_),
    .A2(_15394_),
    .A3(_15463_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24604_ (.A1(_15398_),
    .A2(_15246_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24605_ (.A1(_00622_),
    .A2(_15259_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24606_ (.A1(_15244_),
    .A2(_15229_),
    .A3(_00623_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24607_ (.A1(_00621_),
    .A2(_00624_),
    .A3(_15191_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24608_ (.A1(_15257_),
    .A2(_15222_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24609_ (.A1(_00626_),
    .A2(_00559_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24610_ (.A1(_15426_),
    .A2(_00627_),
    .B(_15217_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24611_ (.A1(_15371_),
    .A2(_15290_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24612_ (.A1(_15269_),
    .A2(_00629_),
    .A3(_15358_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24613_ (.A1(_00628_),
    .A2(_00630_),
    .B(_15239_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24614_ (.A1(_00631_),
    .A2(_00625_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24615_ (.A1(_15296_),
    .A2(_15219_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24616_ (.A1(_00633_),
    .A2(_15259_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24617_ (.A1(_00634_),
    .A2(_15381_),
    .A3(_15358_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24618_ (.A1(_15213_),
    .A2(_15347_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24619_ (.A1(_00636_),
    .A2(_15267_),
    .B(_15190_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24620_ (.A1(_00635_),
    .A2(_00637_),
    .B(_15340_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24621_ (.A1(_00598_),
    .A2(_15404_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24622_ (.A1(_15350_),
    .A2(_15427_),
    .A3(_15305_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24623_ (.A1(_00639_),
    .A2(_15394_),
    .A3(_00640_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24624_ (.A1(_15500_),
    .A2(_15399_),
    .A3(_15173_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24625_ (.A1(_00641_),
    .A2(_00642_),
    .A3(_15353_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24626_ (.A1(_00638_),
    .A2(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24627_ (.A1(_00632_),
    .A2(_00644_),
    .A3(_15288_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24628_ (.A1(_00645_),
    .A2(_00619_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24629_ (.A1(net10),
    .A2(_15248_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24630_ (.A1(_00599_),
    .A2(_15173_),
    .A3(_00646_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24631_ (.A1(net548),
    .A2(_15274_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24632_ (.A1(_15367_),
    .A2(_15383_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24633_ (.A1(_00649_),
    .A2(_15313_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24634_ (.A1(_00648_),
    .A2(_15259_),
    .B(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24635_ (.A1(_00647_),
    .A2(_00651_),
    .B(_15278_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24636_ (.A1(_00611_),
    .A2(_15225_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24637_ (.A1(_00653_),
    .A2(_00626_),
    .B(_15313_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24638_ (.A1(_15226_),
    .A2(_15442_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _24639_ (.A1(_15176_),
    .A2(_15211_),
    .B(_00655_),
    .C(_15347_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24640_ (.A1(_00654_),
    .A2(_00656_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24641_ (.A1(_00657_),
    .A2(_15191_),
    .B(_15240_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24642_ (.A1(_00652_),
    .A2(_00658_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24643_ (.A1(_15316_),
    .A2(_15313_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24644_ (.A1(_00660_),
    .A2(_00582_),
    .B(_15261_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24645_ (.A1(_15388_),
    .A2(_15431_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24646_ (.A1(_00661_),
    .A2(_00662_),
    .B(_15340_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24647_ (.A1(_15406_),
    .A2(_15207_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24648_ (.A1(_15343_),
    .A2(_00664_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24649_ (.A1(net1051),
    .A2(_00553_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24650_ (.A1(_15223_),
    .A2(_15872_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24651_ (.A1(_15273_),
    .A2(_00666_),
    .A3(_00667_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24652_ (.A1(_00665_),
    .A2(_00668_),
    .A3(_15278_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24653_ (.A1(_00663_),
    .A2(_00669_),
    .B(_15287_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24654_ (.A1(_00659_),
    .A2(_00670_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24655_ (.A1(net1218),
    .A2(_15427_),
    .B(_15410_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24656_ (.A1(_15321_),
    .A2(_00672_),
    .B(_15217_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24657_ (.A1(_15330_),
    .A2(_15177_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24658_ (.A1(_00553_),
    .A2(_15350_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24659_ (.A1(_00674_),
    .A2(_00675_),
    .A3(_15324_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24660_ (.A1(_00673_),
    .A2(_00676_),
    .B(_15340_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24661_ (.A1(_15200_),
    .A2(_15204_),
    .A3(_00591_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24662_ (.A1(_15203_),
    .A2(_15215_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24663_ (.A1(_15221_),
    .A2(_15427_),
    .B(_15347_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24664_ (.A1(_00679_),
    .A2(_00565_),
    .B(_00680_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24665_ (.A1(_00678_),
    .A2(_00681_),
    .A3(_15353_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24666_ (.A1(_00677_),
    .A2(_00682_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24667_ (.I(_15406_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24668_ (.A1(_15426_),
    .A2(_00684_),
    .B(_15217_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24669_ (.I(net548),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24670_ (.A1(_00564_),
    .A2(_15199_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24671_ (.A1(_15472_),
    .A2(_00686_),
    .B(_00687_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24672_ (.A1(_00685_),
    .A2(_00688_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24673_ (.A1(_15310_),
    .A2(_15427_),
    .B(_15410_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24674_ (.A1(_00679_),
    .A2(_00690_),
    .B(_15261_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24675_ (.A1(_15376_),
    .A2(_15337_),
    .A3(_15349_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24676_ (.A1(_15177_),
    .A2(_15274_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24677_ (.A1(_00692_),
    .A2(_00693_),
    .A3(_15324_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24678_ (.A1(_00691_),
    .A2(_00694_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24679_ (.A1(_00689_),
    .A2(_00695_),
    .A3(_15280_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24680_ (.A1(_00683_),
    .A2(_00696_),
    .A3(_15287_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24681_ (.A1(_00671_),
    .A2(_00697_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24682_ (.A1(_15123_),
    .A2(_15124_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _24683_ (.A1(_00698_),
    .A2(_15197_),
    .A3(_15254_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24684_ (.A1(_00699_),
    .A2(_15258_),
    .A3(_00591_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24685_ (.A1(_15386_),
    .A2(_15383_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24686_ (.A1(_15345_),
    .A2(_15197_),
    .A3(_15266_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24687_ (.A1(_00701_),
    .A2(_00702_),
    .A3(_15272_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24688_ (.A1(_00703_),
    .A2(_15173_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24689_ (.A1(_00700_),
    .A2(_00704_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24690_ (.A1(_00705_),
    .A2(_15191_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24691_ (.A1(_15254_),
    .A2(_00559_),
    .B(_15427_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24692_ (.A1(_00605_),
    .A2(_00707_),
    .B(_15217_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24693_ (.A1(_15531_),
    .A2(_15322_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24694_ (.A1(_15884_),
    .A2(_15893_),
    .B(_15215_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24695_ (.A1(_00709_),
    .A2(_15229_),
    .A3(_00710_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24696_ (.A1(_00708_),
    .A2(_00711_),
    .B(_15340_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24697_ (.A1(_00706_),
    .A2(_00712_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24698_ (.A1(_15330_),
    .A2(_15404_),
    .A3(_15175_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24699_ (.A1(_00714_),
    .A2(_15394_),
    .A3(_15492_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24700_ (.A1(_15330_),
    .A2(_15259_),
    .A3(_15350_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24701_ (.A1(_00611_),
    .A2(_15376_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24702_ (.A1(_00716_),
    .A2(_00717_),
    .A3(_15229_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24703_ (.A1(_00715_),
    .A2(_00718_),
    .A3(_15278_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24704_ (.A1(_15322_),
    .A2(_15398_),
    .A3(_15427_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24705_ (.A1(_15303_),
    .A2(_15252_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24706_ (.A1(_00720_),
    .A2(_00721_),
    .B(_15261_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24707_ (.A1(_15416_),
    .A2(_00563_),
    .B(_15410_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24708_ (.A1(net1051),
    .A2(_15223_),
    .A3(_15245_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24709_ (.A1(_00723_),
    .A2(_00724_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24710_ (.A1(_00722_),
    .A2(_00725_),
    .B(_15239_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24711_ (.A1(_00719_),
    .A2(_00726_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24712_ (.A1(_00713_),
    .A2(_15288_),
    .A3(_00727_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24713_ (.I(_15275_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24714_ (.A1(_00589_),
    .A2(_00729_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24715_ (.A1(_00730_),
    .A2(_15313_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24716_ (.A1(_15467_),
    .A2(_15173_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24717_ (.A1(_00731_),
    .A2(_00732_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24718_ (.A1(_00733_),
    .A2(_15191_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24719_ (.A1(_15406_),
    .A2(_15376_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24720_ (.A1(_00735_),
    .A2(_15324_),
    .A3(_15362_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24721_ (.I(_15885_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24722_ (.A1(_00737_),
    .A2(_15223_),
    .B(_15410_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24723_ (.A1(_00738_),
    .A2(_00675_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24724_ (.A1(_00736_),
    .A2(_00739_),
    .A3(_15262_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24725_ (.A1(_00734_),
    .A2(_15280_),
    .A3(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24726_ (.A1(_15883_),
    .A2(_15881_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24727_ (.A1(_00581_),
    .A2(_00742_),
    .B(_15349_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24728_ (.A1(_15320_),
    .A2(_15427_),
    .A3(_15245_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24729_ (.A1(_00743_),
    .A2(_00744_),
    .A3(_15324_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24730_ (.A1(net10),
    .A2(_15214_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24731_ (.A1(_00550_),
    .A2(_00746_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24732_ (.A1(_00745_),
    .A2(_00747_),
    .A3(_15262_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24733_ (.A1(_15398_),
    .A2(_15223_),
    .B(_15347_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24734_ (.A1(_00749_),
    .A2(_15335_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24735_ (.A1(_15375_),
    .A2(_15215_),
    .B(_15252_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24736_ (.A1(_00582_),
    .A2(_00751_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24737_ (.A1(_00750_),
    .A2(_00752_),
    .A3(_15353_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24738_ (.A1(_00748_),
    .A2(_15240_),
    .A3(_00753_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24739_ (.A1(_00741_),
    .A2(_00754_),
    .A3(_15287_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24740_ (.A1(_00728_),
    .A2(_00755_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24741_ (.A1(_15255_),
    .A2(_15199_),
    .A3(_15246_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24742_ (.A1(_15386_),
    .A2(net10),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24743_ (.A1(_00756_),
    .A2(_00757_),
    .B(_15262_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24744_ (.A1(_15404_),
    .A2(_15872_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24745_ (.A1(_00709_),
    .A2(_15394_),
    .A3(_00759_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24746_ (.A1(_00758_),
    .A2(_00760_),
    .B(_15280_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _24747_ (.A1(_15299_),
    .A2(_15221_),
    .A3(_15215_),
    .B1(_15519_),
    .B2(_00581_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24748_ (.A1(_00762_),
    .A2(_15486_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _24749_ (.A1(_15268_),
    .A2(_00563_),
    .B1(_15404_),
    .B2(_00581_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24750_ (.A1(_00746_),
    .A2(_15252_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24751_ (.A1(_00764_),
    .A2(_00765_),
    .B(_15217_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24752_ (.A1(_00763_),
    .A2(_00766_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24753_ (.A1(_00761_),
    .A2(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24754_ (.A1(_15291_),
    .A2(_15376_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24755_ (.A1(_15328_),
    .A2(_15450_),
    .B(_15307_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24756_ (.A1(_15515_),
    .A2(_00559_),
    .B(_15215_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24757_ (.A1(_15893_),
    .A2(_15248_),
    .B(_15410_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24758_ (.A1(_00771_),
    .A2(_00772_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _24759_ (.A1(_00769_),
    .A2(_00770_),
    .B(_00773_),
    .C(_15353_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24760_ (.A1(_00593_),
    .A2(_15427_),
    .B(_15410_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24761_ (.A1(_00775_),
    .A2(_15255_),
    .B(_15190_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24762_ (.A1(_15357_),
    .A2(_00765_),
    .A3(_00591_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24763_ (.A1(_00776_),
    .A2(_00777_),
    .B(_15239_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24764_ (.A1(_00774_),
    .A2(_00778_),
    .B(_15287_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24765_ (.A1(_00768_),
    .A2(_00779_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24766_ (.A1(_15367_),
    .A2(_15242_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24767_ (.A1(_15512_),
    .A2(_00781_),
    .A3(_00701_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24768_ (.A1(_15371_),
    .A2(_15313_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24769_ (.A1(_00783_),
    .A2(_00589_),
    .B(_15340_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24770_ (.A1(_00782_),
    .A2(_00784_),
    .B(_15353_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24771_ (.A1(_15315_),
    .A2(_15404_),
    .A3(_15350_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24772_ (.A1(_00786_),
    .A2(_15229_),
    .A3(_15500_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24773_ (.A1(_15215_),
    .A2(net1221),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _24774_ (.A1(_00633_),
    .A2(_15404_),
    .B(_15307_),
    .C(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24775_ (.A1(_00787_),
    .A2(_00789_),
    .A3(_15280_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24776_ (.A1(_00785_),
    .A2(_00790_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24777_ (.A1(_15291_),
    .A2(_15345_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24778_ (.A1(_00562_),
    .A2(_00792_),
    .A3(_15324_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24779_ (.A1(_15507_),
    .A2(_15358_),
    .A3(_00702_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24780_ (.A1(_00793_),
    .A2(_00794_),
    .A3(_15240_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24781_ (.A1(_15300_),
    .A2(_15199_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24782_ (.A1(_00796_),
    .A2(_15384_),
    .B(_15239_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24783_ (.A1(_15242_),
    .A2(_15223_),
    .B(_15347_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24784_ (.A1(_15315_),
    .A2(_15349_),
    .A3(_15376_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24785_ (.A1(_00798_),
    .A2(_00799_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24786_ (.A1(_00797_),
    .A2(_00800_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24787_ (.A1(_00795_),
    .A2(_00801_),
    .A3(_15191_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24788_ (.A1(_00802_),
    .A2(_00791_),
    .A3(_15287_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24789_ (.A1(_00780_),
    .A2(_00803_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _24790_ (.I(\sa21_sub[7] ),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24791_ (.A1(_12815_),
    .A2(_00804_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24792_ (.A1(\sa21_sub[0] ),
    .A2(\sa21_sub[7] ),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24793_ (.A1(_00806_),
    .A2(_00805_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _24794_ (.A1(_00807_),
    .A2(_12770_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24795_ (.A1(_00804_),
    .A2(\sa21_sub[0] ),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24796_ (.A1(_12815_),
    .A2(\sa21_sub[7] ),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24797_ (.A1(_00810_),
    .A2(_00809_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24798_ (.A1(_00811_),
    .A2(_12777_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24799_ (.A1(_00812_),
    .A2(_00808_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24800_ (.A1(_12785_),
    .A2(net531),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24801_ (.A1(_12789_),
    .A2(_12830_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24802_ (.A1(_00814_),
    .A2(_00815_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24803_ (.A1(_00816_),
    .A2(_00813_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24804_ (.A1(_12777_),
    .A2(_00811_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24805_ (.A1(_12770_),
    .A2(_00807_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24806_ (.A1(_00818_),
    .A2(_00819_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24807_ (.A1(_12785_),
    .A2(_12830_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24808_ (.A1(_12789_),
    .A2(net738),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24809_ (.A1(_00822_),
    .A2(_00821_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24810_ (.A1(_00823_),
    .A2(_00820_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24811_ (.A1(_00817_),
    .A2(_00824_),
    .A3(_10522_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24812_ (.A1(_10525_),
    .A2(\text_in_r[17] ),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24813_ (.A1(_00825_),
    .A2(_00826_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24814_ (.I(\u0.tmp_w[17] ),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24815_ (.A1(_00828_),
    .A2(net1268),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24816_ (.A1(net527),
    .A2(\u0.tmp_w[17] ),
    .A3(_00826_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24817_ (.A1(_00829_),
    .A2(_00830_),
    .ZN(_15903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24818_ (.A1(_12783_),
    .A2(net746),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24819_ (.A1(_12811_),
    .A2(_12781_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24820_ (.A1(_00831_),
    .A2(_00832_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24821_ (.A1(_00833_),
    .A2(net727),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24822_ (.A1(_00831_),
    .A2(_00832_),
    .A3(_12762_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24823_ (.A1(_00834_),
    .A2(_00835_),
    .A3(net993),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24824_ (.A1(net715),
    .A2(_12781_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24825_ (.I(_00837_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24826_ (.A1(\sa03_sr[0] ),
    .A2(_12781_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24827_ (.A1(_00838_),
    .A2(_00839_),
    .B(net746),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24828_ (.A1(_12762_),
    .A2(net931),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24829_ (.A1(_00841_),
    .A2(_12811_),
    .A3(_00837_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24830_ (.A1(_00840_),
    .A2(_00842_),
    .A3(net1227),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24831_ (.A1(_00836_),
    .A2(_00843_),
    .B(_10586_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24832_ (.I(\text_in_r[16] ),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24833_ (.A1(_00845_),
    .A2(_10482_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24834_ (.A1(_00844_),
    .A2(_00846_),
    .B(\u0.tmp_w[16] ),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24835_ (.A1(_00836_),
    .A2(_00843_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24836_ (.A1(_00848_),
    .A2(_10479_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24837_ (.I(\u0.tmp_w[16] ),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24838_ (.I(_00846_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24839_ (.A1(_00849_),
    .A2(_00850_),
    .A3(_00851_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24840_ (.A1(_00852_),
    .A2(_00847_),
    .ZN(_15906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24841_ (.A1(_12836_),
    .A2(\sa32_sub[2] ),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24842_ (.A1(_12836_),
    .A2(\sa32_sub[2] ),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24843_ (.A1(_00853_),
    .A2(_00854_),
    .B(\sa03_sr[2] ),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24844_ (.A1(_12834_),
    .A2(_12839_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24845_ (.A1(_12836_),
    .A2(\sa32_sub[2] ),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24846_ (.A1(_00856_),
    .A2(_12864_),
    .A3(_00857_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24847_ (.A1(_00855_),
    .A2(_00858_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24848_ (.A1(net735),
    .A2(net529),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24849_ (.I(_00860_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24850_ (.A1(_00859_),
    .A2(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24851_ (.A1(_00855_),
    .A2(_00858_),
    .A3(_00860_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24852_ (.A1(_00862_),
    .A2(_00863_),
    .B(_10381_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24853_ (.I(\text_in_r[18] ),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24854_ (.A1(_00865_),
    .A2(net596),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24855_ (.I(\u0.tmp_w[18] ),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _24856_ (.A1(_00864_),
    .A2(_00866_),
    .B(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24857_ (.A1(_00862_),
    .A2(_00863_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24858_ (.A1(_00869_),
    .A2(_10402_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24859_ (.I(_00866_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24860_ (.A1(_00870_),
    .A2(\u0.tmp_w[18] ),
    .A3(_00871_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24861_ (.A1(_00868_),
    .A2(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24862_ (.I(_00873_),
    .Z(_15922_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _24863_ (.A1(_00844_),
    .A2(_00846_),
    .B(_00850_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24864_ (.A1(_00849_),
    .A2(\u0.tmp_w[16] ),
    .A3(_00851_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24865_ (.A1(_00874_),
    .A2(_00875_),
    .ZN(_15897_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _24866_ (.A1(_00864_),
    .A2(_00866_),
    .B(\u0.tmp_w[18] ),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24867_ (.A1(_00870_),
    .A2(_00867_),
    .A3(_00871_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24868_ (.A1(_00876_),
    .A2(_00877_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24869_ (.I(_00878_),
    .Z(_15915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24870_ (.A1(_12834_),
    .A2(_00804_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24871_ (.A1(_12836_),
    .A2(net745),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24872_ (.A1(_00880_),
    .A2(_00879_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24873_ (.A1(_12872_),
    .A2(net755),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24874_ (.A1(_00804_),
    .A2(_12836_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24875_ (.A1(_12834_),
    .A2(net50),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24876_ (.A1(_00883_),
    .A2(_00884_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24877_ (.A1(_12879_),
    .A2(_00885_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24878_ (.A1(_00882_),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24879_ (.I(_00887_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24880_ (.A1(_12898_),
    .A2(\sa03_sr[3] ),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24881_ (.I(\sa03_sr[3] ),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24882_ (.A1(_12896_),
    .A2(_00890_),
    .A3(_12897_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24883_ (.A1(_00889_),
    .A2(_00891_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24884_ (.I(_00892_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24885_ (.A1(_00888_),
    .A2(_00893_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24886_ (.A1(_00887_),
    .A2(_00892_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24887_ (.A1(_00894_),
    .A2(_10489_),
    .A3(_00895_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24888_ (.A1(_12193_),
    .A2(\text_in_r[19] ),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24889_ (.A1(_00896_),
    .A2(_00897_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24890_ (.A1(_00898_),
    .A2(\u0.tmp_w[19] ),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24891_ (.I(\u0.tmp_w[19] ),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24892_ (.A1(_00896_),
    .A2(_00900_),
    .A3(_00897_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24893_ (.A1(_00899_),
    .A2(_00901_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24894_ (.I(_00902_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24895_ (.I(_00903_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24896_ (.I(_15900_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24897_ (.A1(net1222),
    .A2(net1226),
    .A3(_00905_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24898_ (.I(net1223),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24899_ (.A1(_15922_),
    .A2(net1232),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _24900_ (.I(_00878_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24901_ (.A1(_00909_),
    .A2(_15909_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24902_ (.A1(_00908_),
    .A2(_00910_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24903_ (.I(_00902_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24904_ (.A1(_00911_),
    .A2(_00912_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24905_ (.A1(_12870_),
    .A2(_00804_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24906_ (.A1(\sa21_sub[3] ),
    .A2(net50),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24907_ (.A1(_00914_),
    .A2(_00915_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24908_ (.I(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24909_ (.I(\sa32_sub[4] ),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24910_ (.A1(_12928_),
    .A2(_00918_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24911_ (.A1(\sa21_sub[4] ),
    .A2(\sa32_sub[4] ),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24912_ (.A1(_00919_),
    .A2(_00920_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24913_ (.A1(_00917_),
    .A2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24914_ (.I(_00921_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24915_ (.A1(_00923_),
    .A2(_00916_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24916_ (.A1(_00922_),
    .A2(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24917_ (.I(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24918_ (.A1(\sa03_sr[4] ),
    .A2(_12889_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24919_ (.A1(_00926_),
    .A2(_00927_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24920_ (.A1(_12889_),
    .A2(\sa03_sr[4] ),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24921_ (.A1(_12889_),
    .A2(\sa03_sr[4] ),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24922_ (.A1(_00929_),
    .A2(_00930_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24923_ (.A1(_00925_),
    .A2(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24924_ (.A1(_00928_),
    .A2(_00932_),
    .A3(_10479_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24925_ (.A1(_10483_),
    .A2(\text_in_r[20] ),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24926_ (.A1(_00933_),
    .A2(_00934_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24927_ (.A1(_00935_),
    .A2(\u0.tmp_w[20] ),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24928_ (.I(\u0.tmp_w[20] ),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24929_ (.A1(_00933_),
    .A2(_00937_),
    .A3(_00934_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24930_ (.A1(_00936_),
    .A2(_00938_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24931_ (.I(_00939_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24932_ (.I(_00940_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _24933_ (.A1(_00904_),
    .A2(net1011),
    .B(_00913_),
    .C(_00941_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24934_ (.A1(net1269),
    .A2(_15906_),
    .A3(_15915_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24935_ (.A1(_00898_),
    .A2(_00900_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24936_ (.A1(_00896_),
    .A2(\u0.tmp_w[19] ),
    .A3(_00897_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24937_ (.A1(_00944_),
    .A2(_00945_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24938_ (.I(_00946_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24939_ (.A1(net941),
    .A2(net484),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24940_ (.A1(_00943_),
    .A2(_00947_),
    .A3(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24941_ (.I(_00908_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _24942_ (.I(_00902_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24943_ (.I(_00951_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24944_ (.I(_00940_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24945_ (.A1(_00950_),
    .A2(_00952_),
    .B(_00953_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24946_ (.A1(_00949_),
    .A2(_00954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24947_ (.I(\sa03_sr[5] ),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24948_ (.A1(_00956_),
    .A2(_12958_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24949_ (.A1(\sa10_sub[4] ),
    .A2(\sa21_sub[4] ),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24950_ (.I(_00958_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24951_ (.A1(_00957_),
    .A2(_00959_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24952_ (.A1(_00957_),
    .A2(_00959_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24953_ (.A1(_00960_),
    .A2(_00961_),
    .A3(_11348_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24954_ (.A1(_10587_),
    .A2(\text_in_r[21] ),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24955_ (.A1(_00962_),
    .A2(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24956_ (.A1(_00964_),
    .A2(\u0.tmp_w[21] ),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24957_ (.I(\u0.tmp_w[21] ),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24958_ (.A1(_00962_),
    .A2(_00966_),
    .A3(_00963_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24959_ (.A1(_00965_),
    .A2(_00967_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24960_ (.I(_00968_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24961_ (.A1(_00942_),
    .A2(_00955_),
    .A3(_00969_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24962_ (.A1(_00909_),
    .A2(_15901_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24963_ (.I(_00971_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24964_ (.I(_15899_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24965_ (.A1(_15922_),
    .A2(_00973_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24966_ (.A1(_00972_),
    .A2(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24967_ (.I(_00903_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24968_ (.A1(_00975_),
    .A2(_00976_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24969_ (.I(_15904_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24970_ (.A1(_00978_),
    .A2(_00909_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _24971_ (.I(_00946_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24972_ (.A1(net1094),
    .A2(_00979_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24973_ (.I(_00939_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24974_ (.I(_00982_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24975_ (.A1(_00981_),
    .A2(_00983_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24976_ (.I(_00968_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24977_ (.A1(_00977_),
    .A2(_00984_),
    .B(_00985_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24978_ (.A1(_00909_),
    .A2(_15906_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24979_ (.I(_00987_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24980_ (.I(_15907_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24981_ (.A1(_15922_),
    .A2(_00989_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _24982_ (.I(_00946_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _24983_ (.I(_00991_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24984_ (.A1(_00988_),
    .A2(_00990_),
    .B(_00992_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24985_ (.A1(net1269),
    .A2(_15915_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24986_ (.A1(_15900_),
    .A2(net1090),
    .A3(net1224),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24987_ (.A1(_00994_),
    .A2(_00952_),
    .A3(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _24988_ (.I(_00982_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24989_ (.A1(_00993_),
    .A2(_00996_),
    .A3(_00997_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24990_ (.A1(\sa10_sub[5] ),
    .A2(\sa21_sub[5] ),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24991_ (.I(\sa03_sr[6] ),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24992_ (.A1(_01000_),
    .A2(_13007_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24993_ (.A1(_00999_),
    .A2(_01001_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24994_ (.A1(_10587_),
    .A2(\text_in_r[22] ),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24995_ (.A1(_01002_),
    .A2(_10585_),
    .B(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24996_ (.I(\u0.tmp_w[22] ),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24997_ (.A1(_01004_),
    .A2(_01005_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24998_ (.A1(_01004_),
    .A2(_01005_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24999_ (.A1(_01006_),
    .A2(_01007_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25000_ (.I(_01008_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25001_ (.A1(_00986_),
    .A2(_00998_),
    .B(_01009_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25002_ (.A1(_00970_),
    .A2(_01010_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25003_ (.A1(net39),
    .A2(\sa10_sub[6] ),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25004_ (.A1(\sa21_sub[6] ),
    .A2(_01012_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _25005_ (.A1(net50),
    .A2(net54),
    .A3(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _25006_ (.I0(_01014_),
    .I1(\text_in_r[23] ),
    .S(_10587_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _25007_ (.A1(\u0.tmp_w[23] ),
    .A2(_01015_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25008_ (.I(_01016_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _25009_ (.I(_01017_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25010_ (.A1(_15922_),
    .A2(net535),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25011_ (.A1(_00909_),
    .A2(_00973_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25012_ (.A1(_01019_),
    .A2(_01020_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25013_ (.I(_00940_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25014_ (.A1(_01021_),
    .A2(_00947_),
    .B(_01022_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25015_ (.A1(net16),
    .A2(net34),
    .A3(_00909_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25016_ (.A1(net1091),
    .A2(net1225),
    .A3(_00978_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25017_ (.A1(_01024_),
    .A2(_00952_),
    .A3(_01025_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25018_ (.A1(net1091),
    .A2(net1225),
    .A3(_15901_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25019_ (.I(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25020_ (.A1(_01028_),
    .A2(_00952_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25021_ (.A1(_01023_),
    .A2(_01026_),
    .A3(_01029_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25022_ (.I(_00995_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25023_ (.A1(_01031_),
    .A2(_00912_),
    .B(_00982_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25024_ (.A1(_00992_),
    .A2(_15920_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25025_ (.I(_00968_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25026_ (.I(_01034_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25027_ (.A1(_01032_),
    .A2(_01033_),
    .B(_01035_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25028_ (.A1(_01030_),
    .A2(_01036_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25029_ (.A1(_00971_),
    .A2(_00976_),
    .B(_01022_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25030_ (.I(_15909_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25031_ (.A1(net1091),
    .A2(net1224),
    .A3(_01039_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25032_ (.A1(_01040_),
    .A2(_00980_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25033_ (.A1(_01041_),
    .A2(_01024_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25034_ (.I(_00968_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25035_ (.A1(_01038_),
    .A2(_01042_),
    .B(_01043_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25036_ (.A1(net941),
    .A2(_15907_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25037_ (.A1(_01045_),
    .A2(_00951_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25038_ (.A1(_01046_),
    .A2(_01024_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25039_ (.I(_00946_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25040_ (.A1(_00971_),
    .A2(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25041_ (.A1(_01047_),
    .A2(_00941_),
    .A3(_01049_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25042_ (.A1(_01044_),
    .A2(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25043_ (.I(_01008_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25044_ (.A1(_01037_),
    .A2(_01051_),
    .A3(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25045_ (.A1(_01011_),
    .A2(_01018_),
    .A3(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25046_ (.A1(_00948_),
    .A2(_00951_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25047_ (.A1(_01055_),
    .A2(_00982_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25048_ (.A1(net940),
    .A2(net34),
    .A3(net497),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25049_ (.A1(_00981_),
    .A2(net498),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25050_ (.A1(_01056_),
    .A2(_01058_),
    .B(_01043_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25051_ (.A1(_00909_),
    .A2(net34),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25052_ (.A1(net498),
    .A2(_00952_),
    .A3(_01060_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25053_ (.A1(_00906_),
    .A2(net1094),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25054_ (.I(_15913_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25055_ (.A1(_01063_),
    .A2(net941),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25056_ (.A1(net1095),
    .A2(_01062_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25057_ (.I(_00940_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25058_ (.A1(_01061_),
    .A2(_01066_),
    .A3(_01065_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25059_ (.A1(_01059_),
    .A2(_01067_),
    .B(_01009_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25060_ (.A1(_01057_),
    .A2(_00903_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25061_ (.A1(\u0.tmp_w[17] ),
    .A2(_00827_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25062_ (.A1(net502),
    .A2(_00828_),
    .A3(_00826_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25063_ (.A1(_01071_),
    .A2(_01070_),
    .ZN(_15898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25064_ (.A1(net21),
    .A2(_00909_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25065_ (.I(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25066_ (.A1(_01069_),
    .A2(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25067_ (.A1(_00948_),
    .A2(_01048_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25068_ (.A1(_00909_),
    .A2(_01063_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25069_ (.I(_00939_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25070_ (.A1(_01075_),
    .A2(_01076_),
    .B(_01077_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25071_ (.A1(_01074_),
    .A2(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25072_ (.A1(net16),
    .A2(_00909_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25073_ (.A1(_01080_),
    .A2(_00971_),
    .B(_00952_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25074_ (.I(_00982_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25075_ (.A1(_00949_),
    .A2(_01081_),
    .A3(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25076_ (.I(_00968_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25077_ (.A1(_01079_),
    .A2(_01083_),
    .A3(_01084_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25078_ (.A1(_01085_),
    .A2(_01068_),
    .B(_01018_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25079_ (.I(_01020_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25080_ (.I(_00903_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25081_ (.A1(_00990_),
    .A2(_01087_),
    .B(_01088_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25082_ (.A1(_15922_),
    .A2(_15899_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25083_ (.A1(_01062_),
    .A2(_01090_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25084_ (.A1(_01089_),
    .A2(_01091_),
    .B(_01066_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25085_ (.A1(_15922_),
    .A2(_00905_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25086_ (.A1(_01093_),
    .A2(_00980_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25087_ (.A1(_01094_),
    .A2(_00982_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25088_ (.A1(net1222),
    .A2(net1226),
    .A3(_15900_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25089_ (.A1(_01096_),
    .A2(_00951_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25090_ (.I(_01097_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25091_ (.A1(net499),
    .A2(net941),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25092_ (.A1(_01098_),
    .A2(_01099_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25093_ (.A1(_01095_),
    .A2(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25094_ (.A1(_01092_),
    .A2(_01101_),
    .B(_00969_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25095_ (.A1(_00987_),
    .A2(_00951_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25096_ (.A1(net21),
    .A2(net34),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25097_ (.A1(_01103_),
    .A2(_01104_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25098_ (.A1(net496),
    .A2(net485),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25099_ (.A1(net1266),
    .A2(_01048_),
    .A3(_01019_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25100_ (.A1(_01105_),
    .A2(_00941_),
    .A3(_01107_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25101_ (.A1(net1097),
    .A2(_00951_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25102_ (.A1(net16),
    .A2(net536),
    .A3(_15922_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25103_ (.A1(_01109_),
    .A2(_01110_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25104_ (.A1(_15915_),
    .A2(_00989_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25105_ (.A1(_00974_),
    .A2(_01112_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25106_ (.A1(_01113_),
    .A2(_00992_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25107_ (.A1(_01111_),
    .A2(_01114_),
    .A3(_00983_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25108_ (.I(_01034_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25109_ (.A1(_01108_),
    .A2(_01115_),
    .A3(_01116_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25110_ (.A1(_01102_),
    .A2(_01117_),
    .A3(_01052_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25111_ (.A1(_01118_),
    .A2(_01086_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25112_ (.A1(_01119_),
    .A2(_01054_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25113_ (.A1(net1089),
    .A2(net941),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25114_ (.A1(_00981_),
    .A2(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25115_ (.A1(_00987_),
    .A2(_01090_),
    .A3(_01088_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25116_ (.A1(_01121_),
    .A2(_01082_),
    .A3(_01122_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25117_ (.A1(_00971_),
    .A2(_01088_),
    .B(_01077_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25118_ (.I(_01019_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25119_ (.A1(_01125_),
    .A2(_01088_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25120_ (.A1(_01020_),
    .A2(_00995_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _25121_ (.I(_00991_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25122_ (.A1(_01127_),
    .A2(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25123_ (.A1(_01124_),
    .A2(_01126_),
    .A3(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25124_ (.A1(_01123_),
    .A2(_01130_),
    .A3(_01116_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25125_ (.A1(_01110_),
    .A2(_00991_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25126_ (.I(_01096_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25127_ (.A1(_01132_),
    .A2(_01133_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25128_ (.A1(_01076_),
    .A2(_00903_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25129_ (.I(_15901_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25130_ (.A1(_15922_),
    .A2(_01136_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25131_ (.A1(_01135_),
    .A2(_01137_),
    .B(_01077_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25132_ (.A1(_01134_),
    .A2(_01138_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25133_ (.I(_01055_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25134_ (.A1(_01140_),
    .A2(_00943_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25135_ (.A1(_01062_),
    .A2(_01022_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25136_ (.A1(_01141_),
    .A2(_01142_),
    .B(_01035_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25137_ (.A1(_01139_),
    .A2(_01143_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25138_ (.A1(_01144_),
    .A2(_01131_),
    .B(_01052_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25139_ (.A1(_01103_),
    .A2(_01099_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25140_ (.A1(_01146_),
    .A2(_01121_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25141_ (.A1(_01147_),
    .A2(_01084_),
    .B(_00997_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25142_ (.A1(_00943_),
    .A2(_01057_),
    .A3(_00992_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25143_ (.A1(_01060_),
    .A2(_01090_),
    .A3(_01088_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25144_ (.A1(_01149_),
    .A2(_01150_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25145_ (.A1(_01151_),
    .A2(_01116_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25146_ (.I(_15923_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25147_ (.A1(_01048_),
    .A2(_01153_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25148_ (.A1(_01154_),
    .A2(_00968_),
    .B(_01022_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25149_ (.A1(_01046_),
    .A2(_00943_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25150_ (.A1(_01155_),
    .A2(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25151_ (.A1(_01157_),
    .A2(_01009_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25152_ (.A1(_01148_),
    .A2(_01152_),
    .B(_01158_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25153_ (.A1(_01145_),
    .A2(_01159_),
    .B(_01017_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25154_ (.A1(_15915_),
    .A2(net1232),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25155_ (.I(_00940_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25156_ (.A1(_01161_),
    .A2(_00904_),
    .B(_01162_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25157_ (.A1(_01134_),
    .A2(_01163_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25158_ (.A1(_01064_),
    .A2(_00991_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25159_ (.A1(_01165_),
    .A2(_01073_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25160_ (.A1(net16),
    .A2(net536),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25161_ (.A1(_01167_),
    .A2(_15915_),
    .A3(_01088_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25162_ (.A1(_01166_),
    .A2(_01168_),
    .A3(_00941_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25163_ (.A1(_01164_),
    .A2(_01169_),
    .A3(_01116_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25164_ (.A1(_00950_),
    .A2(net1011),
    .B(_01128_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25165_ (.A1(_01021_),
    .A2(_00904_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25166_ (.A1(_01171_),
    .A2(_01172_),
    .A3(_00941_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25167_ (.A1(_01167_),
    .A2(_01060_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25168_ (.A1(_01174_),
    .A2(_00992_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25169_ (.A1(_00995_),
    .A2(_00951_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25170_ (.A1(_01176_),
    .A2(_01060_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25171_ (.A1(_01175_),
    .A2(_01177_),
    .A3(_00983_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25172_ (.A1(_01173_),
    .A2(_01178_),
    .A3(_01084_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25173_ (.I(_01008_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25174_ (.I(_01180_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25175_ (.A1(_01170_),
    .A2(_01179_),
    .A3(_01181_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25176_ (.A1(_01094_),
    .A2(_01076_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25177_ (.A1(_01026_),
    .A2(_01183_),
    .A3(_01082_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25178_ (.A1(_00950_),
    .A2(_00952_),
    .B(_00982_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25179_ (.A1(_01099_),
    .A2(_00980_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25180_ (.A1(_01185_),
    .A2(net1229),
    .A3(_01186_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25181_ (.A1(_01184_),
    .A2(_01084_),
    .A3(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25182_ (.A1(_00979_),
    .A2(_00903_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25183_ (.A1(_01189_),
    .A2(_01125_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25184_ (.A1(_01062_),
    .A2(_00948_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25185_ (.A1(_01190_),
    .A2(_01066_),
    .A3(_01191_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25186_ (.A1(_00994_),
    .A2(_01104_),
    .A3(_00952_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25187_ (.A1(_00991_),
    .A2(_15922_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25188_ (.A1(_01194_),
    .A2(net1266),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25189_ (.A1(_01193_),
    .A2(_01195_),
    .A3(_00983_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25190_ (.A1(_01192_),
    .A2(_01196_),
    .A3(_01035_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25191_ (.A1(_01188_),
    .A2(_01197_),
    .A3(_01052_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25192_ (.A1(_01182_),
    .A2(_01198_),
    .A3(_01018_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25193_ (.A1(_01160_),
    .A2(_01199_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25194_ (.A1(_01060_),
    .A2(_01025_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25195_ (.A1(_01200_),
    .A2(_00947_),
    .A3(_01072_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25196_ (.A1(_01201_),
    .A2(_00996_),
    .A3(_00983_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25197_ (.A1(_00994_),
    .A2(net1266),
    .A3(_01048_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25198_ (.A1(_00979_),
    .A2(_01064_),
    .A3(_00912_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25199_ (.A1(_01203_),
    .A2(_01204_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25200_ (.A1(_01205_),
    .A2(_01162_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25201_ (.A1(_01202_),
    .A2(_01206_),
    .A3(_01084_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25202_ (.A1(_01057_),
    .A2(_00912_),
    .B(_00940_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25203_ (.A1(_01110_),
    .A2(_00947_),
    .A3(_01076_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25204_ (.A1(_01208_),
    .A2(_01209_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25205_ (.A1(_01097_),
    .A2(_01080_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25206_ (.A1(_01027_),
    .A2(net1094),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25207_ (.A1(_01212_),
    .A2(_00988_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25208_ (.A1(_01211_),
    .A2(_01213_),
    .B(_00953_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25209_ (.A1(_01210_),
    .A2(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25210_ (.A1(_01215_),
    .A2(_01035_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25211_ (.A1(_01207_),
    .A2(_01216_),
    .A3(_01052_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25212_ (.A1(net1091),
    .A2(net1225),
    .A3(_15913_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25213_ (.A1(_00987_),
    .A2(_01218_),
    .A3(_00951_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25214_ (.A1(_01219_),
    .A2(_00940_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25215_ (.A1(_00910_),
    .A2(net1092),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25216_ (.A1(_01221_),
    .A2(_01080_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25217_ (.A1(_01220_),
    .A2(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25218_ (.A1(_01060_),
    .A2(_01040_),
    .A3(_00903_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25219_ (.A1(_00906_),
    .A2(_00995_),
    .A3(net1092),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25220_ (.A1(_01224_),
    .A2(_01225_),
    .B(_00953_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25221_ (.A1(_01223_),
    .A2(_01226_),
    .B(_01034_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25222_ (.A1(_01072_),
    .A2(_01048_),
    .A3(_01025_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25223_ (.A1(_00913_),
    .A2(_01228_),
    .A3(_01077_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25224_ (.I(_01218_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25225_ (.A1(_01230_),
    .A2(_00903_),
    .B(_00982_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25226_ (.I(_00910_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25227_ (.A1(_01232_),
    .A2(_00912_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25228_ (.A1(_01060_),
    .A2(_01025_),
    .A3(net1092),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25229_ (.A1(_01231_),
    .A2(_01233_),
    .A3(_01234_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25230_ (.A1(_01229_),
    .A2(_01235_),
    .A3(_01043_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25231_ (.A1(_01227_),
    .A2(_01236_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25232_ (.A1(_01237_),
    .A2(_01181_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25233_ (.A1(_01217_),
    .A2(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25234_ (.A1(_01239_),
    .A2(_01017_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25235_ (.I(_00940_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25236_ (.A1(_00951_),
    .A2(_15918_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25237_ (.A1(_01242_),
    .A2(_01069_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25238_ (.A1(_15927_),
    .A2(_01088_),
    .B(_01077_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25239_ (.A1(_01203_),
    .A2(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25240_ (.A1(_01241_),
    .A2(_01243_),
    .B(_01245_),
    .C(_01084_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25241_ (.A1(_01087_),
    .A2(_00912_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25242_ (.A1(_01247_),
    .A2(_01077_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25243_ (.A1(_01062_),
    .A2(_01025_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25244_ (.A1(_01249_),
    .A2(_01248_),
    .B(_00985_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25245_ (.A1(_00980_),
    .A2(_15915_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25246_ (.I(_01251_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25247_ (.A1(_01136_),
    .A2(_00978_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25248_ (.I(_01253_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25249_ (.A1(_01252_),
    .A2(_01254_),
    .B(_01077_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25250_ (.A1(_01120_),
    .A2(_00948_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25251_ (.A1(_01256_),
    .A2(net1092),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25252_ (.A1(_01255_),
    .A2(_01156_),
    .A3(_01257_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25253_ (.A1(_01250_),
    .A2(_01258_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25254_ (.A1(_01246_),
    .A2(_01259_),
    .A3(_01052_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25255_ (.A1(_15920_),
    .A2(_00976_),
    .B(_01022_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25256_ (.A1(_01094_),
    .A2(_01024_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25257_ (.A1(_01261_),
    .A2(_01262_),
    .B(_01043_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25258_ (.A1(_01120_),
    .A2(net1094),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25259_ (.A1(_01264_),
    .A2(_01060_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25260_ (.A1(_01265_),
    .A2(_00941_),
    .A3(_00996_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25261_ (.A1(_01263_),
    .A2(_01266_),
    .B(_01009_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25262_ (.A1(_01104_),
    .A2(net1094),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25263_ (.A1(_01268_),
    .A2(_00994_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25264_ (.A1(_00904_),
    .A2(_01153_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25265_ (.A1(_01269_),
    .A2(_00997_),
    .A3(_01270_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25266_ (.A1(_00994_),
    .A2(_00974_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25267_ (.A1(_01272_),
    .A2(_01128_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25268_ (.A1(_01112_),
    .A2(_00947_),
    .A3(net1271),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25269_ (.A1(_01273_),
    .A2(_01274_),
    .B(_01066_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25270_ (.A1(_01271_),
    .A2(_01275_),
    .A3(_01084_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25271_ (.A1(_01267_),
    .A2(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25272_ (.A1(_01260_),
    .A2(_01277_),
    .A3(_01018_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25273_ (.A1(_01240_),
    .A2(_01278_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25274_ (.A1(_01046_),
    .A2(_00994_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25275_ (.I(_01093_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25276_ (.A1(_01280_),
    .A2(_01048_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25277_ (.A1(_01279_),
    .A2(_01281_),
    .B(_00968_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25278_ (.A1(_00907_),
    .A2(_00951_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _25279_ (.A1(_01283_),
    .A2(_01034_),
    .B1(_00992_),
    .B2(_00971_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25280_ (.A1(_01282_),
    .A2(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25281_ (.A1(_01285_),
    .A2(_01241_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25282_ (.A1(_01232_),
    .A2(_01128_),
    .B(_00968_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25283_ (.A1(_01224_),
    .A2(_01287_),
    .B(_01066_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25284_ (.A1(_01140_),
    .A2(_00906_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25285_ (.A1(_15915_),
    .A2(_01253_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25286_ (.A1(_01290_),
    .A2(net1092),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25287_ (.A1(_01291_),
    .A2(net1096),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25288_ (.A1(_01289_),
    .A2(_01292_),
    .A3(_00985_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25289_ (.A1(_01288_),
    .A2(_01293_),
    .B(_01181_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25290_ (.A1(_01286_),
    .A2(_01294_),
    .B(_01018_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25291_ (.A1(_01291_),
    .A2(_01040_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25292_ (.A1(_01156_),
    .A2(_01296_),
    .B(_00941_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25293_ (.I(_01220_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25294_ (.A1(_01297_),
    .A2(_01298_),
    .B(_00969_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25295_ (.A1(_01023_),
    .A2(_01193_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25296_ (.A1(net1233),
    .A2(net1095),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25297_ (.A1(_00948_),
    .A2(_00910_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25298_ (.A1(_01302_),
    .A2(_00947_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25299_ (.A1(_01301_),
    .A2(_01303_),
    .A3(_00941_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25300_ (.A1(_01300_),
    .A2(_01304_),
    .A3(_01116_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25301_ (.A1(_01299_),
    .A2(_01305_),
    .A3(_01181_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25302_ (.A1(_01295_),
    .A2(_01306_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25303_ (.A1(_01106_),
    .A2(_00987_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25304_ (.A1(_01308_),
    .A2(_00982_),
    .A3(_01251_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25305_ (.A1(_01309_),
    .A2(_01009_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25306_ (.A1(_01098_),
    .A2(_01040_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25307_ (.A1(_01166_),
    .A2(_01311_),
    .A3(_01066_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25308_ (.A1(_01310_),
    .A2(_01312_),
    .B(_01116_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _25309_ (.A1(_01103_),
    .A2(net1267),
    .B1(_01120_),
    .B2(_01062_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25310_ (.A1(_01314_),
    .A2(_00997_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25311_ (.A1(_01120_),
    .A2(_00976_),
    .A3(_01060_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25312_ (.A1(_01095_),
    .A2(_01316_),
    .B(_01180_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25313_ (.A1(_01315_),
    .A2(_01317_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25314_ (.A1(_01318_),
    .A2(_01313_),
    .B(_01017_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25315_ (.A1(_01025_),
    .A2(_00980_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25316_ (.A1(_01320_),
    .A2(_01076_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _25317_ (.A1(_01321_),
    .A2(_01162_),
    .A3(_01211_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25318_ (.A1(_01019_),
    .A2(_01112_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25319_ (.A1(_01323_),
    .A2(_00947_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25320_ (.A1(_01252_),
    .A2(_00973_),
    .B(_00982_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25321_ (.I(_01281_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25322_ (.A1(_01324_),
    .A2(_01325_),
    .A3(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25323_ (.A1(_01322_),
    .A2(_01327_),
    .A3(_01009_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25324_ (.A1(_01264_),
    .A2(_01323_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25325_ (.A1(_01167_),
    .A2(_15915_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25326_ (.A1(_01330_),
    .A2(_01176_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25327_ (.A1(_01329_),
    .A2(_00983_),
    .A3(_01331_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25328_ (.I(_00990_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25329_ (.A1(_01109_),
    .A2(_01333_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25330_ (.A1(_01334_),
    .A2(_01107_),
    .A3(_01162_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25331_ (.A1(_01332_),
    .A2(_01335_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25332_ (.A1(_01336_),
    .A2(_01181_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25333_ (.A1(_01328_),
    .A2(_01116_),
    .A3(_01337_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25334_ (.A1(_01319_),
    .A2(_01338_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25335_ (.A1(_01307_),
    .A2(_01339_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25336_ (.A1(_01269_),
    .A2(_01077_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25337_ (.A1(_01340_),
    .A2(_01146_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25338_ (.A1(_01106_),
    .A2(_01120_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25339_ (.A1(_01342_),
    .A2(_00904_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25340_ (.A1(_01272_),
    .A2(_00992_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25341_ (.A1(_01343_),
    .A2(_01344_),
    .A3(_01241_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25342_ (.A1(_01341_),
    .A2(_00969_),
    .A3(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25343_ (.I(_01186_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25344_ (.A1(_01347_),
    .A2(_01060_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25345_ (.A1(_01348_),
    .A2(_00997_),
    .A3(_01150_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25346_ (.A1(_00972_),
    .A2(_00953_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25347_ (.I(_01041_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25348_ (.A1(_01350_),
    .A2(_01351_),
    .B(_01043_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25349_ (.A1(_01349_),
    .A2(_01352_),
    .B(_01009_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25350_ (.A1(_01346_),
    .A2(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25351_ (.A1(_01048_),
    .A2(_01031_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25352_ (.A1(_01355_),
    .A2(_00910_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25353_ (.A1(_01356_),
    .A2(_01185_),
    .B(_00985_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25354_ (.A1(_01135_),
    .A2(_01093_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25355_ (.A1(_01358_),
    .A2(_01042_),
    .A3(_01082_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25356_ (.A1(_01359_),
    .A2(_01357_),
    .B(_01181_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25357_ (.A1(_01264_),
    .A2(_01024_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25358_ (.A1(_01361_),
    .A2(_01241_),
    .A3(_01204_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25359_ (.A1(_01099_),
    .A2(_01020_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25360_ (.A1(_01363_),
    .A2(_00992_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25361_ (.A1(_01026_),
    .A2(_00997_),
    .A3(_01364_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25362_ (.A1(_01362_),
    .A2(_01365_),
    .A3(_00969_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25363_ (.A1(_01360_),
    .A2(_01366_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25364_ (.A1(_01367_),
    .A2(_01354_),
    .A3(_01018_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25365_ (.A1(_01041_),
    .A2(_01072_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25366_ (.A1(_01073_),
    .A2(_00976_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25367_ (.A1(_00988_),
    .A2(_00912_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25368_ (.A1(_01035_),
    .A2(_01370_),
    .A3(_01369_),
    .A4(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25369_ (.A1(_01342_),
    .A2(_01048_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25370_ (.A1(_01041_),
    .A2(_00987_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25371_ (.A1(_01373_),
    .A2(_01374_),
    .A3(_00985_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25372_ (.A1(_01372_),
    .A2(_01375_),
    .A3(_01241_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25373_ (.A1(_00977_),
    .A2(_01107_),
    .A3(_00985_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25374_ (.I(_15911_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25375_ (.A1(_01378_),
    .A2(_01088_),
    .B(_00968_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25376_ (.A1(_00995_),
    .A2(_01128_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25377_ (.A1(_01379_),
    .A2(_01380_),
    .B(_01066_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25378_ (.A1(_01377_),
    .A2(_01381_),
    .B(_01180_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25379_ (.A1(_01376_),
    .A2(_01382_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25380_ (.A1(_01247_),
    .A2(_00953_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25381_ (.A1(_01080_),
    .A2(_00904_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25382_ (.A1(_01384_),
    .A2(_01385_),
    .A3(_01121_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25383_ (.A1(_01103_),
    .A2(_01064_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25384_ (.A1(_01194_),
    .A2(_01162_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25385_ (.A1(_01387_),
    .A2(_01388_),
    .B(_01035_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25386_ (.A1(_01386_),
    .A2(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25387_ (.A1(_01189_),
    .A2(_01031_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25388_ (.A1(_00949_),
    .A2(_01391_),
    .A3(_01082_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25389_ (.A1(_01137_),
    .A2(_00912_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25390_ (.A1(_01393_),
    .A2(_00953_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25391_ (.A1(_01394_),
    .A2(_01132_),
    .B(_01043_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25392_ (.A1(_01392_),
    .A2(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25393_ (.A1(_01390_),
    .A2(_01396_),
    .A3(_01181_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25394_ (.A1(_01383_),
    .A2(_01397_),
    .A3(_01017_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25395_ (.A1(_01368_),
    .A2(_01398_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25396_ (.A1(_01330_),
    .A2(_01333_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25397_ (.A1(_01140_),
    .A2(_01167_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25398_ (.A1(_00904_),
    .A2(_01399_),
    .B(_01400_),
    .C(_01162_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25399_ (.A1(net21),
    .A2(_00947_),
    .B(_00953_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25400_ (.A1(_01373_),
    .A2(_01402_),
    .B(_00968_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25401_ (.A1(_01401_),
    .A2(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25402_ (.A1(_00974_),
    .A2(net1097),
    .B(_00952_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25403_ (.A1(_01230_),
    .A2(_00912_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _25404_ (.A1(_01405_),
    .A2(_01162_),
    .A3(_01406_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25405_ (.A1(_00994_),
    .A2(_00912_),
    .A3(_01137_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25406_ (.A1(_01355_),
    .A2(_00953_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25407_ (.A1(_01408_),
    .A2(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25408_ (.A1(_01407_),
    .A2(_01410_),
    .B(_01084_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25409_ (.A1(_01404_),
    .A2(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25410_ (.A1(_01412_),
    .A2(_01052_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25411_ (.A1(_01189_),
    .A2(_00953_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25412_ (.A1(_01414_),
    .A2(_01195_),
    .B(_01035_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25413_ (.A1(net1233),
    .A2(_01162_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25414_ (.A1(_01416_),
    .A2(_01303_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25415_ (.A1(_01415_),
    .A2(_01417_),
    .B(_01009_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25416_ (.A1(_00981_),
    .A2(net1096),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25417_ (.A1(_01081_),
    .A2(_01419_),
    .A3(_00997_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25418_ (.A1(_01040_),
    .A2(_00902_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25419_ (.A1(_01421_),
    .A2(_01024_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25420_ (.A1(_01320_),
    .A2(_01254_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25421_ (.A1(_01422_),
    .A2(_01423_),
    .A3(_00941_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25422_ (.A1(_01420_),
    .A2(_01424_),
    .A3(_01116_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25423_ (.A1(_01418_),
    .A2(_01425_),
    .B(_01017_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25424_ (.A1(_01413_),
    .A2(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25425_ (.I(_00943_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25426_ (.I(_01291_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25427_ (.A1(_01069_),
    .A2(_01428_),
    .B(_01429_),
    .C(_00983_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25428_ (.A1(_01185_),
    .A2(_01165_),
    .B(_00985_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25429_ (.A1(_01430_),
    .A2(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25430_ (.A1(_00989_),
    .A2(_01128_),
    .B(_01022_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25431_ (.A1(_00943_),
    .A2(_00976_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25432_ (.A1(_01433_),
    .A2(_01434_),
    .B(_01035_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25433_ (.A1(_01062_),
    .A2(_01045_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25434_ (.I(_01283_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25435_ (.A1(_01437_),
    .A2(_01231_),
    .A3(_01436_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25436_ (.A1(_01435_),
    .A2(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25437_ (.A1(_01439_),
    .A2(_01052_),
    .A3(_01432_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25438_ (.A1(_00943_),
    .A2(_00976_),
    .A3(net1095),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25439_ (.A1(_00990_),
    .A2(_01128_),
    .B(_01077_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25440_ (.A1(_01441_),
    .A2(_01442_),
    .B(_01035_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25441_ (.A1(_00949_),
    .A2(_00954_),
    .A3(_01371_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25442_ (.A1(_01443_),
    .A2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25443_ (.A1(net537),
    .A2(_01128_),
    .B(_01022_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25444_ (.A1(_01446_),
    .A2(_01105_),
    .B(_01043_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25445_ (.A1(_01062_),
    .A2(net498),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25446_ (.A1(_01421_),
    .A2(_01072_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25447_ (.A1(_01448_),
    .A2(_01449_),
    .A3(_01066_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25448_ (.A1(_01450_),
    .A2(_01447_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25449_ (.A1(_01445_),
    .A2(_01451_),
    .A3(_01181_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25450_ (.A1(_01440_),
    .A2(_01017_),
    .A3(_01452_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25451_ (.A1(_01453_),
    .A2(_01427_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25452_ (.A1(_01133_),
    .A2(_01165_),
    .B(_01126_),
    .C(_01066_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25453_ (.A1(_00952_),
    .A2(_15917_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25454_ (.A1(_01449_),
    .A2(_00997_),
    .A3(_01455_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25455_ (.A1(_01454_),
    .A2(_01116_),
    .A3(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25456_ (.A1(_01201_),
    .A2(_00983_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25457_ (.I(_01046_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25458_ (.A1(_01369_),
    .A2(_01459_),
    .B(_00983_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25459_ (.A1(_01458_),
    .A2(_01460_),
    .B(_00969_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25460_ (.A1(_01457_),
    .A2(_01461_),
    .A3(_01052_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25461_ (.A1(_00903_),
    .A2(net21),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25462_ (.A1(_01308_),
    .A2(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25463_ (.A1(_01464_),
    .A2(_00997_),
    .B(_00985_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25464_ (.A1(_01268_),
    .A2(_01135_),
    .B(_01019_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25465_ (.A1(_01466_),
    .A2(_01241_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25466_ (.A1(_01465_),
    .A2(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25467_ (.A1(_01186_),
    .A2(_00953_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25468_ (.A1(_01469_),
    .A2(_01061_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25469_ (.A1(_01133_),
    .A2(_00976_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25470_ (.A1(_01303_),
    .A2(_01082_),
    .A3(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25471_ (.A1(_01470_),
    .A2(_01472_),
    .A3(_01084_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25472_ (.A1(_01468_),
    .A2(_01473_),
    .A3(_01181_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25473_ (.A1(_01462_),
    .A2(_01474_),
    .A3(_01017_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25474_ (.A1(_01347_),
    .A2(net1267),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25475_ (.A1(_00990_),
    .A2(_01088_),
    .B(_01077_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25476_ (.A1(_01476_),
    .A2(_01477_),
    .B(_01035_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25477_ (.A1(_01024_),
    .A2(_01048_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25478_ (.A1(_01479_),
    .A2(_01125_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25479_ (.A1(_01176_),
    .A2(_01290_),
    .B(_01022_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25480_ (.A1(_01480_),
    .A2(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25481_ (.A1(_01478_),
    .A2(_01482_),
    .B(_01180_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25482_ (.A1(_01393_),
    .A2(_01133_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25483_ (.A1(_01484_),
    .A2(_01162_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25484_ (.A1(_01057_),
    .A2(_00992_),
    .A3(net1229),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25485_ (.A1(_01485_),
    .A2(_01486_),
    .B(_00985_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25486_ (.A1(_01437_),
    .A2(_01243_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25487_ (.A1(_01488_),
    .A2(_01241_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25488_ (.A1(_01487_),
    .A2(_01489_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25489_ (.A1(_01483_),
    .A2(_01490_),
    .B(_01017_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25490_ (.A1(_00911_),
    .A2(_01212_),
    .B(_01032_),
    .C(_01371_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25491_ (.A1(_01421_),
    .A2(_01076_),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25492_ (.A1(_01493_),
    .A2(_01049_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25493_ (.I(_01257_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25494_ (.A1(_01494_),
    .A2(_01495_),
    .B(_00983_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25495_ (.A1(_01492_),
    .A2(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25496_ (.A1(_01497_),
    .A2(_00969_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25497_ (.A1(_01264_),
    .A2(net1266),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25498_ (.A1(_15916_),
    .A2(_15925_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25499_ (.A1(_00976_),
    .A2(_01500_),
    .B(_01022_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25500_ (.A1(_01499_),
    .A2(_01501_),
    .B(_00985_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25501_ (.A1(_01232_),
    .A2(_01028_),
    .B(_00992_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25502_ (.A1(_01384_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25503_ (.A1(_01502_),
    .A2(_01504_),
    .B(_01009_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25504_ (.A1(_01498_),
    .A2(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25505_ (.A1(_01506_),
    .A2(_01491_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25506_ (.A1(_01507_),
    .A2(_01475_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25507_ (.A1(_01110_),
    .A2(_00904_),
    .A3(net1229),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25508_ (.A1(_01340_),
    .A2(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25509_ (.A1(_00903_),
    .A2(net34),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25510_ (.A1(_01348_),
    .A2(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25511_ (.A1(_01511_),
    .A2(_01241_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25512_ (.A1(_01509_),
    .A2(_01116_),
    .A3(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25513_ (.A1(_00904_),
    .A2(_01330_),
    .B(_01437_),
    .C(_01082_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25514_ (.A1(_01098_),
    .A2(_01110_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25515_ (.A1(_01515_),
    .A2(_01479_),
    .A3(_01241_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25516_ (.A1(_01516_),
    .A2(_00969_),
    .A3(_01514_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25517_ (.A1(_01513_),
    .A2(_01517_),
    .A3(_01052_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25518_ (.A1(_01140_),
    .A2(_01024_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25519_ (.A1(_01325_),
    .A2(_01257_),
    .A3(_01519_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25520_ (.A1(_01135_),
    .A2(_01162_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25521_ (.A1(_01521_),
    .A2(_01369_),
    .B(_01043_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25522_ (.A1(_01520_),
    .A2(_01522_),
    .B(_01009_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25523_ (.A1(_01265_),
    .A2(_01493_),
    .A3(_01082_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25524_ (.A1(_01289_),
    .A2(_01183_),
    .A3(_00941_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25525_ (.A1(_01524_),
    .A2(_01525_),
    .A3(_00969_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25526_ (.A1(_01523_),
    .A2(_01526_),
    .B(_01018_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25527_ (.A1(_01518_),
    .A2(_01527_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25528_ (.A1(_00904_),
    .A2(net1231),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25529_ (.A1(_01499_),
    .A2(_01529_),
    .A3(_01241_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25530_ (.A1(_01080_),
    .A2(_01128_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25531_ (.A1(_01082_),
    .A2(_01531_),
    .A3(_01029_),
    .A4(_01020_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25532_ (.A1(_01530_),
    .A2(_01532_),
    .A3(_00969_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25533_ (.A1(_01256_),
    .A2(_01087_),
    .B(_00976_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25534_ (.A1(_01045_),
    .A2(_01096_),
    .A3(_01128_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25535_ (.A1(_01534_),
    .A2(_00997_),
    .A3(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25536_ (.A1(_01510_),
    .A2(_15915_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25537_ (.A1(_01463_),
    .A2(_00940_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25538_ (.A1(_01537_),
    .A2(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25539_ (.A1(_01539_),
    .A2(_01296_),
    .B(_01043_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25540_ (.A1(_01536_),
    .A2(_01540_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25541_ (.A1(_01533_),
    .A2(_01541_),
    .A3(_01181_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25542_ (.A1(_01378_),
    .A2(_00947_),
    .B(_01022_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25543_ (.A1(_01543_),
    .A2(_01029_),
    .B(_01043_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25544_ (.I(_01538_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25545_ (.A1(_01121_),
    .A2(_01371_),
    .A3(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25546_ (.A1(_01544_),
    .A2(_01546_),
    .B(_01180_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25547_ (.A1(_01280_),
    .A2(_01088_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25548_ (.A1(_00947_),
    .A2(_15925_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25549_ (.A1(_01082_),
    .A2(_01233_),
    .A3(_01548_),
    .A4(_01549_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25550_ (.A1(_01140_),
    .A2(net1229),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25551_ (.A1(_01094_),
    .A2(_01096_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25552_ (.A1(_01551_),
    .A2(_01552_),
    .A3(_01066_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25553_ (.A1(_01550_),
    .A2(_01553_),
    .A3(_01084_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25554_ (.A1(_01547_),
    .A2(_01554_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25555_ (.A1(_01542_),
    .A2(_01018_),
    .A3(_01555_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25556_ (.A1(_01528_),
    .A2(_01556_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25557_ (.I(\sa30_sr[7] ),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25558_ (.A1(_01557_),
    .A2(\sa30_sr[0] ),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25559_ (.A1(_10391_),
    .A2(_10635_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25560_ (.A1(_01558_),
    .A2(_01559_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25561_ (.A1(net607),
    .A2(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25562_ (.A1(_10416_),
    .A2(_10415_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25563_ (.A1(_01562_),
    .A2(_13583_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25564_ (.A1(_10420_),
    .A2(_10419_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25565_ (.A1(_01564_),
    .A2(_13587_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25566_ (.A1(_01565_),
    .A2(_01563_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25567_ (.I(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25568_ (.A1(_01567_),
    .A2(_01561_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25569_ (.A1(_10343_),
    .A2(_01560_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25570_ (.A1(_01569_),
    .A2(_01566_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25571_ (.A1(_01570_),
    .A2(_01568_),
    .B(_10586_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25572_ (.I(\text_in_r[105] ),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25573_ (.A1(_01572_),
    .A2(_10482_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _25574_ (.A1(_01573_),
    .A2(_01571_),
    .B(\u0.w[0][9] ),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25575_ (.A1(_01570_),
    .A2(_01568_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25576_ (.A1(_10479_),
    .A2(_01575_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25577_ (.I(\u0.w[0][9] ),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25578_ (.I(_01573_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25579_ (.A1(_01576_),
    .A2(_01577_),
    .A3(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25580_ (.A1(_01574_),
    .A2(_01579_),
    .ZN(_15935_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25581_ (.A1(net1067),
    .A2(net576),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25582_ (.A1(_01580_),
    .A2(_10634_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25583_ (.A1(_10339_),
    .A2(_10357_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25584_ (.A1(net1067),
    .A2(net576),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25585_ (.A1(_01582_),
    .A2(_01583_),
    .B(_13580_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25586_ (.A1(_01581_),
    .A2(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25587_ (.A1(_10391_),
    .A2(_01557_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25588_ (.A1(net580),
    .A2(_10635_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25589_ (.A1(_01587_),
    .A2(_01586_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25590_ (.A1(_01585_),
    .A2(net1085),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25591_ (.A1(_01581_),
    .A2(_01584_),
    .A3(_01560_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25592_ (.A1(_01589_),
    .A2(_01590_),
    .B(_10483_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25593_ (.I(\text_in_r[104] ),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25594_ (.A1(_01592_),
    .A2(_10410_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25595_ (.A1(net885),
    .A2(_01593_),
    .B(\u0.w[0][8] ),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25596_ (.A1(_01589_),
    .A2(_01590_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25597_ (.A1(_01595_),
    .A2(_10403_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25598_ (.I(\u0.w[0][8] ),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25599_ (.I(_01593_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25600_ (.A1(net1119),
    .A2(_01597_),
    .A3(_01598_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25601_ (.A1(_01599_),
    .A2(_01594_),
    .ZN(_15940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25602_ (.A1(_10427_),
    .A2(_10450_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25603_ (.A1(_10424_),
    .A2(_10426_),
    .A3(\sa00_sr[2] ),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25604_ (.A1(_01600_),
    .A2(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25605_ (.A1(_01602_),
    .A2(net691),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25606_ (.A1(_01600_),
    .A2(_01601_),
    .A3(net689),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25607_ (.A1(_01603_),
    .A2(_01604_),
    .B(_10482_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25608_ (.I(\text_in_r[106] ),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25609_ (.A1(_01606_),
    .A2(net594),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25610_ (.I(\u0.w[0][10] ),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25611_ (.A1(_01605_),
    .A2(_01607_),
    .B(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25612_ (.A1(_01603_),
    .A2(_01604_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25613_ (.A1(_01610_),
    .A2(_14333_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25614_ (.I(_01607_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25615_ (.A1(_01611_),
    .A2(\u0.w[0][10] ),
    .A3(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25616_ (.A1(_01613_),
    .A2(_01609_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _25617_ (.I(_01614_),
    .Z(_15956_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _25618_ (.A1(_01573_),
    .A2(_01571_),
    .B(_01577_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25619_ (.A1(_01576_),
    .A2(\u0.w[0][9] ),
    .A3(_01578_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25620_ (.A1(_01615_),
    .A2(_01616_),
    .ZN(_15930_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25621_ (.A1(_01605_),
    .A2(_01607_),
    .B(\u0.w[0][10] ),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25622_ (.A1(_01611_),
    .A2(_01608_),
    .A3(_01612_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25623_ (.A1(_01617_),
    .A2(_01618_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _25624_ (.I(_01619_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _25625_ (.I(_01620_),
    .Z(_15949_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25626_ (.A1(_01593_),
    .A2(_01591_),
    .B(_01597_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25627_ (.A1(_01596_),
    .A2(\u0.w[0][8] ),
    .A3(_01598_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25628_ (.A1(_01622_),
    .A2(_01621_),
    .ZN(_15929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25629_ (.A1(net858),
    .A2(net495),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25630_ (.A1(_10466_),
    .A2(_13689_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25631_ (.A1(\sa10_sr[3] ),
    .A2(\sa00_sr[3] ),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25632_ (.A1(_01624_),
    .A2(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25633_ (.I(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25634_ (.A1(_10423_),
    .A2(_01557_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25635_ (.A1(\sa30_sr[2] ),
    .A2(_10635_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25636_ (.A1(_01628_),
    .A2(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25637_ (.A1(_01627_),
    .A2(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25638_ (.I(_01630_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25639_ (.A1(_01632_),
    .A2(_01626_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25640_ (.A1(_01631_),
    .A2(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25641_ (.A1(\sa30_sr[3] ),
    .A2(_13679_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25642_ (.A1(_01634_),
    .A2(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25643_ (.A1(_10459_),
    .A2(_13679_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25644_ (.A1(_01631_),
    .A2(_01633_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25645_ (.A1(_01637_),
    .A2(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25646_ (.A1(_01636_),
    .A2(_01639_),
    .A3(_14333_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25647_ (.A1(_11203_),
    .A2(\text_in_r[107] ),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25648_ (.A1(_01640_),
    .A2(_01641_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25649_ (.A1(\u0.w[0][11] ),
    .A2(_01642_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25650_ (.I(\u0.w[0][11] ),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25651_ (.A1(_01640_),
    .A2(_01644_),
    .A3(_01641_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25652_ (.A1(_01645_),
    .A2(_01643_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25653_ (.A1(_01623_),
    .A2(net1213),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25654_ (.A1(_13648_),
    .A2(_13655_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25655_ (.I(_10542_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25656_ (.A1(\sa30_sr[3] ),
    .A2(net68),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25657_ (.A1(_01649_),
    .A2(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _25658_ (.A1(\sa30_sr[3] ),
    .A2(_10635_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25659_ (.A1(_01652_),
    .A2(_10542_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25660_ (.A1(_01651_),
    .A2(_01653_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25661_ (.A1(_01648_),
    .A2(_01654_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25662_ (.A1(_01648_),
    .A2(_01654_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25663_ (.A1(_01655_),
    .A2(_01656_),
    .A3(_10523_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25664_ (.A1(_10526_),
    .A2(\text_in_r[108] ),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25665_ (.A1(_01657_),
    .A2(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25666_ (.A1(_01659_),
    .A2(\u0.w[0][12] ),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25667_ (.I(\u0.w[0][12] ),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25668_ (.A1(_01657_),
    .A2(_01661_),
    .A3(_01658_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25669_ (.A1(_01660_),
    .A2(_01662_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25670_ (.I(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25671_ (.A1(_01647_),
    .A2(_01664_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25672_ (.I(_01614_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25673_ (.A1(_01666_),
    .A2(_15936_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25674_ (.A1(_01642_),
    .A2(_01644_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25675_ (.A1(_01640_),
    .A2(\u0.w[0][11] ),
    .A3(_01641_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25676_ (.A1(_01668_),
    .A2(_01669_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25677_ (.I(_01670_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25678_ (.A1(_01667_),
    .A2(_01671_),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25679_ (.I(_15938_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25680_ (.A1(_15949_),
    .A2(_01673_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25681_ (.A1(_01672_),
    .A2(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25682_ (.A1(\sa30_sr[5] ),
    .A2(_13651_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25683_ (.A1(_01676_),
    .A2(_10581_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25684_ (.A1(_01676_),
    .A2(_10581_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25685_ (.A1(_01677_),
    .A2(_01678_),
    .A3(_10403_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25686_ (.A1(_12115_),
    .A2(\text_in_r[109] ),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25687_ (.A1(_01679_),
    .A2(_01680_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25688_ (.A1(_01681_),
    .A2(\u0.w[0][13] ),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25689_ (.A1(_01681_),
    .A2(\u0.w[0][13] ),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25690_ (.A1(_01682_),
    .A2(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25691_ (.I(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25692_ (.I(_01685_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25693_ (.A1(_01665_),
    .A2(_01675_),
    .B(_01686_),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25694_ (.I(_01646_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25695_ (.A1(_01688_),
    .A2(_01667_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25696_ (.I(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25697_ (.A1(net495),
    .A2(net886),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25698_ (.A1(_01690_),
    .A2(_01691_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25699_ (.A1(_01659_),
    .A2(_01661_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25700_ (.A1(_01657_),
    .A2(\u0.w[0][12] ),
    .A3(_01658_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25701_ (.A1(_01693_),
    .A2(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25702_ (.I(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25703_ (.I(_01696_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25704_ (.A1(net621),
    .A2(net886),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25705_ (.A1(_01666_),
    .A2(_15947_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25706_ (.A1(_01698_),
    .A2(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25707_ (.I(_01671_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25708_ (.A1(_01700_),
    .A2(_01701_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25709_ (.A1(_01692_),
    .A2(_01697_),
    .A3(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25710_ (.A1(\sa10_sr[6] ),
    .A2(\sa30_sr[6] ),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25711_ (.A1(_13742_),
    .A2(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25712_ (.A1(_01705_),
    .A2(_10545_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25713_ (.A1(_01705_),
    .A2(_10545_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25714_ (.A1(_10587_),
    .A2(\text_in_r[110] ),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _25715_ (.A1(_01706_),
    .A2(_10639_),
    .A3(_01707_),
    .B(_01708_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25716_ (.A1(_01709_),
    .A2(\u0.w[0][14] ),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25717_ (.A1(_01709_),
    .A2(\u0.w[0][14] ),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25718_ (.A1(_01710_),
    .A2(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25719_ (.I(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25720_ (.A1(_01687_),
    .A2(_01703_),
    .B(_01713_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25721_ (.A1(_15930_),
    .A2(_01614_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25722_ (.I(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25723_ (.I(_01646_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25724_ (.A1(_01716_),
    .A2(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25725_ (.A1(net886),
    .A2(_15933_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25726_ (.A1(_01719_),
    .A2(_01670_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25727_ (.A1(_01720_),
    .A2(_01695_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25728_ (.A1(_15945_),
    .A2(_01619_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25729_ (.A1(_01623_),
    .A2(_01722_),
    .A3(_01671_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25730_ (.A1(_01718_),
    .A2(_01721_),
    .A3(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25731_ (.A1(net27),
    .A2(_15949_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25732_ (.I(_01725_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25733_ (.A1(_01690_),
    .A2(net1137),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25734_ (.I(_01671_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25735_ (.I(_15947_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25736_ (.A1(net886),
    .A2(_01729_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25737_ (.A1(_01623_),
    .A2(_01728_),
    .A3(net1215),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25738_ (.I(_01696_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25739_ (.A1(_01727_),
    .A2(_01731_),
    .A3(_01732_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25740_ (.I(_01685_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25741_ (.A1(_01724_),
    .A2(_01733_),
    .A3(_01734_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _25742_ (.A1(net68),
    .A2(_10389_),
    .A3(_10582_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25743_ (.A1(_10639_),
    .A2(\text_in_r[111] ),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25744_ (.A1(_01736_),
    .A2(_12965_),
    .B(_01737_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _25745_ (.A1(\u0.w[0][15] ),
    .A2(_01738_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25746_ (.I(_01739_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25747_ (.I(_01740_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25748_ (.A1(_01714_),
    .A2(_01735_),
    .B(_01741_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25749_ (.I(_15932_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25750_ (.A1(net886),
    .A2(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25751_ (.I(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25752_ (.A1(_01745_),
    .A2(net1214),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25753_ (.I(_01746_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _25754_ (.I(_01670_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25755_ (.I(_01748_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25756_ (.A1(_01666_),
    .A2(net1139),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25757_ (.A1(_01749_),
    .A2(_01750_),
    .B(_01663_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25758_ (.A1(_01718_),
    .A2(_01747_),
    .A3(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25759_ (.I(_15941_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25760_ (.A1(_15956_),
    .A2(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25761_ (.I(_01754_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25762_ (.I(_15931_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25763_ (.A1(net886),
    .A2(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25764_ (.I(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25765_ (.I(_01688_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25766_ (.A1(_01755_),
    .A2(_01758_),
    .B(_01759_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25767_ (.A1(_01748_),
    .A2(_01744_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _25768_ (.I(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25769_ (.A1(_15956_),
    .A2(_15931_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25770_ (.A1(_01762_),
    .A2(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25771_ (.I(_01695_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25772_ (.A1(_01764_),
    .A2(_01760_),
    .B(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25773_ (.A1(_01752_),
    .A2(_01766_),
    .B(_01734_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25774_ (.A1(net863),
    .A2(net886),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25775_ (.A1(_01768_),
    .A2(_01688_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25776_ (.A1(net1120),
    .A2(net495),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25777_ (.A1(_01769_),
    .A2(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25778_ (.A1(net588),
    .A2(net494),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25779_ (.I(_01748_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25780_ (.A1(net863),
    .A2(net858),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25781_ (.A1(_01772_),
    .A2(_01773_),
    .A3(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25782_ (.A1(_01771_),
    .A2(_01775_),
    .A3(_01732_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _25783_ (.I(_01684_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25784_ (.I(_01777_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25785_ (.A1(_01744_),
    .A2(_01717_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25786_ (.A1(_01666_),
    .A2(_15945_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25787_ (.A1(_01779_),
    .A2(_01780_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25788_ (.I(_01663_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25789_ (.A1(_15949_),
    .A2(_15941_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25790_ (.I(_01748_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25791_ (.A1(_01763_),
    .A2(_01783_),
    .A3(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25792_ (.A1(_01781_),
    .A2(_01782_),
    .A3(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25793_ (.A1(_01776_),
    .A2(_01778_),
    .A3(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25794_ (.A1(_01787_),
    .A2(_01713_),
    .A3(_01767_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25795_ (.A1(_01742_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25796_ (.A1(net621),
    .A2(net857),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25797_ (.A1(_01790_),
    .A2(_01688_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25798_ (.I(net1213),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25799_ (.A1(_01792_),
    .A2(_15954_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25800_ (.A1(_01791_),
    .A2(_01793_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25801_ (.I(_01777_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25802_ (.A1(_01794_),
    .A2(_01697_),
    .B(_01795_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25803_ (.I(_15936_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25804_ (.A1(_01797_),
    .A2(_15949_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25805_ (.A1(net858),
    .A2(_15938_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25806_ (.A1(_01798_),
    .A2(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25807_ (.I(_01646_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25808_ (.A1(_01800_),
    .A2(_01801_),
    .B(_01696_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25809_ (.A1(_01774_),
    .A2(_01757_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25810_ (.A1(_01803_),
    .A2(_01773_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25811_ (.A1(_15956_),
    .A2(_15933_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25812_ (.I(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25813_ (.I(_01717_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25814_ (.A1(_01806_),
    .A2(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25815_ (.A1(_01802_),
    .A2(_01804_),
    .A3(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25816_ (.A1(_01796_),
    .A2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25817_ (.A1(_01755_),
    .A2(_01801_),
    .B(_01663_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25818_ (.I(_01719_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25819_ (.A1(_01812_),
    .A2(_01748_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25820_ (.I(_01798_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25821_ (.A1(_01717_),
    .A2(_01814_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25822_ (.A1(_01811_),
    .A2(_01813_),
    .A3(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25823_ (.I(_15943_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25824_ (.A1(_01817_),
    .A2(_01666_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25825_ (.A1(_01818_),
    .A2(_01748_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25826_ (.A1(_15949_),
    .A2(_15936_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25827_ (.A1(_01819_),
    .A2(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25828_ (.A1(_01821_),
    .A2(_01721_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25829_ (.A1(_01816_),
    .A2(_01822_),
    .A3(_01795_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25830_ (.A1(_01810_),
    .A2(_01823_),
    .A3(_01713_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25831_ (.A1(_01666_),
    .A2(_01756_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25832_ (.A1(_01825_),
    .A2(_01792_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25833_ (.A1(_01674_),
    .A2(_01671_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25834_ (.A1(_01826_),
    .A2(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25835_ (.A1(_01720_),
    .A2(_01664_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25836_ (.A1(_01828_),
    .A2(_01829_),
    .B(_01686_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25837_ (.A1(_01666_),
    .A2(_15941_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25838_ (.A1(net586),
    .A2(_15956_),
    .B(_01831_),
    .C(_01784_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25839_ (.A1(net479),
    .A2(_15949_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25840_ (.A1(_01833_),
    .A2(_01792_),
    .A3(net1113),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25841_ (.A1(_01832_),
    .A2(_01782_),
    .A3(_01834_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25842_ (.A1(_01830_),
    .A2(_01835_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25843_ (.A1(net886),
    .A2(_15943_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25844_ (.I(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25845_ (.A1(_01838_),
    .A2(_01717_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25846_ (.A1(_01839_),
    .A2(_01761_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25847_ (.I(_01799_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25848_ (.A1(_01841_),
    .A2(_01688_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25849_ (.A1(_01842_),
    .A2(_01695_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25850_ (.A1(_01840_),
    .A2(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25851_ (.I(_01663_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25852_ (.A1(_01723_),
    .A2(_01845_),
    .A3(_01842_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25853_ (.A1(_01844_),
    .A2(_01846_),
    .A3(_01686_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _25854_ (.I(_01712_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25855_ (.I(_01848_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25856_ (.A1(_01836_),
    .A2(_01847_),
    .A3(_01849_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25857_ (.A1(_01824_),
    .A2(_01850_),
    .A3(_01741_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25858_ (.A1(_01789_),
    .A2(_01851_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25859_ (.A1(_01792_),
    .A2(_15961_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25860_ (.A1(_01726_),
    .A2(_01749_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25861_ (.A1(_01843_),
    .A2(_01852_),
    .A3(_01853_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25862_ (.A1(_01730_),
    .A2(_01750_),
    .A3(_01749_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25863_ (.A1(_01802_),
    .A2(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25864_ (.A1(_01854_),
    .A2(_01856_),
    .A3(_01734_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25865_ (.A1(_01762_),
    .A2(_01623_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25866_ (.A1(_01674_),
    .A2(_01688_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25867_ (.I(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25868_ (.A1(_01860_),
    .A2(_01774_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25869_ (.A1(_01858_),
    .A2(_01861_),
    .A3(_01732_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25870_ (.A1(_01833_),
    .A2(_01770_),
    .A3(_01717_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25871_ (.A1(_15956_),
    .A2(_01797_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25872_ (.I(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25873_ (.I(_01695_),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25874_ (.A1(_01865_),
    .A2(_01728_),
    .B(_01866_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25875_ (.A1(_01863_),
    .A2(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25876_ (.A1(_01862_),
    .A2(_01868_),
    .A3(_01778_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25877_ (.A1(_01857_),
    .A2(_01713_),
    .A3(_01869_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25878_ (.A1(_01780_),
    .A2(_01748_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25879_ (.A1(_01871_),
    .A2(_01698_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25880_ (.A1(_15949_),
    .A2(_15938_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25881_ (.I(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25882_ (.A1(_01874_),
    .A2(_01759_),
    .B(_01866_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25883_ (.A1(_01872_),
    .A2(_01875_),
    .B(_01686_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25884_ (.A1(_01666_),
    .A2(_01729_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25885_ (.A1(_01877_),
    .A2(_01748_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25886_ (.A1(_01878_),
    .A2(_01726_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25887_ (.I(_15945_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25888_ (.A1(_15949_),
    .A2(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25889_ (.A1(_01881_),
    .A2(_01807_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25890_ (.A1(_01879_),
    .A2(_01732_),
    .A3(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25891_ (.A1(_01876_),
    .A2(_01883_),
    .B(_01712_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25892_ (.A1(net63),
    .A2(net586),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25893_ (.A1(_01885_),
    .A2(_01691_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25894_ (.A1(_01886_),
    .A2(_01701_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25895_ (.A1(_01791_),
    .A2(_01691_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25896_ (.A1(_01887_),
    .A2(_01888_),
    .A3(_01782_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25897_ (.A1(_01841_),
    .A2(_01745_),
    .B(_01728_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25898_ (.A1(_01803_),
    .A2(_01807_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25899_ (.A1(_01890_),
    .A2(_01891_),
    .A3(_01765_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25900_ (.I(_01685_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25901_ (.A1(_01889_),
    .A2(_01892_),
    .A3(_01893_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25902_ (.A1(_01884_),
    .A2(_01894_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25903_ (.A1(_01870_),
    .A2(_01741_),
    .A3(_01895_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25904_ (.A1(_01716_),
    .A2(_01827_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25905_ (.A1(net63),
    .A2(_15956_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25906_ (.A1(_01769_),
    .A2(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25907_ (.A1(_01897_),
    .A2(_01899_),
    .A3(_01686_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25908_ (.A1(_01691_),
    .A2(_01717_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25909_ (.A1(_01901_),
    .A2(_01763_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25910_ (.A1(_01672_),
    .A2(net1114),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25911_ (.A1(_01902_),
    .A2(_01903_),
    .A3(_01795_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25912_ (.A1(_01900_),
    .A2(_01904_),
    .A3(_01697_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25913_ (.A1(_01685_),
    .A2(_01748_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25914_ (.A1(_01722_),
    .A2(_01646_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25915_ (.I(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25916_ (.A1(_01908_),
    .A2(_01831_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25917_ (.A1(_15957_),
    .A2(_01906_),
    .B(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _25918_ (.I(_01663_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25919_ (.A1(_01910_),
    .A2(_01911_),
    .B(_01848_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25920_ (.A1(_01905_),
    .A2(_01912_),
    .B(_01741_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25921_ (.A1(_01701_),
    .A2(_01758_),
    .B(_01720_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25922_ (.I(_01774_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25923_ (.A1(_01915_),
    .A2(_01759_),
    .B(_01664_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25924_ (.A1(_01688_),
    .A2(_01790_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25925_ (.I(_01917_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25926_ (.A1(_01914_),
    .A2(_01916_),
    .A3(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25927_ (.A1(_01769_),
    .A2(_01763_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25928_ (.A1(_01897_),
    .A2(_01920_),
    .A3(_01782_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25929_ (.A1(_01919_),
    .A2(_01921_),
    .A3(_01778_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25930_ (.I(_01647_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25931_ (.A1(_01923_),
    .A2(net1114),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25932_ (.A1(_01924_),
    .A2(_01782_),
    .A3(_01761_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25933_ (.I(_15933_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25934_ (.A1(_01666_),
    .A2(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25935_ (.A1(_01927_),
    .A2(_01688_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25936_ (.I(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25937_ (.A1(_01929_),
    .A2(net1215),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25938_ (.A1(_01872_),
    .A2(_01930_),
    .A3(_01765_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25939_ (.A1(_01925_),
    .A2(_01931_),
    .A3(_01893_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25940_ (.A1(_01922_),
    .A2(_01932_),
    .A3(_01849_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25941_ (.A1(_01913_),
    .A2(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25942_ (.A1(_01934_),
    .A2(_01896_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25943_ (.A1(_01689_),
    .A2(_01664_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25944_ (.A1(_01871_),
    .A2(net1215),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25945_ (.A1(_01935_),
    .A2(_01936_),
    .B(_01848_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25946_ (.A1(_01898_),
    .A2(_01807_),
    .A3(_01744_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25947_ (.A1(_01768_),
    .A2(_01805_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25948_ (.A1(_01939_),
    .A2(_01701_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25949_ (.A1(_01938_),
    .A2(_01940_),
    .A3(_01732_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25950_ (.A1(_01937_),
    .A2(_01941_),
    .B(_01893_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25951_ (.A1(_01818_),
    .A2(net1212),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25952_ (.A1(_01943_),
    .A2(_01691_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25953_ (.A1(_01762_),
    .A2(net1113),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _25954_ (.I(_01695_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25955_ (.A1(_01945_),
    .A2(_01944_),
    .B(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25956_ (.A1(_01715_),
    .A2(_01749_),
    .A3(_01837_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25957_ (.A1(_01768_),
    .A2(_01699_),
    .A3(_01792_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25958_ (.A1(_01949_),
    .A2(_01946_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25959_ (.A1(_01948_),
    .A2(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25960_ (.A1(_01947_),
    .A2(_01951_),
    .B(_01849_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25961_ (.A1(_01942_),
    .A2(_01952_),
    .B(_01741_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25962_ (.A1(_01798_),
    .A2(_01748_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25963_ (.A1(_01954_),
    .A2(_01799_),
    .B(_01695_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25964_ (.A1(_01955_),
    .A2(_01834_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25965_ (.A1(_01956_),
    .A2(_01712_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25966_ (.A1(_01672_),
    .A2(_01833_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25967_ (.A1(_01699_),
    .A2(_01873_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25968_ (.A1(_01959_),
    .A2(_01759_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25969_ (.A1(_01958_),
    .A2(_01960_),
    .B(_01845_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25970_ (.A1(_01957_),
    .A2(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25971_ (.A1(_01666_),
    .A2(_01673_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25972_ (.A1(_01691_),
    .A2(_01728_),
    .A3(_01963_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25973_ (.A1(_01699_),
    .A2(_01749_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25974_ (.A1(_01964_),
    .A2(_01732_),
    .A3(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25975_ (.A1(_01833_),
    .A2(_01807_),
    .B(_01845_),
    .C(_01799_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25976_ (.A1(_01848_),
    .A2(_01839_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25977_ (.A1(_01966_),
    .A2(_01967_),
    .B(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25978_ (.A1(_01962_),
    .A2(_01969_),
    .B(_01734_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25979_ (.A1(_01953_),
    .A2(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25980_ (.A1(net27),
    .A2(_15956_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _25981_ (.A1(_01972_),
    .A2(_01784_),
    .A3(_01825_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25982_ (.A1(_15949_),
    .A2(_01753_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25983_ (.A1(_01645_),
    .A2(_01790_),
    .A3(_01974_),
    .A4(net1216),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25984_ (.A1(_01973_),
    .A2(_01975_),
    .B(_01911_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25985_ (.A1(_01833_),
    .A2(_01770_),
    .A3(_01749_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25986_ (.A1(_01749_),
    .A2(_15957_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25987_ (.A1(_01977_),
    .A2(_01782_),
    .A3(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25988_ (.A1(_01979_),
    .A2(_01734_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25989_ (.A1(_01715_),
    .A2(_01784_),
    .A3(_01691_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25990_ (.A1(_01981_),
    .A2(_01834_),
    .A3(_01765_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25991_ (.A1(_01820_),
    .A2(_01671_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25992_ (.A1(_01983_),
    .A2(_01750_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25993_ (.A1(_15954_),
    .A2(_01801_),
    .B(_01696_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25994_ (.A1(_01984_),
    .A2(_01985_),
    .B(_01685_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25995_ (.A1(_01982_),
    .A2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25996_ (.A1(_01976_),
    .A2(_01980_),
    .B(_01987_),
    .C(_01849_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25997_ (.A1(_01762_),
    .A2(_01963_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25998_ (.A1(_01758_),
    .A2(_01759_),
    .B(_01866_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25999_ (.A1(_01989_),
    .A2(_01990_),
    .B(_01686_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26000_ (.A1(_01926_),
    .A2(_01673_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26001_ (.A1(_01992_),
    .A2(net886),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26002_ (.A1(_01871_),
    .A2(net590),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26003_ (.A1(_01994_),
    .A2(_01909_),
    .A3(_01765_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26004_ (.A1(_01991_),
    .A2(_01995_),
    .B(_01848_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26005_ (.A1(_15952_),
    .A2(_01792_),
    .B(_01689_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26006_ (.A1(_01997_),
    .A2(_01946_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26007_ (.A1(_01759_),
    .A2(_15963_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26008_ (.A1(_01958_),
    .A2(_01765_),
    .A3(_01999_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26009_ (.A1(_01998_),
    .A2(_01893_),
    .A3(_02000_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26010_ (.A1(_01996_),
    .A2(_02001_),
    .B(_01739_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26011_ (.A1(_01988_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26012_ (.A1(_01971_),
    .A2(_02003_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26013_ (.A1(_01754_),
    .A2(_01744_),
    .A3(_01801_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26014_ (.A1(_01775_),
    .A2(_01946_),
    .A3(_02004_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26015_ (.A1(_01783_),
    .A2(_01667_),
    .A3(_01773_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26016_ (.A1(_01722_),
    .A2(_01750_),
    .A3(_01792_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26017_ (.A1(_02006_),
    .A2(_02007_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26018_ (.A1(_02008_),
    .A2(_01845_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26019_ (.A1(_02005_),
    .A2(_02009_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26020_ (.A1(_02010_),
    .A2(_01849_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26021_ (.A1(_01715_),
    .A2(_01807_),
    .A3(_01698_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26022_ (.A1(net1215),
    .A2(_01963_),
    .A3(_01728_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26023_ (.A1(_02012_),
    .A2(_01911_),
    .A3(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26024_ (.A1(_01774_),
    .A2(_01801_),
    .A3(_01974_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26025_ (.A1(_01757_),
    .A2(_01750_),
    .A3(_01749_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26026_ (.A1(_02015_),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26027_ (.A1(_02017_),
    .A2(_01697_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26028_ (.A1(_02014_),
    .A2(_02018_),
    .A3(_01713_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26029_ (.A1(_02011_),
    .A2(_02019_),
    .A3(_01778_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26030_ (.A1(_01715_),
    .A2(_01807_),
    .A3(_01691_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26031_ (.A1(_02021_),
    .A2(_01751_),
    .B(_01848_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26032_ (.A1(_01772_),
    .A2(_01759_),
    .A3(_01768_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26033_ (.A1(_01715_),
    .A2(_01728_),
    .A3(_01744_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26034_ (.A1(_02023_),
    .A2(_02024_),
    .A3(_01782_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26035_ (.A1(_02022_),
    .A2(_02025_),
    .B(_01778_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26036_ (.A1(_01943_),
    .A2(_01698_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26037_ (.A1(_01879_),
    .A2(_02027_),
    .A3(_01697_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26038_ (.I(_01672_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26039_ (.A1(_02023_),
    .A2(_01911_),
    .A3(_02029_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26040_ (.A1(_02028_),
    .A2(_02030_),
    .A3(_01849_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26041_ (.A1(_02026_),
    .A2(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26042_ (.A1(_02020_),
    .A2(_02032_),
    .A3(_01741_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26043_ (.A1(_01906_),
    .A2(_01750_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26044_ (.A1(_01813_),
    .A2(_01695_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26045_ (.A1(_02034_),
    .A2(_02035_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26046_ (.A1(_01831_),
    .A2(_01688_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _26047_ (.A1(_01972_),
    .A2(_01777_),
    .A3(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26048_ (.A1(_01746_),
    .A2(_01777_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26049_ (.A1(_02038_),
    .A2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26050_ (.A1(_02040_),
    .A2(_02036_),
    .B(_01848_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26051_ (.A1(_01878_),
    .A2(net589),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26052_ (.A1(_01623_),
    .A2(_01744_),
    .A3(_01717_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26053_ (.A1(_02042_),
    .A2(_02043_),
    .A3(_01685_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26054_ (.A1(_01838_),
    .A2(_01671_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26055_ (.A1(_01944_),
    .A2(_01777_),
    .A3(_02045_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26056_ (.A1(_02044_),
    .A2(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26057_ (.A1(_02047_),
    .A2(_01911_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26058_ (.A1(_02041_),
    .A2(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26059_ (.A1(_01863_),
    .A2(_01804_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26060_ (.A1(_02050_),
    .A2(_01845_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26061_ (.A1(_01700_),
    .A2(_01792_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26062_ (.A1(_01623_),
    .A2(_01837_),
    .B(_01717_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26063_ (.A1(_02052_),
    .A2(_02053_),
    .B(_01946_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26064_ (.A1(_02051_),
    .A2(_01795_),
    .A3(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26065_ (.A1(_01818_),
    .A2(_01993_),
    .A3(_01671_),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26066_ (.A1(_01909_),
    .A2(_02056_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26067_ (.A1(_02057_),
    .A2(_01664_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26068_ (.A1(_01949_),
    .A2(_01946_),
    .B(_01777_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26069_ (.A1(_02058_),
    .A2(_02059_),
    .B(_01712_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26070_ (.A1(_02055_),
    .A2(_02060_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26071_ (.A1(_02049_),
    .A2(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26072_ (.A1(_02062_),
    .A2(_01739_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26073_ (.A1(_02063_),
    .A2(_02033_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26074_ (.A1(_01918_),
    .A2(_01837_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26075_ (.A1(_01843_),
    .A2(_02064_),
    .B(_01686_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26076_ (.A1(_01730_),
    .A2(_01688_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26077_ (.A1(_02066_),
    .A2(_01750_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26078_ (.A1(_02067_),
    .A2(_01821_),
    .A3(_01911_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26079_ (.A1(_02065_),
    .A2(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26080_ (.A1(_01983_),
    .A2(_01715_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26081_ (.A1(_02070_),
    .A2(_01697_),
    .A3(_01960_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26082_ (.A1(_01898_),
    .A2(_01757_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26083_ (.A1(_02072_),
    .A2(_01701_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26084_ (.A1(_01802_),
    .A2(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26085_ (.A1(_02071_),
    .A2(_02074_),
    .A3(_01893_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26086_ (.A1(_02069_),
    .A2(_02075_),
    .A3(_01713_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26087_ (.A1(_01715_),
    .A2(_01768_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26088_ (.A1(_02077_),
    .A2(_01701_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26089_ (.A1(_02078_),
    .A2(_01902_),
    .A3(_01911_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26090_ (.I(_01819_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26091_ (.A1(_01696_),
    .A2(_01719_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26092_ (.A1(_02081_),
    .A2(_02080_),
    .B(_01686_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26093_ (.A1(_02079_),
    .A2(_02082_),
    .B(_01712_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26094_ (.A1(_01899_),
    .A2(_01977_),
    .A3(_01911_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26095_ (.A1(net1137),
    .A2(_01885_),
    .A3(_01807_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26096_ (.A1(net1137),
    .A2(_01728_),
    .A3(_01763_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26097_ (.A1(_02085_),
    .A2(_02086_),
    .A3(_01732_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26098_ (.A1(_02084_),
    .A2(_02087_),
    .A3(_01734_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26099_ (.A1(_02083_),
    .A2(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26100_ (.A1(_02076_),
    .A2(_02089_),
    .A3(_01741_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26101_ (.A1(_01790_),
    .A2(_01671_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26102_ (.A1(_01792_),
    .A2(_01880_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26103_ (.A1(_02091_),
    .A2(_01663_),
    .A3(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26104_ (.A1(_02093_),
    .A2(_01848_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26105_ (.A1(_01815_),
    .A2(_01696_),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26106_ (.A1(_01819_),
    .A2(_01725_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26107_ (.A1(_02095_),
    .A2(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26108_ (.A1(_02094_),
    .A2(_02097_),
    .B(_01893_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26109_ (.A1(_01723_),
    .A2(_01663_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26110_ (.A1(_01860_),
    .A2(net1113),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26111_ (.A1(_02099_),
    .A2(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26112_ (.A1(_01871_),
    .A2(_01929_),
    .A3(_01664_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26113_ (.A1(_02101_),
    .A2(_02102_),
    .A3(_01849_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26114_ (.A1(_02098_),
    .A2(_02103_),
    .B(_01740_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26115_ (.A1(_01769_),
    .A2(_01877_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26116_ (.A1(_01671_),
    .A2(_15956_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26117_ (.A1(_02106_),
    .A2(_01866_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26118_ (.A1(_02105_),
    .A2(_02107_),
    .B(_01712_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26119_ (.A1(_01758_),
    .A2(_01801_),
    .B(_01663_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26120_ (.A1(_01897_),
    .A2(_02109_),
    .A3(_01718_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26121_ (.A1(_02108_),
    .A2(_02110_),
    .B(_01778_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26122_ (.A1(_01772_),
    .A2(_01715_),
    .A3(_01792_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26123_ (.A1(_01819_),
    .A2(_01768_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26124_ (.A1(_02112_),
    .A2(_02113_),
    .A3(_01697_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26125_ (.A1(_01775_),
    .A2(_01721_),
    .A3(_01826_),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26126_ (.A1(_02114_),
    .A2(_02115_),
    .A3(_01713_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26127_ (.A1(_02111_),
    .A2(_02116_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26128_ (.A1(_02117_),
    .A2(_02104_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26129_ (.A1(_02118_),
    .A2(_02090_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26130_ (.A1(_01943_),
    .A2(_01820_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26131_ (.I(_01992_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26132_ (.A1(_01963_),
    .A2(_01773_),
    .A3(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26133_ (.A1(_02119_),
    .A2(_01866_),
    .A3(_02121_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26134_ (.A1(_01959_),
    .A2(_01773_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26135_ (.A1(_01718_),
    .A2(_01721_),
    .A3(_02123_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26136_ (.A1(_02122_),
    .A2(_02124_),
    .B(_01795_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26137_ (.A1(_02053_),
    .A2(_01779_),
    .B(_01664_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26138_ (.A1(_01859_),
    .A2(_01864_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26139_ (.A1(_02127_),
    .A2(_01946_),
    .B(_01795_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26140_ (.A1(_02126_),
    .A2(_02128_),
    .B(_01712_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26141_ (.A1(_02125_),
    .A2(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26142_ (.A1(net27),
    .A2(_01749_),
    .B(_01696_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26143_ (.A1(_02112_),
    .A2(_02131_),
    .B(_01685_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26144_ (.A1(_01923_),
    .A2(_01885_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26145_ (.A1(_01722_),
    .A2(_01831_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26146_ (.A1(_02134_),
    .A2(_01784_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26147_ (.A1(_02133_),
    .A2(_01946_),
    .A3(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26148_ (.A1(_02132_),
    .A2(_02136_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26149_ (.A1(_01761_),
    .A2(_01825_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26150_ (.A1(_01699_),
    .A2(_01801_),
    .B(_01696_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26151_ (.A1(_02138_),
    .A2(_02139_),
    .B(_01795_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26152_ (.A1(_01972_),
    .A2(_01928_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26153_ (.A1(_02141_),
    .A2(_01917_),
    .B(_01946_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26154_ (.A1(_02140_),
    .A2(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26155_ (.A1(_02143_),
    .A2(_01713_),
    .A3(_02137_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26156_ (.A1(_02130_),
    .A2(_02144_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26157_ (.A1(_01741_),
    .A2(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26158_ (.A1(_01901_),
    .A2(_01963_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26159_ (.A1(_02099_),
    .A2(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26160_ (.A1(_01908_),
    .A2(_01877_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26161_ (.A1(_01755_),
    .A2(_01784_),
    .B(_01664_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26162_ (.A1(_02149_),
    .A2(_02150_),
    .B(_01795_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26163_ (.A1(_02148_),
    .A2(_02151_),
    .B(_01712_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26164_ (.A1(_01701_),
    .A2(net864),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26165_ (.A1(_01771_),
    .A2(_01911_),
    .A3(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26166_ (.A1(_01943_),
    .A2(_01726_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26167_ (.A1(_01762_),
    .A2(_01667_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26168_ (.A1(_02155_),
    .A2(_02156_),
    .A3(_01732_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26169_ (.A1(_02154_),
    .A2(_02157_),
    .A3(_01778_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26170_ (.A1(_02158_),
    .A2(_02152_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26171_ (.I(_01878_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26172_ (.A1(_01843_),
    .A2(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26173_ (.A1(_01690_),
    .A2(_01722_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26174_ (.A1(_01728_),
    .A2(net589),
    .B(_01866_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26175_ (.A1(_02162_),
    .A2(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26176_ (.A1(_02161_),
    .A2(_01795_),
    .A3(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26177_ (.A1(_01773_),
    .A2(_01753_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26178_ (.A1(_01907_),
    .A2(_02166_),
    .A3(_01663_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26179_ (.A1(_02167_),
    .A2(_01685_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26180_ (.I(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26181_ (.A1(_01762_),
    .A2(_01831_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26182_ (.A1(_01698_),
    .A2(_01877_),
    .A3(_01801_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26183_ (.A1(_02170_),
    .A2(_01765_),
    .A3(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26184_ (.A1(_02169_),
    .A2(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26185_ (.A1(_02165_),
    .A2(_02173_),
    .A3(_01713_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26186_ (.A1(_02174_),
    .A2(_01739_),
    .A3(_02159_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26187_ (.A1(_02175_),
    .A2(_02146_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26188_ (.A1(_01770_),
    .A2(_01749_),
    .A3(_01774_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26189_ (.A1(_01726_),
    .A2(_01801_),
    .A3(_01864_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26190_ (.A1(_02176_),
    .A2(_02177_),
    .A3(_01664_),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26191_ (.A1(_02066_),
    .A2(_01774_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26192_ (.A1(_02176_),
    .A2(_02179_),
    .B(_01845_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26193_ (.A1(_02178_),
    .A2(_02180_),
    .B(_01778_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _26194_ (.A1(_01698_),
    .A2(_01773_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26195_ (.A1(_02053_),
    .A2(_01946_),
    .A3(_02182_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26196_ (.A1(_01692_),
    .A2(_01697_),
    .A3(_01852_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26197_ (.A1(_02183_),
    .A2(_01734_),
    .A3(_02184_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26198_ (.A1(_02181_),
    .A2(_02185_),
    .A3(_01849_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26199_ (.I(_15951_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26200_ (.A1(_02187_),
    .A2(_01784_),
    .B(_01866_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26201_ (.A1(_02188_),
    .A2(_02155_),
    .B(_01686_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26202_ (.A1(_01878_),
    .A2(_01698_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26203_ (.A1(_01916_),
    .A2(_02190_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26204_ (.A1(_02189_),
    .A2(_02191_),
    .B(_01848_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26205_ (.A1(_02096_),
    .A2(_02037_),
    .B(_01845_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26206_ (.A1(_02193_),
    .A2(_01955_),
    .B(_01893_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26207_ (.A1(_02194_),
    .A2(_02192_),
    .B(_01741_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26208_ (.A1(_02186_),
    .A2(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26209_ (.A1(_01772_),
    .A2(_01715_),
    .A3(_01784_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26210_ (.A1(_15950_),
    .A2(_15959_),
    .B(_01759_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26211_ (.A1(_02197_),
    .A2(_01782_),
    .A3(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26212_ (.A1(_01806_),
    .A2(_01838_),
    .B(_01784_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26213_ (.A1(_02200_),
    .A2(_02109_),
    .B(_01685_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26214_ (.A1(_02199_),
    .A2(_02201_),
    .B(_01712_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26215_ (.A1(_02045_),
    .A2(_01696_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26216_ (.A1(_01791_),
    .A2(_01768_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26217_ (.A1(_02106_),
    .A2(_02120_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26218_ (.A1(_02203_),
    .A2(_02204_),
    .A3(_02205_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26219_ (.A1(_01943_),
    .A2(_01730_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26220_ (.A1(_15956_),
    .A2(_01880_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26221_ (.A1(_01719_),
    .A2(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26222_ (.A1(_02209_),
    .A2(_01728_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26223_ (.A1(_02207_),
    .A2(_01845_),
    .A3(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26224_ (.A1(_02206_),
    .A2(_02211_),
    .A3(_01893_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26225_ (.A1(_02212_),
    .A2(_02202_),
    .B(_01739_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26226_ (.A1(_01997_),
    .A2(_01747_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26227_ (.A1(_02214_),
    .A2(_01697_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26228_ (.A1(_01672_),
    .A2(net1137),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26229_ (.A1(_01929_),
    .A2(_01698_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26230_ (.A1(_02216_),
    .A2(_02217_),
    .A3(_01845_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26231_ (.A1(_02215_),
    .A2(_01778_),
    .A3(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26232_ (.A1(_01791_),
    .A2(net590),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26233_ (.A1(_01983_),
    .A2(_01774_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26234_ (.A1(_02220_),
    .A2(_02221_),
    .A3(_01782_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26235_ (.A1(_01983_),
    .A2(_01898_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26236_ (.A1(_02223_),
    .A2(_01811_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26237_ (.A1(_02222_),
    .A2(_01893_),
    .A3(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26238_ (.A1(_02219_),
    .A2(_02225_),
    .A3(_01713_),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26239_ (.A1(_02213_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26240_ (.A1(_02227_),
    .A2(_02196_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26241_ (.A1(_01897_),
    .A2(_02095_),
    .A3(_01718_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26242_ (.A1(_01806_),
    .A2(_01801_),
    .B(_01696_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26243_ (.A1(_01701_),
    .A2(_01880_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26244_ (.A1(_02229_),
    .A2(_02230_),
    .B(_01686_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26245_ (.A1(_02228_),
    .A2(_02231_),
    .B(_01739_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26246_ (.A1(_01837_),
    .A2(_01750_),
    .B(_01773_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26247_ (.A1(_01773_),
    .A2(_15959_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26248_ (.A1(_02233_),
    .A2(_01866_),
    .A3(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26249_ (.A1(_01923_),
    .A2(net1137),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26250_ (.A1(_01750_),
    .A2(_01698_),
    .A3(_01728_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26251_ (.A1(_02236_),
    .A2(_02237_),
    .A3(_01732_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26252_ (.A1(_02235_),
    .A2(_02238_),
    .A3(_01734_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26253_ (.A1(_02232_),
    .A2(_02239_),
    .B(_01849_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26254_ (.A1(_01780_),
    .A2(_01717_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26255_ (.A1(_01983_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26256_ (.A1(_02242_),
    .A2(_02182_),
    .B(_01697_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26257_ (.A1(_01881_),
    .A2(_01773_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26258_ (.A1(_01746_),
    .A2(_02244_),
    .A3(_01866_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26259_ (.A1(_02243_),
    .A2(_01734_),
    .A3(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26260_ (.A1(_01759_),
    .A2(net587),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26261_ (.A1(_02077_),
    .A2(_01807_),
    .B(_01765_),
    .C(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26262_ (.A1(_02241_),
    .A2(_01726_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26263_ (.A1(_01977_),
    .A2(_01911_),
    .A3(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26264_ (.A1(_02248_),
    .A2(_02250_),
    .A3(_01778_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26265_ (.A1(_01739_),
    .A2(_02251_),
    .A3(_02246_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26266_ (.A1(_02252_),
    .A2(_02240_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26267_ (.A1(_01716_),
    .A2(_01701_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26268_ (.A1(_02229_),
    .A2(_02254_),
    .A3(_01757_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26269_ (.A1(_15938_),
    .A2(_01759_),
    .B(_01664_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26270_ (.A1(_02197_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26271_ (.A1(_02255_),
    .A2(_01734_),
    .A3(_02257_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26272_ (.A1(_02241_),
    .A2(_01833_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26273_ (.A1(_02259_),
    .A2(_01732_),
    .A3(_02056_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26274_ (.A1(_01757_),
    .A2(_02208_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26275_ (.A1(_02261_),
    .A2(_01807_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26276_ (.A1(_01831_),
    .A2(_01698_),
    .A3(_01784_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26277_ (.A1(_02262_),
    .A2(_02263_),
    .A3(_01845_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26278_ (.A1(_02260_),
    .A2(_02264_),
    .A3(_01795_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26279_ (.A1(_02258_),
    .A2(_02265_),
    .A3(_01741_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26280_ (.A1(_01923_),
    .A2(_01820_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26281_ (.A1(_02261_),
    .A2(_01701_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26282_ (.A1(_02267_),
    .A2(_02268_),
    .A3(_01765_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26283_ (.A1(_02066_),
    .A2(_01866_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26284_ (.A1(_02270_),
    .A2(_02096_),
    .B(_01685_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26285_ (.A1(_02269_),
    .A2(_02271_),
    .B(_01740_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26286_ (.A1(_01981_),
    .A2(_02207_),
    .A3(_01782_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26287_ (.A1(_02043_),
    .A2(_01855_),
    .A3(_01765_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26288_ (.A1(_02273_),
    .A2(_01893_),
    .A3(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26289_ (.A1(_02272_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26290_ (.A1(_02266_),
    .A2(_02276_),
    .A3(_01849_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26291_ (.A1(_02253_),
    .A2(_02277_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _26292_ (.I(\sa30_sub[7] ),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26293_ (.A1(_02278_),
    .A2(net518),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26294_ (.A1(_11190_),
    .A2(\sa30_sub[7] ),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26295_ (.A1(_02279_),
    .A2(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26296_ (.A1(_02281_),
    .A2(_11158_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26297_ (.A1(_11190_),
    .A2(_02278_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26298_ (.A1(net518),
    .A2(net816),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26299_ (.A1(_02283_),
    .A2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26300_ (.A1(_02285_),
    .A2(\sa30_sub[1] ),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26301_ (.A1(_02282_),
    .A2(_02286_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26302_ (.A1(\sa11_sr[1] ),
    .A2(\sa01_sr[1] ),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26303_ (.A1(_02288_),
    .A2(_14317_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26304_ (.A1(_11215_),
    .A2(_14327_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26305_ (.A1(_02289_),
    .A2(_02290_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26306_ (.A1(_02287_),
    .A2(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26307_ (.A1(_02288_),
    .A2(_14327_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26308_ (.A1(_11215_),
    .A2(_14317_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26309_ (.A1(_02293_),
    .A2(_02294_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26310_ (.A1(_02282_),
    .A2(_02286_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26311_ (.A1(_02295_),
    .A2(_02296_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26312_ (.A1(_02292_),
    .A2(_02297_),
    .B(_12115_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26313_ (.I(\text_in_r[73] ),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26314_ (.A1(_02299_),
    .A2(_10586_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _26315_ (.A1(_02298_),
    .A2(_02300_),
    .B(\u0.w[1][9] ),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26316_ (.A1(_02292_),
    .A2(_02297_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26317_ (.A1(_11348_),
    .A2(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _26318_ (.I(_02300_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26319_ (.A1(net809),
    .A2(_07833_),
    .A3(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26320_ (.A1(_02305_),
    .A2(_02301_),
    .ZN(_15971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26321_ (.A1(_11149_),
    .A2(_11166_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26322_ (.A1(net800),
    .A2(net796),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26323_ (.A1(_02306_),
    .A2(_02307_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26324_ (.A1(_02308_),
    .A2(_14314_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26325_ (.A1(_02306_),
    .A2(_11436_),
    .A3(_02307_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26326_ (.A1(_02309_),
    .A2(_02310_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26327_ (.A1(_02311_),
    .A2(_02285_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26328_ (.A1(_02309_),
    .A2(_02310_),
    .A3(_02281_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26329_ (.A1(_02312_),
    .A2(_02313_),
    .B(_12193_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26330_ (.I(\text_in_r[72] ),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26331_ (.A1(_02315_),
    .A2(_10482_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26332_ (.A1(_02314_),
    .A2(_02316_),
    .B(\u0.w[1][8] ),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26333_ (.A1(_02312_),
    .A2(_02313_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26334_ (.A1(_02318_),
    .A2(_11279_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26335_ (.I(_02316_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26336_ (.A1(_02319_),
    .A2(_07828_),
    .A3(_02320_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26337_ (.A1(_02317_),
    .A2(_02321_),
    .ZN(_15976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26338_ (.A1(_11222_),
    .A2(_11224_),
    .A3(\sa01_sr[2] ),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26339_ (.A1(_11223_),
    .A2(_11221_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26340_ (.A1(\sa11_sr[2] ),
    .A2(\sa30_sub[2] ),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26341_ (.A1(_02323_),
    .A2(_11250_),
    .A3(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26342_ (.A1(_02322_),
    .A2(_02325_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26343_ (.A1(_02326_),
    .A2(net1146),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26344_ (.A1(_02322_),
    .A2(_02325_),
    .A3(net1028),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26345_ (.A1(_02327_),
    .A2(_02328_),
    .B(_10482_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26346_ (.I(\text_in_r[74] ),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26347_ (.A1(_02330_),
    .A2(_11202_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26348_ (.A1(_02329_),
    .A2(_02331_),
    .B(_07839_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26349_ (.A1(_02327_),
    .A2(_02328_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26350_ (.A1(_02333_),
    .A2(_14333_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26351_ (.I(_02331_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26352_ (.A1(_02334_),
    .A2(\u0.w[1][10] ),
    .A3(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26353_ (.A1(_02332_),
    .A2(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26354_ (.I(_02337_),
    .Z(_15992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _26355_ (.A1(_02298_),
    .A2(_02300_),
    .B(_07833_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26356_ (.A1(_02304_),
    .A2(\u0.w[1][9] ),
    .A3(_02303_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26357_ (.A1(_02338_),
    .A2(_02339_),
    .ZN(_15966_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26358_ (.A1(_02329_),
    .A2(_02331_),
    .B(\u0.w[1][10] ),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26359_ (.A1(_02334_),
    .A2(_07839_),
    .A3(_02335_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26360_ (.A1(_02340_),
    .A2(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26361_ (.I(_02342_),
    .Z(_15985_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _26362_ (.I(_02342_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26363_ (.A1(_02343_),
    .A2(_15969_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _26364_ (.I(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26365_ (.A1(_11266_),
    .A2(_14400_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26366_ (.A1(\sa11_sr[3] ),
    .A2(\sa01_sr[3] ),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26367_ (.A1(_02346_),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26368_ (.I(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26369_ (.A1(_11221_),
    .A2(_02278_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26370_ (.A1(\sa30_sub[2] ),
    .A2(net62),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26371_ (.A1(_02350_),
    .A2(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26372_ (.A1(_02349_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26373_ (.I(_02352_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26374_ (.A1(_02354_),
    .A2(_02348_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26375_ (.A1(_02353_),
    .A2(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26376_ (.A1(\sa30_sub[3] ),
    .A2(_14393_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26377_ (.A1(_02356_),
    .A2(_02357_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26378_ (.A1(_11259_),
    .A2(_14393_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26379_ (.A1(_02353_),
    .A2(_02355_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26380_ (.A1(_02359_),
    .A2(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26381_ (.A1(_10522_),
    .A2(_02361_),
    .A3(_02358_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26382_ (.A1(_10525_),
    .A2(\text_in_r[75] ),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26383_ (.A1(_02362_),
    .A2(_02363_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26384_ (.A1(_02364_),
    .A2(\u0.w[1][11] ),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26385_ (.A1(_02362_),
    .A2(_07843_),
    .A3(_02363_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26386_ (.A1(_02365_),
    .A2(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26387_ (.I(_02367_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26388_ (.I(_02368_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26389_ (.A1(\sa30_sub[3] ),
    .A2(net818),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26390_ (.A1(_11342_),
    .A2(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26391_ (.I(_02370_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26392_ (.A1(_02372_),
    .A2(_11341_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26393_ (.A1(_02371_),
    .A2(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26394_ (.I(\sa30_sub[4] ),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26395_ (.A1(_02375_),
    .A2(_14419_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26396_ (.A1(_02374_),
    .A2(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26397_ (.A1(_02374_),
    .A2(_02376_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26398_ (.A1(_02378_),
    .A2(_13010_),
    .A3(_02377_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26399_ (.A1(_11385_),
    .A2(\text_in_r[76] ),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26400_ (.A1(_02379_),
    .A2(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26401_ (.A1(_02381_),
    .A2(_07849_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26402_ (.A1(_02379_),
    .A2(\u0.w[1][12] ),
    .A3(_02380_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26403_ (.A1(_02383_),
    .A2(_02382_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _26404_ (.I(_02384_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26405_ (.A1(_02345_),
    .A2(_02369_),
    .B(net943),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _26406_ (.I(_02337_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26407_ (.A1(_02387_),
    .A2(net797),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26408_ (.A1(_07843_),
    .A2(_02364_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26409_ (.A1(_02362_),
    .A2(\u0.w[1][11] ),
    .A3(_02363_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26410_ (.A1(_02389_),
    .A2(_02390_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26411_ (.I(net70),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26412_ (.A1(_02388_),
    .A2(_02392_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26413_ (.A1(_02316_),
    .A2(_02314_),
    .B(_07828_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26414_ (.A1(_02319_),
    .A2(\u0.w[1][8] ),
    .A3(_02320_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26415_ (.A1(_02395_),
    .A2(_02394_),
    .ZN(_15965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26416_ (.A1(_15965_),
    .A2(_02337_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26417_ (.A1(_02343_),
    .A2(_15981_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _26418_ (.I(_02391_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26419_ (.A1(_02396_),
    .A2(_02397_),
    .A3(_02398_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26420_ (.A1(_02386_),
    .A2(_02393_),
    .A3(_02399_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26421_ (.A1(_15985_),
    .A2(net31),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26422_ (.I(_02401_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26423_ (.I(_02367_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26424_ (.I(_02403_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _26425_ (.I(_02404_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26426_ (.A1(_02337_),
    .A2(_15972_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26427_ (.A1(net810),
    .A2(_02405_),
    .A3(_02406_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _26428_ (.I(_02385_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26429_ (.I(_15983_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26430_ (.A1(_02343_),
    .A2(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26431_ (.I(_02398_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26432_ (.A1(_02396_),
    .A2(_02410_),
    .A3(_02411_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26433_ (.A1(_02407_),
    .A2(_02408_),
    .A3(_02412_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26434_ (.A1(\sa11_sr[6] ),
    .A2(\sa30_sub[6] ),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26435_ (.A1(_14478_),
    .A2(_02414_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26436_ (.A1(_02415_),
    .A2(_11339_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26437_ (.A1(_02415_),
    .A2(_11339_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26438_ (.A1(_10411_),
    .A2(\text_in_r[78] ),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _26439_ (.A1(_02416_),
    .A2(_10526_),
    .A3(_02417_),
    .B(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26440_ (.A1(_02419_),
    .A2(\u0.w[1][14] ),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26441_ (.A1(_02419_),
    .A2(\u0.w[1][14] ),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26442_ (.A1(_02420_),
    .A2(_02421_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26443_ (.A1(_02400_),
    .A2(_02413_),
    .B(_02422_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _26444_ (.I(_15968_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26445_ (.A1(_02342_),
    .A2(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26446_ (.I(_02425_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26447_ (.A1(_02426_),
    .A2(net70),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _26448_ (.I(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26449_ (.A1(_15992_),
    .A2(_15967_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26450_ (.A1(_02428_),
    .A2(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26451_ (.A1(_02343_),
    .A2(_15967_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26452_ (.A1(_02431_),
    .A2(net69),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26453_ (.A1(_02387_),
    .A2(_15977_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26454_ (.A1(_02432_),
    .A2(_02433_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26455_ (.I(_02384_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26456_ (.A1(_02430_),
    .A2(_02434_),
    .B(_02435_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26457_ (.A1(_02387_),
    .A2(_02424_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26458_ (.A1(_02381_),
    .A2(\u0.w[1][12] ),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26459_ (.A1(_02379_),
    .A2(_07849_),
    .A3(_02380_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26460_ (.A1(_02438_),
    .A2(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _26461_ (.I(_02440_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26462_ (.A1(_02392_),
    .A2(_02437_),
    .B(_02441_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26463_ (.A1(net92),
    .A2(_15992_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26464_ (.I(_02403_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26465_ (.A1(_15985_),
    .A2(net802),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26466_ (.A1(_02443_),
    .A2(_02444_),
    .A3(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26467_ (.A1(_02442_),
    .A2(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26468_ (.A1(_02447_),
    .A2(_02422_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26469_ (.A1(_02436_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26470_ (.A1(\sa30_sub[5] ),
    .A2(_11304_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26471_ (.A1(_02450_),
    .A2(_11379_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26472_ (.A1(_02450_),
    .A2(_11379_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26473_ (.A1(_02451_),
    .A2(_02452_),
    .A3(_10405_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26474_ (.A1(_12193_),
    .A2(\text_in_r[77] ),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26475_ (.A1(_02453_),
    .A2(_02454_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26476_ (.A1(_02455_),
    .A2(\u0.w[1][13] ),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26477_ (.A1(_02455_),
    .A2(\u0.w[1][13] ),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26478_ (.A1(_02456_),
    .A2(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26479_ (.I(_02458_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26480_ (.I(_02459_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26481_ (.A1(_02423_),
    .A2(_02449_),
    .B(_02460_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26482_ (.A1(net31),
    .A2(_15965_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26483_ (.A1(_15976_),
    .A2(_02343_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26484_ (.A1(_02462_),
    .A2(_02463_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26485_ (.A1(_02464_),
    .A2(_02392_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26486_ (.A1(_02463_),
    .A2(net69),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26487_ (.I(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26488_ (.A1(_02467_),
    .A2(_02462_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26489_ (.I(_02385_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26490_ (.A1(_02465_),
    .A2(_02468_),
    .A3(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26491_ (.A1(_02387_),
    .A2(_15981_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26492_ (.A1(_02471_),
    .A2(_02403_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26493_ (.A1(_02472_),
    .A2(net66),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26494_ (.I(_02441_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26495_ (.A1(_15985_),
    .A2(_15977_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26496_ (.A1(_02429_),
    .A2(_02475_),
    .A3(_02411_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26497_ (.A1(_02473_),
    .A2(_02474_),
    .A3(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26498_ (.I(_02422_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26499_ (.A1(_02470_),
    .A2(_02477_),
    .A3(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26500_ (.A1(net794),
    .A2(_02343_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26501_ (.A1(_02480_),
    .A2(_02406_),
    .A3(_02369_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26502_ (.A1(_02409_),
    .A2(_02387_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _26503_ (.I(_02398_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26504_ (.A1(net66),
    .A2(_02482_),
    .A3(_02483_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _26505_ (.I(_02441_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26506_ (.A1(_02481_),
    .A2(_02484_),
    .B(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _26507_ (.I(_15974_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26508_ (.A1(_02343_),
    .A2(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26509_ (.A1(_02488_),
    .A2(_02406_),
    .A3(_02411_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26510_ (.A1(_02396_),
    .A2(net69),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26511_ (.I(_02384_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26512_ (.A1(_02489_),
    .A2(_02490_),
    .B(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _26513_ (.I(_02422_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26514_ (.I(_02493_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26515_ (.A1(_02486_),
    .A2(_02492_),
    .B(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _26516_ (.I(_02458_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26517_ (.I(_02496_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26518_ (.I(_02497_),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26519_ (.A1(_02479_),
    .A2(_02495_),
    .A3(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _26520_ (.A1(net819),
    .A2(_11189_),
    .A3(_11382_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26521_ (.A1(_12961_),
    .A2(\text_in_r[79] ),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26522_ (.A1(_02500_),
    .A2(_12965_),
    .B(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _26523_ (.A1(\u0.w[1][15] ),
    .A2(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26524_ (.I(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26525_ (.A1(_02461_),
    .A2(_02499_),
    .A3(_02504_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26526_ (.A1(_15971_),
    .A2(_02343_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26527_ (.A1(_02506_),
    .A2(_02403_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26528_ (.A1(_02387_),
    .A2(net801),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26529_ (.A1(_02507_),
    .A2(_02508_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26530_ (.A1(_02480_),
    .A2(_02433_),
    .A3(_02411_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26531_ (.A1(_02509_),
    .A2(_02510_),
    .B(_02435_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26532_ (.I(_15967_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26533_ (.A1(_15992_),
    .A2(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26534_ (.A1(_02513_),
    .A2(_02345_),
    .B(_02444_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26535_ (.A1(_02488_),
    .A2(_02391_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26536_ (.I(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _26537_ (.I(_02441_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26538_ (.A1(_02514_),
    .A2(_02516_),
    .B(_02517_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26539_ (.A1(_02511_),
    .A2(_02518_),
    .B(_02494_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26540_ (.A1(_02345_),
    .A2(_02398_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26541_ (.A1(_02520_),
    .A2(_02384_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26542_ (.A1(_02343_),
    .A2(_15972_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26543_ (.A1(_02433_),
    .A2(_02522_),
    .A3(_02369_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26544_ (.A1(_02521_),
    .A2(_02523_),
    .B(_02493_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26545_ (.A1(_02522_),
    .A2(net70),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26546_ (.I(_15979_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26547_ (.A1(_02387_),
    .A2(_02526_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26548_ (.A1(_02525_),
    .A2(_02527_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26549_ (.A1(_02345_),
    .A2(_02405_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26550_ (.A1(_02528_),
    .A2(_02474_),
    .A3(_02529_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26551_ (.I(_02458_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26552_ (.A1(_02524_),
    .A2(_02530_),
    .B(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26553_ (.A1(_02519_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26554_ (.A1(_02387_),
    .A2(_15974_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26555_ (.I(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26556_ (.A1(_02535_),
    .A2(_02368_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26557_ (.A1(_02399_),
    .A2(_02441_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26558_ (.A1(_02343_),
    .A2(_15979_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26559_ (.A1(_02534_),
    .A2(_02538_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26560_ (.A1(_02539_),
    .A2(_02444_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26561_ (.A1(_02540_),
    .A2(_02491_),
    .A3(_02427_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26562_ (.A1(_02536_),
    .A2(_02537_),
    .B(_02541_),
    .C(_02494_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _26563_ (.I(_02508_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26564_ (.A1(_02543_),
    .A2(_02444_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26565_ (.A1(_02392_),
    .A2(_15990_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26566_ (.A1(_02544_),
    .A2(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26567_ (.A1(_02546_),
    .A2(_02408_),
    .B(_02493_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26568_ (.I(_15972_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26569_ (.A1(_02548_),
    .A2(_15985_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26570_ (.A1(_02549_),
    .A2(_02398_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26571_ (.A1(_02550_),
    .A2(_02441_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26572_ (.A1(_02551_),
    .A2(_02536_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26573_ (.A1(_02396_),
    .A2(_02431_),
    .A3(_02398_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26574_ (.A1(_15992_),
    .A2(_15969_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26575_ (.A1(_02554_),
    .A2(_02398_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26576_ (.A1(_02553_),
    .A2(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26577_ (.A1(_02552_),
    .A2(_02556_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26578_ (.I(_02496_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26579_ (.A1(_02547_),
    .A2(_02557_),
    .B(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26580_ (.A1(_02542_),
    .A2(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _26581_ (.I(_02503_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26582_ (.A1(_02533_),
    .A2(_02560_),
    .A3(_02561_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26583_ (.A1(_02505_),
    .A2(_02562_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26584_ (.A1(_02515_),
    .A2(_02388_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26585_ (.A1(_02463_),
    .A2(_02429_),
    .A3(_02369_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26586_ (.A1(_02563_),
    .A2(_02474_),
    .A3(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26587_ (.A1(_15976_),
    .A2(_02387_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26588_ (.A1(_02566_),
    .A2(_02344_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26589_ (.I(_02404_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26590_ (.A1(_02567_),
    .A2(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26591_ (.A1(_02431_),
    .A2(_02437_),
    .A3(_02411_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26592_ (.A1(_02569_),
    .A2(_02570_),
    .A3(_02435_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26593_ (.A1(_02565_),
    .A2(_02571_),
    .A3(_02558_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26594_ (.A1(_02471_),
    .A2(_02398_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26595_ (.A1(_02573_),
    .A2(_02445_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26596_ (.I(_15969_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26597_ (.A1(_02387_),
    .A2(_02575_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26598_ (.A1(_02410_),
    .A2(_02576_),
    .A3(_02369_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26599_ (.A1(_02574_),
    .A2(_02408_),
    .A3(_02577_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26600_ (.A1(_02396_),
    .A2(_02397_),
    .A3(_02369_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26601_ (.A1(_02579_),
    .A2(_02517_),
    .A3(_02427_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26602_ (.A1(_02578_),
    .A2(_02531_),
    .A3(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26603_ (.A1(_02572_),
    .A2(_02581_),
    .B(_02478_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26604_ (.A1(_02480_),
    .A2(_02368_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26605_ (.A1(_02583_),
    .A2(_02429_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26606_ (.A1(_02406_),
    .A2(net820),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26607_ (.I(_02585_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26608_ (.A1(_02586_),
    .A2(_02397_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26609_ (.A1(_02584_),
    .A2(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26610_ (.I(_02440_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26611_ (.I(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26612_ (.A1(_02588_),
    .A2(_02558_),
    .B(_02590_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26613_ (.A1(_02467_),
    .A2(_02443_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26614_ (.A1(_02592_),
    .A2(_02563_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26615_ (.A1(_02593_),
    .A2(_02460_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26616_ (.I(_15993_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26617_ (.A1(_02458_),
    .A2(_02595_),
    .A3(_02411_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26618_ (.A1(_02397_),
    .A2(_02403_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26619_ (.A1(_02597_),
    .A2(_02433_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26620_ (.A1(_02596_),
    .A2(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26621_ (.A1(_02599_),
    .A2(_02469_),
    .B(_02422_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26622_ (.A1(_02591_),
    .A2(_02594_),
    .B(_02600_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26623_ (.A1(_02582_),
    .A2(_02601_),
    .B(_02504_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26624_ (.A1(_02507_),
    .A2(_02462_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _26625_ (.I(_02391_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26626_ (.A1(_02604_),
    .A2(_15992_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26627_ (.A1(_02605_),
    .A2(_02548_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26628_ (.A1(_02603_),
    .A2(_02590_),
    .A3(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26629_ (.A1(_02488_),
    .A2(net69),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26630_ (.I(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26631_ (.A1(_02609_),
    .A2(_02566_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26632_ (.A1(_02428_),
    .A2(_02396_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26633_ (.A1(_02610_),
    .A2(_02611_),
    .A3(_02408_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26634_ (.A1(_02607_),
    .A2(_02612_),
    .A3(_02498_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26635_ (.A1(_02535_),
    .A2(_02369_),
    .B(_02589_),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26636_ (.A1(_02401_),
    .A2(_02483_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26637_ (.A1(_02368_),
    .A2(_15997_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26638_ (.A1(_02614_),
    .A2(_02615_),
    .A3(_02616_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26639_ (.A1(_02534_),
    .A2(net944),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26640_ (.A1(_02618_),
    .A2(_02568_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26641_ (.A1(_02437_),
    .A2(_02410_),
    .A3(_02483_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26642_ (.A1(_02619_),
    .A2(_02620_),
    .A3(_02517_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26643_ (.A1(_02617_),
    .A2(_02621_),
    .A3(_02531_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26644_ (.A1(_02613_),
    .A2(_02478_),
    .A3(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26645_ (.A1(net92),
    .A2(_15976_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26646_ (.A1(_02624_),
    .A2(_02480_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26647_ (.I(_02604_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26648_ (.A1(_02625_),
    .A2(_02626_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26649_ (.A1(_02508_),
    .A2(_02404_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26650_ (.A1(_02628_),
    .A2(_02480_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26651_ (.A1(_02627_),
    .A2(_02629_),
    .A3(_02517_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26652_ (.A1(_02534_),
    .A2(net66),
    .A3(_02392_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26653_ (.A1(_15985_),
    .A2(_02512_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26654_ (.A1(_02566_),
    .A2(_02632_),
    .A3(_02444_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26655_ (.A1(_02631_),
    .A2(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26656_ (.A1(_02634_),
    .A2(_02469_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26657_ (.A1(_02630_),
    .A2(_02635_),
    .A3(_02531_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _26658_ (.I(_02493_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26659_ (.A1(_15985_),
    .A2(_15974_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26660_ (.A1(_02638_),
    .A2(_02369_),
    .B(net943),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26661_ (.A1(_02639_),
    .A2(_02574_),
    .B(_02459_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26662_ (.A1(_02482_),
    .A2(net70),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26663_ (.A1(_02641_),
    .A2(_02402_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _26664_ (.I(_15981_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26665_ (.A1(_15985_),
    .A2(_02643_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26666_ (.I(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26667_ (.A1(_02645_),
    .A2(_02405_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26668_ (.A1(_02642_),
    .A2(_02435_),
    .A3(_02646_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26669_ (.A1(_02640_),
    .A2(_02647_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26670_ (.A1(_02636_),
    .A2(_02637_),
    .A3(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26671_ (.A1(_02623_),
    .A2(_02649_),
    .A3(_02561_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26672_ (.A1(_02602_),
    .A2(_02650_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26673_ (.A1(net944),
    .A2(_02398_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26674_ (.A1(_02651_),
    .A2(_02534_),
    .B(net943),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26675_ (.A1(_02652_),
    .A2(_02509_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26676_ (.I(_02506_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26677_ (.A1(_02654_),
    .A2(_02585_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26678_ (.I(_02482_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26679_ (.A1(_02608_),
    .A2(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26680_ (.A1(_02655_),
    .A2(_02657_),
    .B(_02491_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26681_ (.A1(_02653_),
    .A2(_02658_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26682_ (.A1(_02659_),
    .A2(_02460_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26683_ (.A1(_02388_),
    .A2(_02444_),
    .A3(_02445_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26684_ (.I(_02661_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26685_ (.A1(_02463_),
    .A2(_02554_),
    .A3(_02392_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26686_ (.A1(_02662_),
    .A2(_02663_),
    .B(_02469_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26687_ (.A1(_02406_),
    .A2(_02404_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26688_ (.A1(_02665_),
    .A2(_02589_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26689_ (.A1(_02573_),
    .A2(_02410_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26690_ (.A1(_02666_),
    .A2(_02667_),
    .B(_02459_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26691_ (.A1(_02664_),
    .A2(_02668_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26692_ (.A1(_02660_),
    .A2(_02478_),
    .A3(_02669_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26693_ (.A1(_15992_),
    .A2(_15983_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26694_ (.I(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26695_ (.A1(_02466_),
    .A2(_02672_),
    .B(_02384_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26696_ (.A1(_02388_),
    .A2(_02392_),
    .A3(_02538_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26697_ (.A1(_02673_),
    .A2(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26698_ (.A1(_02426_),
    .A2(_02508_),
    .A3(_02392_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26699_ (.A1(_02480_),
    .A2(_02527_),
    .A3(_02404_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26700_ (.A1(_02676_),
    .A2(_02677_),
    .B(_02435_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26701_ (.A1(_02675_),
    .A2(_02678_),
    .B(_02498_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26702_ (.A1(_15992_),
    .A2(_02487_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26703_ (.A1(_02680_),
    .A2(_02604_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26704_ (.A1(_02681_),
    .A2(net810),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26705_ (.A1(_02682_),
    .A2(_02474_),
    .A3(_02540_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26706_ (.A1(_02534_),
    .A2(_02392_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26707_ (.I(_02463_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26708_ (.A1(_02671_),
    .A2(_02368_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26709_ (.A1(_02684_),
    .A2(_02685_),
    .B(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26710_ (.I(_02538_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26711_ (.A1(_02688_),
    .A2(_02404_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26712_ (.A1(_02689_),
    .A2(_02485_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26713_ (.A1(_02687_),
    .A2(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26714_ (.A1(_02683_),
    .A2(_02691_),
    .A3(_02531_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26715_ (.A1(_02679_),
    .A2(_02692_),
    .A3(_02637_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26716_ (.A1(_02670_),
    .A2(_02693_),
    .A3(_02504_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26717_ (.A1(_02632_),
    .A2(_02398_),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26718_ (.A1(_02695_),
    .A2(_02589_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26719_ (.A1(_02428_),
    .A2(_02680_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26720_ (.A1(_02697_),
    .A2(_02696_),
    .B(_02459_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26721_ (.A1(_02575_),
    .A2(_02487_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26722_ (.A1(_15985_),
    .A2(_02699_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26723_ (.A1(_02573_),
    .A2(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26724_ (.A1(_02598_),
    .A2(_02701_),
    .A3(_02435_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26725_ (.A1(_02698_),
    .A2(_02702_),
    .B(_02494_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26726_ (.A1(_02404_),
    .A2(_15999_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26727_ (.A1(_02655_),
    .A2(_02485_),
    .A3(_02704_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26728_ (.A1(_02368_),
    .A2(_15988_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26729_ (.A1(_02706_),
    .A2(_02665_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26730_ (.I(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26731_ (.A1(_02708_),
    .A2(_02474_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26732_ (.A1(_02705_),
    .A2(_02531_),
    .A3(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26733_ (.A1(_02710_),
    .A2(_02703_),
    .B(_02504_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26734_ (.A1(_02506_),
    .A2(_02462_),
    .A3(_02483_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26735_ (.A1(_15993_),
    .A2(_02626_),
    .B(_02712_),
    .C(_02517_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26736_ (.I(_02513_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26737_ (.A1(_02507_),
    .A2(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26738_ (.A1(_02508_),
    .A2(_02604_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26739_ (.I(_15977_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26740_ (.A1(_15985_),
    .A2(_02717_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26741_ (.A1(_02716_),
    .A2(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26742_ (.A1(_02715_),
    .A2(_02719_),
    .B(_02408_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26743_ (.A1(_02713_),
    .A2(_02720_),
    .A3(_02460_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26744_ (.A1(_02388_),
    .A2(_02483_),
    .A3(_02480_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26745_ (.A1(_02509_),
    .A2(_02469_),
    .A3(_02722_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26746_ (.A1(_15990_),
    .A2(_02405_),
    .B(_02491_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26747_ (.A1(_02525_),
    .A2(_02437_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26748_ (.A1(_02724_),
    .A2(_02725_),
    .B(_02459_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26749_ (.A1(_02723_),
    .A2(_02726_),
    .B(_02422_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26750_ (.A1(_02721_),
    .A2(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26751_ (.A1(_02711_),
    .A2(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26752_ (.A1(_02694_),
    .A2(_02729_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26753_ (.A1(_02586_),
    .A2(_02475_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26754_ (.A1(_02597_),
    .A2(_02437_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26755_ (.A1(_02730_),
    .A2(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26756_ (.A1(_02732_),
    .A2(_02485_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26757_ (.A1(_02426_),
    .A2(_02368_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26758_ (.A1(_15992_),
    .A2(_02717_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26759_ (.A1(_02734_),
    .A2(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26760_ (.A1(_02465_),
    .A2(_02736_),
    .A3(_02491_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26761_ (.A1(_02733_),
    .A2(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26762_ (.A1(_02738_),
    .A2(_02637_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26763_ (.A1(_02681_),
    .A2(_02410_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26764_ (.A1(_02740_),
    .A2(_02661_),
    .A3(_02474_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26765_ (.I(_02566_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26766_ (.A1(_02742_),
    .A2(_02718_),
    .B(_02405_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26767_ (.A1(_02632_),
    .A2(_02437_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26768_ (.A1(_02744_),
    .A2(_02626_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26769_ (.A1(_02743_),
    .A2(_02408_),
    .A3(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26770_ (.A1(_02741_),
    .A2(_02746_),
    .A3(_02422_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26771_ (.A1(_02739_),
    .A2(_02498_),
    .A3(_02747_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26772_ (.A1(net803),
    .A2(_02405_),
    .A3(_02480_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26773_ (.A1(_02442_),
    .A2(_02749_),
    .B(_02494_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26774_ (.A1(_02462_),
    .A2(_02566_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26775_ (.A1(_02751_),
    .A2(_02405_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26776_ (.A1(_02388_),
    .A2(_02626_),
    .A3(net66),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26777_ (.A1(_02752_),
    .A2(_02753_),
    .A3(_02474_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26778_ (.A1(_02750_),
    .A2(_02754_),
    .B(_02558_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26779_ (.A1(_02527_),
    .A2(_02368_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26780_ (.A1(_02756_),
    .A2(_02445_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26781_ (.A1(_02642_),
    .A2(_02757_),
    .A3(_02469_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26782_ (.A1(_02752_),
    .A2(_02590_),
    .A3(_02585_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26783_ (.A1(_02758_),
    .A2(_02759_),
    .A3(_02637_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26784_ (.A1(_02755_),
    .A2(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26785_ (.A1(_02748_),
    .A2(_02761_),
    .A3(_02561_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26786_ (.A1(_02553_),
    .A2(_02441_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26787_ (.A1(_02763_),
    .A2(_02603_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26788_ (.A1(_02734_),
    .A2(_02482_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26789_ (.A1(_02396_),
    .A2(_02538_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26790_ (.A1(_02766_),
    .A2(_02604_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26791_ (.A1(_02765_),
    .A2(net943),
    .A3(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26792_ (.A1(_02768_),
    .A2(_02764_),
    .B(_02558_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26793_ (.A1(_02673_),
    .A2(_02458_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26794_ (.A1(_02527_),
    .A2(_02391_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26795_ (.A1(_02771_),
    .A2(_02700_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26796_ (.A1(_02598_),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26797_ (.A1(_02773_),
    .A2(_02485_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26798_ (.A1(_02770_),
    .A2(_02774_),
    .B(_02422_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26799_ (.A1(_02775_),
    .A2(_02769_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26800_ (.A1(_02433_),
    .A2(_02368_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _26801_ (.A1(_02496_),
    .A2(_02654_),
    .A3(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26802_ (.I(_02425_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26803_ (.A1(_02779_),
    .A2(_02368_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26804_ (.A1(_02780_),
    .A2(_02496_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26805_ (.A1(_02778_),
    .A2(_02781_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26806_ (.I(_02521_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26807_ (.I(_02437_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26808_ (.A1(_02458_),
    .A2(_02604_),
    .A3(_02784_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26809_ (.A1(_02783_),
    .A2(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26810_ (.A1(_02782_),
    .A2(_02786_),
    .B(_02494_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26811_ (.I(_02490_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26812_ (.A1(_02788_),
    .A2(_02426_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26813_ (.A1(_02641_),
    .A2(_02700_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26814_ (.A1(_02789_),
    .A2(_02790_),
    .A3(_02458_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26815_ (.A1(_02688_),
    .A2(_02604_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26816_ (.A1(_02677_),
    .A2(_02496_),
    .A3(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26817_ (.A1(_02791_),
    .A2(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26818_ (.A1(_02794_),
    .A2(_02590_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26819_ (.A1(_02787_),
    .A2(_02795_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26820_ (.A1(_02796_),
    .A2(_02776_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26821_ (.A1(_02797_),
    .A2(_02504_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26822_ (.A1(_02798_),
    .A2(_02762_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26823_ (.A1(_02388_),
    .A2(_02463_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26824_ (.A1(_02799_),
    .A2(_02626_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26825_ (.A1(_02800_),
    .A2(_02584_),
    .A3(_02590_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26826_ (.A1(_02771_),
    .A2(_02485_),
    .A3(_02345_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26827_ (.A1(_02801_),
    .A2(_02498_),
    .A3(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26828_ (.A1(_02592_),
    .A2(_02712_),
    .A3(_02590_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26829_ (.A1(_02402_),
    .A2(_02624_),
    .A3(_02405_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26830_ (.A1(_02402_),
    .A2(_02411_),
    .A3(_02429_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26831_ (.A1(_02805_),
    .A2(_02806_),
    .A3(_02408_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26832_ (.A1(_02804_),
    .A2(_02807_),
    .A3(_02460_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26833_ (.A1(_02803_),
    .A2(_02808_),
    .A3(_02637_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26834_ (.A1(net803),
    .A2(_02626_),
    .A3(_02431_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26835_ (.A1(_02552_),
    .A2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26836_ (.I(_02657_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26837_ (.A1(_02525_),
    .A2(net803),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26838_ (.A1(_02812_),
    .A2(_02813_),
    .A3(_02408_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26839_ (.A1(_02811_),
    .A2(_02814_),
    .A3(_02460_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26840_ (.A1(_02688_),
    .A2(_02483_),
    .B(_02589_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26841_ (.A1(_02543_),
    .A2(_02604_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26842_ (.I(_02817_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26843_ (.A1(_02816_),
    .A2(_02818_),
    .A3(_02540_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26844_ (.A1(_02437_),
    .A2(_02410_),
    .A3(_02369_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26845_ (.A1(_02528_),
    .A2(_02517_),
    .A3(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26846_ (.A1(_02819_),
    .A2(_02821_),
    .A3(_02558_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26847_ (.A1(_02815_),
    .A2(_02822_),
    .A3(_02478_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26848_ (.A1(_02809_),
    .A2(_02823_),
    .A3(_02561_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26849_ (.A1(_02467_),
    .A2(_02482_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26850_ (.A1(_02825_),
    .A2(_02605_),
    .B(_02485_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26851_ (.A1(_02432_),
    .A2(_02443_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26852_ (.I(_02563_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26853_ (.A1(_02827_),
    .A2(_02828_),
    .B(_02491_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26854_ (.A1(_02826_),
    .A2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26855_ (.A1(_02830_),
    .A2(_02637_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26856_ (.A1(_02401_),
    .A2(_02624_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26857_ (.A1(_02832_),
    .A2(_02444_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26858_ (.A1(_02771_),
    .A2(_02463_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26859_ (.A1(_02833_),
    .A2(_02834_),
    .B(_02517_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26860_ (.A1(_02465_),
    .A2(_02514_),
    .B(_02435_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26861_ (.A1(_02835_),
    .A2(_02836_),
    .B(_02478_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26862_ (.A1(_02831_),
    .A2(_02837_),
    .A3(_02460_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26863_ (.A1(_02404_),
    .A2(_02643_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26864_ (.A1(_02716_),
    .A2(_02839_),
    .A3(_02441_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26865_ (.A1(_02840_),
    .A2(_02494_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26866_ (.A1(_02550_),
    .A2(_02385_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26867_ (.A1(_02771_),
    .A2(_02402_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26868_ (.A1(_02842_),
    .A2(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26869_ (.A1(_02841_),
    .A2(_02844_),
    .B(_02531_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26870_ (.A1(_02609_),
    .A2(_02508_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26871_ (.A1(_02537_),
    .A2(_02846_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26872_ (.A1(_02576_),
    .A2(net69),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26873_ (.I(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26874_ (.A1(_02849_),
    .A2(_02573_),
    .A3(_02589_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26875_ (.A1(_02847_),
    .A2(_02850_),
    .A3(_02494_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26876_ (.A1(_02845_),
    .A2(_02851_),
    .B(_02561_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26877_ (.A1(_02838_),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26878_ (.A1(_02824_),
    .A2(_02853_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26879_ (.A1(_02426_),
    .A2(_02671_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _26880_ (.A1(_02428_),
    .A2(_02433_),
    .B1(_02854_),
    .B2(_02568_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26881_ (.A1(_02855_),
    .A2(_02469_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26882_ (.A1(_02604_),
    .A2(_02717_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _26883_ (.A1(_02597_),
    .A2(_02857_),
    .A3(_02491_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26884_ (.A1(_02858_),
    .A2(_02558_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26885_ (.A1(_02856_),
    .A2(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26886_ (.A1(_02597_),
    .A2(_02406_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26887_ (.A1(_02700_),
    .A2(_02626_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26888_ (.A1(_02861_),
    .A2(_02474_),
    .A3(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26889_ (.I(_02641_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26890_ (.A1(_02614_),
    .A2(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26891_ (.A1(_02863_),
    .A2(_02498_),
    .A3(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26892_ (.A1(_02860_),
    .A2(_02504_),
    .A3(_02866_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26893_ (.A1(_02849_),
    .A2(_02506_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26894_ (.A1(_02868_),
    .A2(_02817_),
    .B(_02491_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26895_ (.A1(_02686_),
    .A2(_02441_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26896_ (.A1(_02428_),
    .A2(_02714_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26897_ (.A1(_02870_),
    .A2(_02871_),
    .B(_02497_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26898_ (.A1(_02869_),
    .A2(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26899_ (.A1(net31),
    .A2(_02483_),
    .B(_02385_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26900_ (.A1(_02833_),
    .A2(_02874_),
    .B(_02459_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26901_ (.A1(_02788_),
    .A2(_02624_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26902_ (.A1(_02644_),
    .A2(_02735_),
    .A3(_02483_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26903_ (.A1(_02876_),
    .A2(_02877_),
    .A3(_02491_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26904_ (.A1(_02875_),
    .A2(_02878_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26905_ (.A1(_02873_),
    .A2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26906_ (.A1(_02880_),
    .A2(_02561_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26907_ (.A1(_02867_),
    .A2(_02881_),
    .A3(_02478_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26908_ (.A1(_15992_),
    .A2(_02548_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26909_ (.A1(_02608_),
    .A2(net943),
    .A3(_02883_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26910_ (.A1(_02884_),
    .A2(_02497_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26911_ (.A1(net66),
    .A2(_02444_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26912_ (.A1(_02767_),
    .A2(_02517_),
    .A3(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26913_ (.A1(_02885_),
    .A2(_02887_),
    .B(_02504_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26914_ (.A1(_02756_),
    .A2(_02522_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26915_ (.I(_02699_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26916_ (.A1(_02681_),
    .A2(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26917_ (.A1(_02889_),
    .A2(_02891_),
    .A3(_02408_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26918_ (.A1(_02641_),
    .A2(_02488_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26919_ (.A1(_02386_),
    .A2(_02893_),
    .A3(_02393_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26920_ (.A1(_02892_),
    .A2(_02894_),
    .A3(_02498_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26921_ (.A1(_02888_),
    .A2(_02895_),
    .B(_02478_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26922_ (.A1(_15965_),
    .A2(_02568_),
    .B(_02468_),
    .C(_02517_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26923_ (.A1(_02756_),
    .A2(_02402_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26924_ (.A1(_02779_),
    .A2(_02585_),
    .B(_02898_),
    .C(_02435_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26925_ (.A1(_02897_),
    .A2(_02899_),
    .A3(_02498_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26926_ (.A1(_02605_),
    .A2(_02717_),
    .B(_02589_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26927_ (.A1(_02597_),
    .A2(_02482_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26928_ (.A1(_02901_),
    .A2(_02902_),
    .B(_02497_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26929_ (.A1(_02583_),
    .A2(_02680_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26930_ (.A1(_02904_),
    .A2(_02537_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26931_ (.A1(_02903_),
    .A2(_02905_),
    .B(_02561_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26932_ (.A1(_02900_),
    .A2(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26933_ (.A1(_02896_),
    .A2(_02907_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26934_ (.A1(_02882_),
    .A2(_02908_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26935_ (.A1(_02520_),
    .A2(_02589_),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26936_ (.A1(_02756_),
    .A2(_02410_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26937_ (.A1(_02605_),
    .A2(_02643_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26938_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26939_ (.A1(_02628_),
    .A2(_02463_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26940_ (.A1(_02605_),
    .A2(_02890_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26941_ (.A1(_02816_),
    .A2(_02913_),
    .A3(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26942_ (.A1(_02912_),
    .A2(_02915_),
    .A3(_02460_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26943_ (.A1(_02832_),
    .A2(_02626_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26944_ (.A1(_15986_),
    .A2(_15995_),
    .B(_02405_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26945_ (.A1(_02917_),
    .A2(_02590_),
    .A3(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26946_ (.A1(_02605_),
    .A2(_15969_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26947_ (.A1(_02816_),
    .A2(_02920_),
    .A3(_02695_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26948_ (.A1(_02919_),
    .A2(_02921_),
    .A3(_02498_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26949_ (.A1(_02916_),
    .A2(_02922_),
    .A3(_02637_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26950_ (.A1(_02849_),
    .A2(_02445_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26951_ (.A1(_02586_),
    .A2(net810),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26952_ (.A1(_02924_),
    .A2(_02925_),
    .A3(_02497_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26953_ (.A1(_02628_),
    .A2(_02700_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26954_ (.A1(_02525_),
    .A2(_02566_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26955_ (.A1(_02927_),
    .A2(_02928_),
    .A3(_02531_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26956_ (.A1(_02926_),
    .A2(_02929_),
    .A3(_02590_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26957_ (.A1(_02443_),
    .A2(_02626_),
    .A3(_02522_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26958_ (.A1(_02735_),
    .A2(_02483_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26959_ (.A1(_02931_),
    .A2(_02531_),
    .A3(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26960_ (.A1(_02708_),
    .A2(_02558_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26961_ (.A1(_02780_),
    .A2(_02497_),
    .B(_02485_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26962_ (.A1(_02933_),
    .A2(_02934_),
    .A3(_02935_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26963_ (.A1(_02930_),
    .A2(_02936_),
    .A3(_02478_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26964_ (.A1(_02923_),
    .A2(_02937_),
    .A3(_02561_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26965_ (.I(_02445_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _26966_ (.A1(_02939_),
    .A2(_02405_),
    .B1(_02456_),
    .B2(_02457_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26967_ (.A1(_02940_),
    .A2(_02767_),
    .B(_02408_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26968_ (.A1(_02751_),
    .A2(_02404_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26969_ (.A1(net810),
    .A2(_02444_),
    .A3(_02883_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26970_ (.A1(_02942_),
    .A2(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26971_ (.A1(_02944_),
    .A2(_02558_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26972_ (.A1(_02941_),
    .A2(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26973_ (.A1(_02616_),
    .A2(_02458_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26974_ (.A1(_02947_),
    .A2(_02481_),
    .B(_02517_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26975_ (.A1(_02410_),
    .A2(_02404_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26976_ (.A1(_02949_),
    .A2(_02742_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26977_ (.A1(_02942_),
    .A2(_02497_),
    .A3(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26978_ (.A1(_02948_),
    .A2(_02951_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26979_ (.A1(_02946_),
    .A2(_02952_),
    .A3(_02637_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26980_ (.I(_15987_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26981_ (.A1(_02954_),
    .A2(_02411_),
    .B(_02491_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26982_ (.A1(_02955_),
    .A2(_02898_),
    .B(_02459_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26983_ (.A1(_02742_),
    .A2(_02568_),
    .B(_02589_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26984_ (.A1(_02854_),
    .A2(_02626_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26985_ (.A1(_02957_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26986_ (.A1(_02956_),
    .A2(_02959_),
    .B(_02494_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26987_ (.A1(_02843_),
    .A2(_02777_),
    .B(_02485_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26988_ (.A1(_02961_),
    .A2(_02652_),
    .B(_02531_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26989_ (.A1(_02960_),
    .A2(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26990_ (.A1(_02953_),
    .A2(_02963_),
    .A3(_02504_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26991_ (.A1(_02938_),
    .A2(_02964_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26992_ (.A1(_02568_),
    .A2(_15976_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26993_ (.A1(_02799_),
    .A2(_02568_),
    .B(_02435_),
    .C(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26994_ (.A1(_02472_),
    .A2(net810),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26995_ (.A1(_02712_),
    .A2(_02967_),
    .A3(_02590_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26996_ (.A1(_02966_),
    .A2(_02968_),
    .A3(_02498_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26997_ (.A1(_02568_),
    .A2(_02645_),
    .B(_02886_),
    .C(_02485_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26998_ (.A1(_02525_),
    .A2(_02472_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26999_ (.A1(_02939_),
    .A2(_02444_),
    .B(_02441_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27000_ (.A1(_02971_),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27001_ (.A1(_02970_),
    .A2(_02973_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27002_ (.A1(_02974_),
    .A2(_02460_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27003_ (.A1(_02969_),
    .A2(_02975_),
    .A3(_02478_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27004_ (.A1(_02789_),
    .A2(_02469_),
    .A3(_02620_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27005_ (.A1(_02910_),
    .A2(_02722_),
    .A3(_02474_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27006_ (.A1(_02977_),
    .A2(_02978_),
    .A3(_02460_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27007_ (.A1(_02843_),
    .A2(_02474_),
    .A3(_02949_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27008_ (.A1(_02396_),
    .A2(_02522_),
    .A3(_02369_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27009_ (.A1(_02431_),
    .A2(_02471_),
    .A3(_02483_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27010_ (.A1(_02981_),
    .A2(_02982_),
    .A3(_02435_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27011_ (.A1(_02980_),
    .A2(_02983_),
    .A3(_02558_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27012_ (.A1(_02979_),
    .A2(_02637_),
    .A3(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27013_ (.A1(_02976_),
    .A2(_02985_),
    .A3(_02504_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27014_ (.A1(_02443_),
    .A2(_02392_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27015_ (.A1(_02987_),
    .A2(_02848_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27016_ (.A1(_02988_),
    .A2(_02459_),
    .A3(_02431_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27017_ (.A1(_02432_),
    .A2(_02471_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27018_ (.A1(_02433_),
    .A2(_02445_),
    .A3(_02411_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27019_ (.A1(_02990_),
    .A2(_02991_),
    .B(_02459_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27020_ (.A1(_02989_),
    .A2(_02992_),
    .B(_02590_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27021_ (.A1(_15974_),
    .A2(_02568_),
    .B(_02497_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27022_ (.A1(_02994_),
    .A2(_02917_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27023_ (.A1(_02472_),
    .A2(_02506_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27024_ (.A1(_02772_),
    .A2(_02996_),
    .A3(_02497_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27025_ (.A1(_02995_),
    .A2(_02997_),
    .A3(_02469_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27026_ (.A1(_02993_),
    .A2(_02637_),
    .A3(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27027_ (.A1(_02842_),
    .A2(_02393_),
    .A3(_02563_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27028_ (.A1(_02643_),
    .A2(_02411_),
    .B(_02385_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27029_ (.A1(_03001_),
    .A2(_02555_),
    .B(_02459_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27030_ (.A1(_03000_),
    .A2(_03002_),
    .B(_02494_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27031_ (.A1(_02507_),
    .A2(_02566_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27032_ (.A1(_03004_),
    .A2(_02676_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27033_ (.A1(_03005_),
    .A2(_02469_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27034_ (.A1(_02604_),
    .A2(_15995_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27035_ (.A1(_03007_),
    .A2(_02589_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27036_ (.A1(_03008_),
    .A2(_02689_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27037_ (.A1(_02784_),
    .A2(_02568_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27038_ (.A1(_03009_),
    .A2(_03010_),
    .B(_02497_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27039_ (.A1(_03006_),
    .A2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27040_ (.A1(_03003_),
    .A2(_03012_),
    .B(_02504_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27041_ (.A1(_02999_),
    .A2(_03013_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27042_ (.A1(_02986_),
    .A2(_03014_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _27043_ (.I(\sa31_sub[7] ),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27044_ (.A1(_03015_),
    .A2(\sa31_sub[0] ),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27045_ (.A1(_12002_),
    .A2(_12251_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27046_ (.A1(_03017_),
    .A2(_03016_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27047_ (.A1(_03018_),
    .A2(net1168),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27048_ (.A1(_12002_),
    .A2(_03015_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27049_ (.A1(net789),
    .A2(_12251_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27050_ (.A1(_03021_),
    .A2(_03020_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27051_ (.A1(_03022_),
    .A2(\sa31_sub[1] ),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27052_ (.A1(_03023_),
    .A2(_03019_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27053_ (.I(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27054_ (.A1(\sa12_sr[1] ),
    .A2(\sa02_sr[1] ),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27055_ (.A1(net1192),
    .A2(_15064_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27056_ (.A1(_12024_),
    .A2(_15062_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27057_ (.A1(_03027_),
    .A2(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27058_ (.A1(_03025_),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27059_ (.A1(_15064_),
    .A2(_12024_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27060_ (.A1(net1192),
    .A2(_15062_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27061_ (.A1(_03031_),
    .A2(_03032_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27062_ (.A1(_03024_),
    .A2(_03033_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27063_ (.A1(_03034_),
    .A2(_03030_),
    .B(_10526_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27064_ (.I(\text_in_r[41] ),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27065_ (.A1(_03036_),
    .A2(_10586_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27066_ (.A1(_03037_),
    .A2(_03035_),
    .B(\u0.w[2][9] ),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27067_ (.A1(_03034_),
    .A2(_03030_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27068_ (.A1(_03039_),
    .A2(_11348_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27069_ (.I(\u0.w[2][9] ),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27070_ (.I(_03037_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27071_ (.A1(_03040_),
    .A2(_03041_),
    .A3(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27072_ (.A1(_03038_),
    .A2(_03043_),
    .ZN(_16007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27073_ (.A1(net1177),
    .A2(net1180),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27074_ (.A1(net1177),
    .A2(\sa12_sr[0] ),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27075_ (.A1(_03044_),
    .A2(_03045_),
    .B(_15059_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27076_ (.I(_03045_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27077_ (.A1(net1177),
    .A2(net1178),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27078_ (.A1(_03047_),
    .A2(_12250_),
    .A3(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27079_ (.A1(_03046_),
    .A2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27080_ (.A1(_03050_),
    .A2(_03022_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27081_ (.A1(_03046_),
    .A2(_03049_),
    .A3(_03018_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27082_ (.A1(_03051_),
    .A2(_03052_),
    .B(_10525_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27083_ (.I(\text_in_r[40] ),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27084_ (.A1(_03054_),
    .A2(_10381_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27085_ (.A1(_03053_),
    .A2(_03055_),
    .B(\u0.w[2][8] ),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27086_ (.A1(_03051_),
    .A2(_03052_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27087_ (.A1(_03057_),
    .A2(_10405_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27088_ (.I(\u0.w[2][8] ),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27089_ (.I(_03055_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27090_ (.A1(_03058_),
    .A2(_03059_),
    .A3(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27091_ (.A1(_03056_),
    .A2(_03061_),
    .ZN(_16012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27092_ (.A1(_12031_),
    .A2(_12033_),
    .A3(\sa02_sr[2] ),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27093_ (.A1(_12032_),
    .A2(_12030_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27094_ (.A1(\sa12_sr[2] ),
    .A2(\sa31_sub[2] ),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27095_ (.A1(_03063_),
    .A2(_12057_),
    .A3(_03064_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27096_ (.A1(_03062_),
    .A2(_03065_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27097_ (.A1(_03066_),
    .A2(_11964_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27098_ (.A1(_03062_),
    .A2(_03065_),
    .A3(net1175),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27099_ (.A1(_03067_),
    .A2(_03068_),
    .B(_10410_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27100_ (.I(\text_in_r[42] ),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27101_ (.A1(_03070_),
    .A2(_11202_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27102_ (.I(\u0.w[2][10] ),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27103_ (.A1(_03069_),
    .A2(_03071_),
    .B(_03072_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27104_ (.A1(_03067_),
    .A2(_03068_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27105_ (.A1(_03074_),
    .A2(_10522_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27106_ (.I(_03071_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27107_ (.A1(_03075_),
    .A2(\u0.w[2][10] ),
    .A3(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27108_ (.A1(_03073_),
    .A2(_03077_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27109_ (.I(_03078_),
    .Z(_16028_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27110_ (.A1(_03037_),
    .A2(_03035_),
    .B(_03041_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27111_ (.A1(_03042_),
    .A2(\u0.w[2][9] ),
    .A3(_03040_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27112_ (.A1(_03079_),
    .A2(_03080_),
    .ZN(_16002_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27113_ (.A1(_03069_),
    .A2(_03071_),
    .B(\u0.w[2][10] ),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27114_ (.A1(_03075_),
    .A2(_03072_),
    .A3(_03076_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27115_ (.A1(_03081_),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _27116_ (.I(_03083_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _27117_ (.I(_03084_),
    .Z(_16021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27118_ (.I(_16003_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27119_ (.A1(_03084_),
    .A2(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27120_ (.A1(net643),
    .A2(\sa31_sub[2] ),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27121_ (.A1(net701),
    .A2(_15131_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27122_ (.A1(_12030_),
    .A2(_03015_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27123_ (.A1(\sa31_sub[2] ),
    .A2(_12251_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27124_ (.A1(_03089_),
    .A2(_03090_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27125_ (.A1(_15135_),
    .A2(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27126_ (.A1(_03092_),
    .A2(_03088_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27127_ (.A1(\sa12_sr[3] ),
    .A2(\sa02_sr[3] ),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27128_ (.A1(_03094_),
    .A2(_12066_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27129_ (.A1(\sa12_sr[3] ),
    .A2(\sa02_sr[3] ),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27130_ (.A1(\sa12_sr[3] ),
    .A2(\sa02_sr[3] ),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27131_ (.A1(_03096_),
    .A2(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27132_ (.A1(_03098_),
    .A2(\sa31_sub[3] ),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27133_ (.A1(_03095_),
    .A2(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27134_ (.A1(_03093_),
    .A2(_03100_),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27135_ (.A1(_03093_),
    .A2(_03100_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27136_ (.A1(_03101_),
    .A2(_10549_),
    .A3(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27137_ (.A1(_12193_),
    .A2(\text_in_r[43] ),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27138_ (.A1(_03104_),
    .A2(\u0.w[2][11] ),
    .A3(_03103_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27139_ (.A1(_03087_),
    .A2(_03098_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27140_ (.A1(_03094_),
    .A2(_03091_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27141_ (.A1(_03107_),
    .A2(_03106_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27142_ (.A1(_15135_),
    .A2(\sa31_sub[3] ),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27143_ (.A1(_15131_),
    .A2(_12066_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27144_ (.A1(_03109_),
    .A2(_03110_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27145_ (.I(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27146_ (.A1(_03108_),
    .A2(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27147_ (.A1(_03094_),
    .A2(_03091_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27148_ (.A1(_03087_),
    .A2(_03098_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27149_ (.A1(_03114_),
    .A2(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27150_ (.A1(_03116_),
    .A2(_03111_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27151_ (.A1(_03117_),
    .A2(_03113_),
    .A3(_10405_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27152_ (.I(\u0.w[2][11] ),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27153_ (.A1(_10522_),
    .A2(\text_in_r[43] ),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27154_ (.A1(_03118_),
    .A2(_03119_),
    .A3(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27155_ (.A1(_03121_),
    .A2(_03105_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27156_ (.I(_03122_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27157_ (.A1(_03086_),
    .A2(_03123_),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _27158_ (.A1(\sa12_sr[4] ),
    .A2(\sa02_sr[4] ),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27159_ (.A1(\sa31_sub[3] ),
    .A2(net642),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27160_ (.A1(_03125_),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _27161_ (.A1(\sa31_sub[3] ),
    .A2(_12251_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27162_ (.A1(_03128_),
    .A2(_12148_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27163_ (.A1(_03127_),
    .A2(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27164_ (.I(\sa31_sub[4] ),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27165_ (.A1(_03131_),
    .A2(_15156_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27166_ (.A1(_03132_),
    .A2(_03130_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27167_ (.A1(\sa31_sub[4] ),
    .A2(_15156_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27168_ (.A1(_03127_),
    .A2(_03129_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27169_ (.A1(_03134_),
    .A2(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27170_ (.A1(_13010_),
    .A2(_03136_),
    .A3(_03133_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27171_ (.A1(_10526_),
    .A2(\text_in_r[44] ),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27172_ (.A1(_03138_),
    .A2(_03137_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27173_ (.A1(_03139_),
    .A2(\u0.w[2][12] ),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27174_ (.I(\u0.w[2][12] ),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27175_ (.A1(_03137_),
    .A2(_03141_),
    .A3(_03138_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27176_ (.A1(_03140_),
    .A2(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _27177_ (.I(_03143_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27178_ (.A1(_03124_),
    .A2(_03144_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27179_ (.I(_03078_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27180_ (.I(_16013_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27181_ (.A1(_03146_),
    .A2(_03147_),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27182_ (.A1(_03103_),
    .A2(_03119_),
    .A3(_03104_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27183_ (.A1(_03120_),
    .A2(\u0.w[2][11] ),
    .A3(_03118_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27184_ (.A1(_03149_),
    .A2(_03150_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27185_ (.I(_03151_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 _27186_ (.I(_03152_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27187_ (.A1(_03148_),
    .A2(net704),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _27188_ (.I(_16004_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27189_ (.A1(_03155_),
    .A2(_03083_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27190_ (.A1(net647),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _27191_ (.I(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27192_ (.A1(_16028_),
    .A2(_16003_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27193_ (.A1(_03158_),
    .A2(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27194_ (.A1(_03145_),
    .A2(_03154_),
    .A3(_03160_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27195_ (.A1(_03146_),
    .A2(net15),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27196_ (.I(_03162_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27197_ (.I(_03152_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27198_ (.A1(_03163_),
    .A2(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27199_ (.I(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27200_ (.I(_03156_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27201_ (.A1(_03167_),
    .A2(net703),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27202_ (.A1(_03078_),
    .A2(_03155_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27203_ (.A1(net647),
    .A2(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27204_ (.A1(_03168_),
    .A2(_03170_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27205_ (.A1(_03139_),
    .A2(_03141_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27206_ (.A1(_03137_),
    .A2(\u0.w[2][12] ),
    .A3(_03138_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27207_ (.A1(_03173_),
    .A2(_03172_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27208_ (.I(_03174_),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27209_ (.I(_03175_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27210_ (.A1(_03166_),
    .A2(_03171_),
    .B(_03176_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27211_ (.A1(\sa31_sub[5] ),
    .A2(_15154_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27212_ (.I(_12187_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27213_ (.A1(_03178_),
    .A2(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27214_ (.I(\sa31_sub[5] ),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27215_ (.A1(_03181_),
    .A2(_15154_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27216_ (.A1(_03182_),
    .A2(_12187_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27217_ (.A1(_03180_),
    .A2(_03183_),
    .A3(_10549_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27218_ (.A1(_10483_),
    .A2(\text_in_r[45] ),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27219_ (.A1(_03184_),
    .A2(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27220_ (.A1(_03186_),
    .A2(\u0.w[2][13] ),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27221_ (.A1(_03186_),
    .A2(\u0.w[2][13] ),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27222_ (.A1(_03187_),
    .A2(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _27223_ (.I(_03189_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27224_ (.A1(_03161_),
    .A2(_03177_),
    .A3(_03190_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _27225_ (.I(_16012_),
    .ZN(_16001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27226_ (.A1(net15),
    .A2(net639),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27227_ (.A1(net29),
    .A2(_03084_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27228_ (.A1(_03192_),
    .A2(_03193_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 _27229_ (.I(_03123_),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27230_ (.A1(_03194_),
    .A2(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27231_ (.A1(_03193_),
    .A2(_03152_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27232_ (.I(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27233_ (.A1(_03198_),
    .A2(_03192_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27234_ (.A1(_03196_),
    .A2(_03199_),
    .A3(_03176_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27235_ (.A1(_03146_),
    .A2(_16017_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27236_ (.I(_03151_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27237_ (.A1(_03201_),
    .A2(_03202_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27238_ (.A1(_03203_),
    .A2(net44),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27239_ (.I(_03144_),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27240_ (.A1(_16021_),
    .A2(_16013_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27241_ (.I(_03123_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27242_ (.A1(_03159_),
    .A2(_03206_),
    .A3(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27243_ (.A1(_03204_),
    .A2(_03205_),
    .A3(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27244_ (.I(_03189_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27245_ (.I(_03210_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _27246_ (.I(_03211_),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27247_ (.A1(_03200_),
    .A2(_03209_),
    .A3(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27248_ (.A1(\sa12_sr[6] ),
    .A2(\sa31_sub[6] ),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27249_ (.A1(_15233_),
    .A2(_03214_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27250_ (.A1(_12151_),
    .A2(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _27251_ (.I0(_03216_),
    .I1(\text_in_r[46] ),
    .S(_12115_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27252_ (.A1(_03217_),
    .A2(\u0.w[2][14] ),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27253_ (.A1(_03217_),
    .A2(\u0.w[2][14] ),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27254_ (.A1(_03218_),
    .A2(_03219_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27255_ (.I(_03220_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27256_ (.A1(_03191_),
    .A2(_03213_),
    .A3(_03221_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27257_ (.A1(_03084_),
    .A2(_16005_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27258_ (.I(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27259_ (.A1(_03224_),
    .A2(_03202_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27260_ (.A1(_03225_),
    .A2(_03144_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27261_ (.A1(net638),
    .A2(_03146_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _27262_ (.I(_03122_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27263_ (.A1(_16017_),
    .A2(_03083_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27264_ (.A1(_03227_),
    .A2(_03228_),
    .A3(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27265_ (.A1(_03226_),
    .A2(_03165_),
    .A3(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27266_ (.A1(_03078_),
    .A2(_16008_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27267_ (.A1(_03232_),
    .A2(_03202_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27268_ (.I(_03233_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27269_ (.A1(net637),
    .A2(_03084_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27270_ (.I(_03235_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27271_ (.A1(_03234_),
    .A2(_03236_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27272_ (.I(_16019_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27273_ (.A1(_16021_),
    .A2(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27274_ (.A1(_03227_),
    .A2(_03207_),
    .A3(_03239_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27275_ (.A1(_03237_),
    .A2(_03240_),
    .A3(_03176_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27276_ (.A1(_03231_),
    .A2(_03241_),
    .A3(_03190_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27277_ (.A1(net638),
    .A2(_03084_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27278_ (.A1(_03234_),
    .A2(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27279_ (.A1(_03146_),
    .A2(_03238_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27280_ (.A1(_03158_),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27281_ (.I(_03174_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27282_ (.A1(_03244_),
    .A2(_03246_),
    .A3(_03247_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27283_ (.A1(_03232_),
    .A2(net647),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _27284_ (.I(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _27285_ (.I(_16010_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27286_ (.A1(_03084_),
    .A2(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27287_ (.A1(_03250_),
    .A2(net705),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27288_ (.A1(_03227_),
    .A2(_03202_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27289_ (.A1(_03253_),
    .A2(_03205_),
    .A3(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27290_ (.A1(_03248_),
    .A2(_03255_),
    .A3(_03212_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _27291_ (.I(_03220_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27292_ (.I(_03257_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27293_ (.A1(_03242_),
    .A2(_03256_),
    .A3(_03258_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _27294_ (.A1(net642),
    .A2(net1174),
    .A3(_12190_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27295_ (.A1(_12961_),
    .A2(\text_in_r[47] ),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27296_ (.A1(_03260_),
    .A2(_12965_),
    .B(_03261_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27297_ (.A1(\u0.w[2][15] ),
    .A2(_03262_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27298_ (.I(_03263_),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27299_ (.A1(_03222_),
    .A2(_03259_),
    .A3(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27300_ (.I(_16008_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27301_ (.A1(_03084_),
    .A2(_03266_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27302_ (.A1(_03267_),
    .A2(_03123_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27303_ (.A1(_03268_),
    .A2(_03154_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27304_ (.A1(_03224_),
    .A2(net703),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27305_ (.A1(_03270_),
    .A2(net644),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27306_ (.A1(_03269_),
    .A2(_03271_),
    .B(_03257_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27307_ (.A1(_16021_),
    .A2(_16008_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27308_ (.A1(_03273_),
    .A2(_03228_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27309_ (.I(_16015_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27310_ (.A1(_03275_),
    .A2(_03078_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27311_ (.A1(_03274_),
    .A2(net883),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27312_ (.I(_03144_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27313_ (.A1(_03277_),
    .A2(_03278_),
    .A3(_03225_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _27314_ (.I(_03189_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27315_ (.A1(_03272_),
    .A2(_03279_),
    .B(_03280_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27316_ (.A1(_03146_),
    .A2(_16013_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27317_ (.I(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27318_ (.A1(net29),
    .A2(_16028_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27319_ (.A1(_03283_),
    .A2(_03284_),
    .A3(_03164_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27320_ (.A1(net48),
    .A2(_03084_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27321_ (.A1(_03146_),
    .A2(_16004_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27322_ (.A1(_03286_),
    .A2(_03287_),
    .A3(net704),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27323_ (.I(_03174_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27324_ (.A1(_03285_),
    .A2(_03288_),
    .B(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27325_ (.A1(_16028_),
    .A2(_03085_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27326_ (.I(_03202_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27327_ (.A1(_03291_),
    .A2(_03224_),
    .B(_03292_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27328_ (.A1(_03252_),
    .A2(net703),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27329_ (.I(_03143_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27330_ (.A1(_03293_),
    .A2(_03294_),
    .B(_03295_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27331_ (.A1(_03290_),
    .A2(_03296_),
    .B(_03258_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27332_ (.A1(_03281_),
    .A2(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27333_ (.A1(_03287_),
    .A2(_03202_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27334_ (.A1(net704),
    .A2(_16026_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27335_ (.A1(_03299_),
    .A2(_03300_),
    .B(net645),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27336_ (.A1(_03301_),
    .A2(_03220_),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27337_ (.A1(_16021_),
    .A2(_16003_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27338_ (.A1(_03227_),
    .A2(_03228_),
    .A3(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27339_ (.A1(_16028_),
    .A2(_16005_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27340_ (.A1(_03305_),
    .A2(net703),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27341_ (.A1(_03304_),
    .A2(_03306_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27342_ (.A1(_03268_),
    .A2(_03144_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27343_ (.A1(_03078_),
    .A2(_16010_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27344_ (.I(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27345_ (.A1(_03310_),
    .A2(_03202_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27346_ (.I(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27347_ (.A1(_03308_),
    .A2(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27348_ (.A1(_03307_),
    .A2(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27349_ (.I(_03210_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27350_ (.A1(_03302_),
    .A2(_03314_),
    .B(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27351_ (.A1(_03230_),
    .A2(_03144_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27352_ (.A1(_03317_),
    .A2(_03311_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27353_ (.A1(_03084_),
    .A2(_16015_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27354_ (.A1(_03309_),
    .A2(_03319_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27355_ (.A1(_03320_),
    .A2(_03164_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27356_ (.A1(_03321_),
    .A2(_03247_),
    .A3(_03157_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27357_ (.A1(_03318_),
    .A2(_03258_),
    .A3(_03322_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27358_ (.A1(_03316_),
    .A2(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _27359_ (.I(_03263_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27360_ (.A1(_03298_),
    .A2(_03324_),
    .A3(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27361_ (.A1(_03265_),
    .A2(_03326_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _27362_ (.I(_03170_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27363_ (.A1(_03327_),
    .A2(_03239_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27364_ (.A1(_03313_),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27365_ (.A1(_03311_),
    .A2(net645),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27366_ (.A1(_03202_),
    .A2(_16033_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27367_ (.I(_03235_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 _27368_ (.I(_03153_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27369_ (.A1(_03332_),
    .A2(_03333_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27370_ (.A1(_03330_),
    .A2(_03331_),
    .A3(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27371_ (.A1(_03329_),
    .A2(_03335_),
    .A3(_03190_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27372_ (.A1(_03158_),
    .A2(_03227_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27373_ (.A1(_03252_),
    .A2(_03202_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27374_ (.I(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27375_ (.A1(net29),
    .A2(_03146_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27376_ (.A1(_03339_),
    .A2(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27377_ (.A1(_03337_),
    .A2(_03341_),
    .A3(_03176_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27378_ (.A1(_03286_),
    .A2(net702),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27379_ (.A1(_03343_),
    .A2(_03192_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27380_ (.A1(net648),
    .A2(_16028_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27381_ (.I(_03174_),
    .Z(_03346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27382_ (.A1(_03345_),
    .A2(_03266_),
    .B(net646),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27383_ (.A1(_03344_),
    .A2(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27384_ (.A1(_03342_),
    .A2(_03348_),
    .A3(_03212_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27385_ (.A1(_03336_),
    .A2(_03349_),
    .A3(_03221_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27386_ (.A1(net48),
    .A2(net29),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27387_ (.I(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27388_ (.I(_03228_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27389_ (.A1(_03352_),
    .A2(_03284_),
    .B(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27390_ (.A1(_03299_),
    .A2(_03243_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27391_ (.A1(_03354_),
    .A2(_03278_),
    .A3(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27392_ (.A1(_03340_),
    .A2(net702),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27393_ (.A1(_03357_),
    .A2(_03086_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27394_ (.A1(_03158_),
    .A2(_03309_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27395_ (.A1(_03358_),
    .A2(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27396_ (.I(_03175_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27397_ (.A1(_03360_),
    .A2(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27398_ (.A1(_03356_),
    .A2(_03362_),
    .A3(_03190_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27399_ (.A1(_16021_),
    .A2(_16010_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27400_ (.A1(_03364_),
    .A2(_03292_),
    .B(net645),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27401_ (.A1(_03201_),
    .A2(_03123_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27402_ (.A1(net634),
    .A2(_16021_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27403_ (.A1(_03366_),
    .A2(net881),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _27404_ (.I(_03189_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27405_ (.A1(_03365_),
    .A2(_03368_),
    .B(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27406_ (.A1(_03245_),
    .A2(net703),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27407_ (.A1(_03371_),
    .A2(_03236_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27408_ (.I(_16017_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27409_ (.A1(_16021_),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27410_ (.A1(_03374_),
    .A2(_03195_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27411_ (.A1(_03372_),
    .A2(_03247_),
    .A3(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27412_ (.A1(_03370_),
    .A2(_03376_),
    .B(_03220_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27413_ (.A1(_03363_),
    .A2(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27414_ (.A1(_03350_),
    .A2(_03325_),
    .A3(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27415_ (.I(_03254_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27416_ (.A1(_03380_),
    .A2(_03229_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27417_ (.A1(_03157_),
    .A2(_03144_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27418_ (.A1(_03381_),
    .A2(_03382_),
    .B(_03211_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27419_ (.I(_16005_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27420_ (.A1(_03146_),
    .A2(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27421_ (.A1(_03385_),
    .A2(_03152_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27422_ (.A1(_03386_),
    .A2(_03239_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27423_ (.A1(_03368_),
    .A2(_03387_),
    .A3(_03176_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27424_ (.A1(_03383_),
    .A2(_03388_),
    .B(_03220_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27425_ (.A1(_03327_),
    .A2(_03303_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27426_ (.A1(_03390_),
    .A2(_03225_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27427_ (.A1(_03195_),
    .A2(_03340_),
    .B(net644),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27428_ (.A1(_03391_),
    .A2(_03392_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _27429_ (.A1(_03163_),
    .A2(_03294_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27430_ (.I(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27431_ (.A1(_03198_),
    .A2(_03159_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27432_ (.A1(_03395_),
    .A2(_03396_),
    .A3(_03205_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27433_ (.A1(_03393_),
    .A2(_03212_),
    .A3(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27434_ (.A1(_03398_),
    .A2(_03389_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27435_ (.A1(_03243_),
    .A2(_03153_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27436_ (.A1(_03400_),
    .A2(_03159_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27437_ (.A1(_03250_),
    .A2(_03229_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27438_ (.A1(_03401_),
    .A2(_03211_),
    .A3(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27439_ (.A1(_03403_),
    .A2(_03361_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27440_ (.A1(net48),
    .A2(_16028_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27441_ (.A1(_03198_),
    .A2(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27442_ (.A1(_03395_),
    .A2(_03369_),
    .A3(_03406_),
    .Z(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27443_ (.I(_16029_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27444_ (.A1(_03189_),
    .A2(_03408_),
    .A3(_03207_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27445_ (.A1(_03229_),
    .A2(_03152_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27446_ (.A1(_03410_),
    .A2(_03282_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27447_ (.A1(_03409_),
    .A2(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27448_ (.A1(_03412_),
    .A2(_03278_),
    .B(_03257_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27449_ (.A1(_03404_),
    .A2(_03407_),
    .B(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27450_ (.A1(_03399_),
    .A2(_03414_),
    .A3(_03264_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27451_ (.A1(_03379_),
    .A2(_03415_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27452_ (.A1(_16028_),
    .A2(_03251_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27453_ (.A1(_03158_),
    .A2(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27454_ (.A1(_03417_),
    .A2(_03145_),
    .B(_03369_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27455_ (.A1(_03384_),
    .A2(_03251_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27456_ (.A1(_03419_),
    .A2(_16021_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27457_ (.A1(_03366_),
    .A2(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27458_ (.A1(_03411_),
    .A2(_03421_),
    .A3(_03176_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27459_ (.A1(_03422_),
    .A2(_03418_),
    .B(_03257_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27460_ (.I(_03286_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _27461_ (.A1(_03424_),
    .A2(_03249_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27462_ (.A1(_03333_),
    .A2(_16035_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27463_ (.A1(_03247_),
    .A2(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27464_ (.I(_16024_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27465_ (.A1(_03228_),
    .A2(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27466_ (.A1(_03233_),
    .A2(_03429_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _27467_ (.A1(_03425_),
    .A2(_03427_),
    .B1(_03430_),
    .B2(_03361_),
    .C(_03280_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27468_ (.A1(_03423_),
    .A2(_03431_),
    .B(_03264_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27469_ (.A1(_03286_),
    .A2(_03192_),
    .A3(_03195_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _27470_ (.A1(_16029_),
    .A2(_03353_),
    .B(_03433_),
    .C(_03205_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27471_ (.A1(_03424_),
    .A2(_03207_),
    .A3(_03291_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27472_ (.A1(_16021_),
    .A2(_03147_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27473_ (.A1(_03287_),
    .A2(_03436_),
    .A3(_03195_),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27474_ (.A1(_03435_),
    .A2(_03437_),
    .B(_03361_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27475_ (.A1(_03434_),
    .A2(_03190_),
    .A3(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27476_ (.A1(net877),
    .A2(_03228_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27477_ (.A1(_03440_),
    .A2(_03243_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27478_ (.A1(_03441_),
    .A2(_03361_),
    .A3(_03288_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27479_ (.A1(_16026_),
    .A2(_03333_),
    .B(net646),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27480_ (.A1(_03274_),
    .A2(net879),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27481_ (.A1(_03443_),
    .A2(_03444_),
    .B(_03369_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27482_ (.A1(_03442_),
    .A2(_03445_),
    .B(_03221_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27483_ (.A1(_03446_),
    .A2(_03439_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27484_ (.A1(_03447_),
    .A2(_03432_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27485_ (.I(_03245_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _27486_ (.A1(_03449_),
    .A2(_03338_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27487_ (.A1(_03425_),
    .A2(_03450_),
    .B(net646),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27488_ (.I(_03143_),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27489_ (.I(_03122_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27490_ (.A1(_03309_),
    .A2(_03267_),
    .A3(_03453_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27491_ (.A1(_03288_),
    .A2(_03452_),
    .A3(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27492_ (.A1(_03451_),
    .A2(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27493_ (.A1(_03456_),
    .A2(_03190_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27494_ (.A1(_03405_),
    .A2(_03167_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27495_ (.A1(_03193_),
    .A2(_03305_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27496_ (.A1(_03459_),
    .A2(_03207_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _27497_ (.A1(_03353_),
    .A2(_03458_),
    .B(_03460_),
    .C(_03289_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27498_ (.A1(_03366_),
    .A2(_03239_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27499_ (.A1(_03233_),
    .A2(_03144_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27500_ (.A1(_03462_),
    .A2(_03463_),
    .B(_03369_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27501_ (.A1(_03461_),
    .A2(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27502_ (.A1(_03457_),
    .A2(_03465_),
    .A3(_03221_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27503_ (.A1(net877),
    .A2(_03195_),
    .A3(_03319_),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27504_ (.A1(_03146_),
    .A2(_16019_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27505_ (.I(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27506_ (.A1(_03197_),
    .A2(_03469_),
    .B(_03174_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27507_ (.A1(_03467_),
    .A2(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27508_ (.A1(_03243_),
    .A2(net704),
    .A3(net883),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27509_ (.A1(net44),
    .A2(_03287_),
    .A3(_03207_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27510_ (.A1(_03473_),
    .A2(_03472_),
    .B(_03289_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27511_ (.A1(_03471_),
    .A2(_03474_),
    .B(_03315_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27512_ (.A1(_03416_),
    .A2(_03228_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27513_ (.A1(_03476_),
    .A2(_03236_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27514_ (.A1(_03477_),
    .A2(_03295_),
    .A3(_03321_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27515_ (.A1(_03309_),
    .A2(_03195_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27516_ (.I(_03193_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27517_ (.A1(_03468_),
    .A2(_03153_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27518_ (.A1(_03479_),
    .A2(_03480_),
    .B(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27519_ (.I(_03319_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27520_ (.A1(_03483_),
    .A2(_03292_),
    .B(_03452_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27521_ (.A1(_03482_),
    .A2(_03484_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27522_ (.A1(_03478_),
    .A2(_03485_),
    .A3(_03280_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27523_ (.A1(_03475_),
    .A2(_03258_),
    .A3(_03486_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27524_ (.A1(_03466_),
    .A2(_03487_),
    .A3(_03264_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27525_ (.A1(_03488_),
    .A2(_03448_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27526_ (.A1(_03410_),
    .A2(net880),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27527_ (.A1(_03250_),
    .A2(_03206_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27528_ (.A1(_03489_),
    .A2(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27529_ (.A1(_03491_),
    .A2(_03295_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27530_ (.A1(_03167_),
    .A2(net702),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27531_ (.A1(_03493_),
    .A2(_03148_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27532_ (.A1(_03196_),
    .A2(_03494_),
    .A3(_03289_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27533_ (.A1(_03492_),
    .A2(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27534_ (.A1(_03496_),
    .A2(_03212_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27535_ (.A1(_03192_),
    .A2(_03340_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27536_ (.A1(_03498_),
    .A2(_03333_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27537_ (.A1(_03499_),
    .A2(_03278_),
    .A3(_03249_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27538_ (.A1(_03276_),
    .A2(net702),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27539_ (.A1(_03501_),
    .A2(net882),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27540_ (.A1(_03372_),
    .A2(_03502_),
    .A3(_03247_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27541_ (.A1(_03500_),
    .A2(_03503_),
    .A3(_03190_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27542_ (.A1(_03497_),
    .A2(_03504_),
    .A3(_03258_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27543_ (.A1(net877),
    .A2(_03353_),
    .A3(net44),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27544_ (.A1(_03499_),
    .A2(_03506_),
    .A3(_03278_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27545_ (.A1(net877),
    .A2(_03243_),
    .A3(_03333_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27546_ (.A1(_03508_),
    .A2(_03176_),
    .A3(_03170_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27547_ (.A1(_03507_),
    .A2(_03509_),
    .A3(_03280_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27548_ (.A1(_03458_),
    .A2(_03333_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27549_ (.A1(_03476_),
    .A2(_03239_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27550_ (.A1(_03511_),
    .A2(_03512_),
    .A3(_03205_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27551_ (.A1(_03340_),
    .A2(_03436_),
    .A3(_03164_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27552_ (.A1(_03086_),
    .A2(net880),
    .A3(_03195_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27553_ (.A1(_03514_),
    .A2(_03515_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27554_ (.A1(_03516_),
    .A2(_03176_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27555_ (.A1(_03513_),
    .A2(_03212_),
    .A3(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27556_ (.A1(_03510_),
    .A2(_03518_),
    .A3(_03221_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27557_ (.A1(_03505_),
    .A2(_03519_),
    .A3(_03325_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27558_ (.I(_03344_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27559_ (.A1(_03304_),
    .A2(_03452_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27560_ (.A1(_03521_),
    .A2(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27561_ (.A1(_03227_),
    .A2(_03319_),
    .B(_03153_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27562_ (.A1(_03493_),
    .A2(_03449_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27563_ (.A1(_03524_),
    .A2(_03452_),
    .A3(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27564_ (.A1(_03523_),
    .A2(_03526_),
    .B(_03315_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27565_ (.A1(_03276_),
    .A2(net648),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27566_ (.I(_03528_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27567_ (.A1(_03529_),
    .A2(_03420_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27568_ (.A1(_03411_),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27569_ (.A1(_03531_),
    .A2(_03295_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27570_ (.A1(_03470_),
    .A2(_03189_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27571_ (.A1(_03532_),
    .A2(_03533_),
    .B(_03220_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27572_ (.A1(_03527_),
    .A2(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27573_ (.A1(_03282_),
    .A2(_03202_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27574_ (.A1(_03211_),
    .A2(_03424_),
    .A3(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _27575_ (.A1(_03189_),
    .A2(_03168_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27576_ (.A1(_03537_),
    .A2(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27577_ (.A1(_03210_),
    .A2(_03164_),
    .A3(net880),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27578_ (.I(_03271_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27579_ (.A1(_03540_),
    .A2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27580_ (.A1(_03539_),
    .A2(_03542_),
    .B(_03257_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27581_ (.A1(_03371_),
    .A2(_03420_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27582_ (.A1(_03227_),
    .A2(net704),
    .A3(_03167_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27583_ (.A1(_03545_),
    .A2(_03544_),
    .A3(_03189_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27584_ (.A1(_03483_),
    .A2(_03453_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27585_ (.A1(_03472_),
    .A2(_03211_),
    .A3(_03547_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27586_ (.A1(_03546_),
    .A2(_03548_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27587_ (.A1(_03549_),
    .A2(_03278_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27588_ (.A1(_03543_),
    .A2(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27589_ (.A1(_03535_),
    .A2(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27590_ (.A1(_03552_),
    .A2(_03264_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27591_ (.A1(_03520_),
    .A2(_03553_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27592_ (.A1(_03405_),
    .A2(_03243_),
    .A3(_03453_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27593_ (.A1(_03401_),
    .A2(_03554_),
    .A3(_03278_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27594_ (.A1(_03529_),
    .A2(_03452_),
    .A3(_03224_),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27595_ (.A1(_03555_),
    .A2(_03212_),
    .A3(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27596_ (.A1(_03433_),
    .A2(_03406_),
    .A3(_03278_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27597_ (.A1(_03236_),
    .A2(_03351_),
    .A3(_03333_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27598_ (.A1(_03236_),
    .A2(_03207_),
    .A3(_03159_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27599_ (.A1(_03559_),
    .A2(_03560_),
    .A3(_03247_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27600_ (.A1(_03558_),
    .A2(_03561_),
    .A3(_03190_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27601_ (.A1(_03557_),
    .A2(_03562_),
    .A3(_03258_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27602_ (.A1(_03440_),
    .A2(_03303_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27603_ (.A1(_03313_),
    .A2(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27604_ (.I(_03450_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27605_ (.A1(_03274_),
    .A2(net878),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27606_ (.A1(_03566_),
    .A2(_03567_),
    .A3(_03247_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27607_ (.A1(_03565_),
    .A2(_03568_),
    .A3(_03280_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27608_ (.A1(_03483_),
    .A2(_03207_),
    .B(_03144_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27609_ (.I(_03287_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27610_ (.A1(_03571_),
    .A2(_03228_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27611_ (.I(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27612_ (.A1(_03570_),
    .A2(_03573_),
    .A3(_03321_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27613_ (.A1(net879),
    .A2(_03239_),
    .A3(_03292_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27614_ (.A1(_03277_),
    .A2(_03205_),
    .A3(_03575_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27615_ (.A1(_03574_),
    .A2(_03576_),
    .A3(_03315_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27616_ (.A1(_03569_),
    .A2(_03577_),
    .A3(_03221_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27617_ (.A1(_03563_),
    .A2(_03578_),
    .A3(_03325_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27618_ (.A1(_03235_),
    .A2(_03351_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27619_ (.A1(_03580_),
    .A2(_03292_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27620_ (.A1(_03529_),
    .A2(_03193_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27621_ (.A1(_03581_),
    .A2(_03582_),
    .B(_03295_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27622_ (.A1(_03196_),
    .A2(_03293_),
    .B(_03289_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27623_ (.A1(_03583_),
    .A2(_03584_),
    .B(_03221_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27624_ (.A1(_03162_),
    .A2(_03086_),
    .B(_03195_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27625_ (.A1(_03586_),
    .A2(_03394_),
    .B(net646),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27626_ (.I(_03345_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27627_ (.A1(_03197_),
    .A2(_03449_),
    .B(_03588_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27628_ (.A1(_03589_),
    .A2(_03295_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27629_ (.A1(_03587_),
    .A2(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27630_ (.A1(_03591_),
    .A2(_03258_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27631_ (.A1(_03585_),
    .A2(_03592_),
    .A3(_03190_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27632_ (.A1(_03287_),
    .A2(_03453_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27633_ (.A1(_03153_),
    .A2(_03373_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27634_ (.A1(_03594_),
    .A2(_03144_),
    .A3(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27635_ (.A1(_03596_),
    .A2(_03257_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27636_ (.A1(_03268_),
    .A2(_03175_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27637_ (.A1(_03529_),
    .A2(_03236_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27638_ (.A1(_03598_),
    .A2(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27639_ (.A1(_03597_),
    .A2(_03600_),
    .B(_03280_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27640_ (.A1(_03339_),
    .A2(_03287_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27641_ (.A1(_03317_),
    .A2(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27642_ (.A1(_03366_),
    .A2(_03386_),
    .A3(_03452_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27643_ (.A1(_03603_),
    .A2(_03257_),
    .A3(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27644_ (.A1(_03601_),
    .A2(_03605_),
    .B(_03325_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27645_ (.A1(_03593_),
    .A2(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27646_ (.A1(_03579_),
    .A2(_03607_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27647_ (.A1(_03374_),
    .A2(_03453_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _27648_ (.A1(_03254_),
    .A2(_03352_),
    .B1(_03608_),
    .B2(_03148_),
    .C(_03346_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27649_ (.A1(net15),
    .A2(_03195_),
    .B(_03175_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27650_ (.A1(_03610_),
    .A2(_03581_),
    .B(_03369_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27651_ (.A1(_03609_),
    .A2(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27652_ (.A1(_03386_),
    .A2(_03286_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27653_ (.A1(_03613_),
    .A2(_03572_),
    .B(_03289_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _27654_ (.A1(_03157_),
    .A2(_03291_),
    .B(_03481_),
    .C(_03452_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27655_ (.A1(_03614_),
    .A2(_03369_),
    .A3(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27656_ (.A1(_03616_),
    .A2(_03612_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27657_ (.A1(_03617_),
    .A2(_03221_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27658_ (.A1(_16028_),
    .A2(_03266_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27659_ (.A1(_03338_),
    .A2(net645),
    .A3(_03619_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27660_ (.A1(_03620_),
    .A2(_03315_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27661_ (.A1(_03493_),
    .A2(_03452_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27662_ (.A1(_03524_),
    .A2(_03622_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27663_ (.A1(_03621_),
    .A2(_03623_),
    .B(_03220_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27664_ (.A1(_03371_),
    .A2(net705),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27665_ (.A1(_03226_),
    .A2(_03625_),
    .A3(_03165_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27666_ (.A1(_03501_),
    .A2(_03273_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27667_ (.I(_03419_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27668_ (.A1(_03476_),
    .A2(_03628_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27669_ (.A1(_03627_),
    .A2(_03629_),
    .A3(_03247_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27670_ (.A1(_03626_),
    .A2(_03630_),
    .A3(_03212_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27671_ (.A1(_03631_),
    .A2(_03624_),
    .B(_03264_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27672_ (.A1(_03632_),
    .A2(_03618_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27673_ (.A1(_03167_),
    .A2(_03468_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _27674_ (.A1(_03158_),
    .A2(_03282_),
    .B1(_03634_),
    .B2(_03333_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27675_ (.A1(_03635_),
    .A2(_03361_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27676_ (.A1(_03228_),
    .A2(_03147_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _27677_ (.A1(_03410_),
    .A2(net646),
    .A3(_03637_),
    .B(_03189_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27678_ (.I(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27679_ (.A1(_03636_),
    .A2(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27680_ (.A1(_03234_),
    .A2(_03229_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27681_ (.A1(_03420_),
    .A2(_03353_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27682_ (.A1(_03641_),
    .A2(_03205_),
    .A3(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27683_ (.I(_03371_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27684_ (.A1(_03330_),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27685_ (.A1(_03643_),
    .A2(_03645_),
    .A3(_03315_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27686_ (.A1(_03640_),
    .A2(_03221_),
    .A3(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27687_ (.A1(_03400_),
    .A2(_03416_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27688_ (.A1(_03317_),
    .A2(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27689_ (.A1(_03148_),
    .A2(_03207_),
    .B(_03452_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27690_ (.A1(_03410_),
    .A2(_03245_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27691_ (.A1(_03650_),
    .A2(_03651_),
    .B(_03211_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27692_ (.A1(_03649_),
    .A2(_03652_),
    .B(_03220_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27693_ (.A1(_03501_),
    .A2(_03235_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27694_ (.A1(_03250_),
    .A2(net44),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27695_ (.A1(_03654_),
    .A2(_03655_),
    .A3(_03176_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27696_ (.A1(_03353_),
    .A2(net29),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27697_ (.A1(_03199_),
    .A2(_03205_),
    .A3(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27698_ (.A1(_03656_),
    .A2(_03658_),
    .A3(_03212_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27699_ (.A1(_03653_),
    .A2(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27700_ (.A1(_03647_),
    .A2(_03660_),
    .A3(_03264_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27701_ (.A1(_03661_),
    .A2(_03633_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27702_ (.A1(_03405_),
    .A2(_03353_),
    .A3(_03273_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27703_ (.A1(_03662_),
    .A2(_03361_),
    .A3(_03154_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27704_ (.A1(_03274_),
    .A2(_03340_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27705_ (.A1(_03287_),
    .A2(_03420_),
    .A3(_03292_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27706_ (.A1(_03664_),
    .A2(_03205_),
    .A3(_03665_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27707_ (.A1(_03663_),
    .A2(_03666_),
    .A3(_03280_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27708_ (.A1(_03250_),
    .A2(_03236_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27709_ (.A1(net881),
    .A2(_03385_),
    .A3(_03292_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27710_ (.A1(_03668_),
    .A2(_03205_),
    .A3(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27711_ (.A1(_03430_),
    .A2(_03168_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27712_ (.A1(_03671_),
    .A2(_03361_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27713_ (.A1(_03670_),
    .A2(_03672_),
    .A3(_03315_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27714_ (.A1(_03667_),
    .A2(_03673_),
    .A3(_03221_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27715_ (.A1(_03193_),
    .A2(_03287_),
    .A3(_03292_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27716_ (.A1(_03345_),
    .A2(_03628_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27717_ (.A1(_03570_),
    .A2(_03675_),
    .A3(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27718_ (.A1(_16028_),
    .A2(_03373_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27719_ (.A1(_03223_),
    .A2(_03678_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27720_ (.A1(_03679_),
    .A2(_03353_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27721_ (.A1(net883),
    .A2(_03239_),
    .A3(_03164_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27722_ (.A1(_03680_),
    .A2(_03681_),
    .A3(_03295_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27723_ (.A1(_03677_),
    .A2(_03280_),
    .A3(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27724_ (.A1(_03580_),
    .A2(_03353_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27725_ (.A1(_16022_),
    .A2(_16031_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27726_ (.A1(_03333_),
    .A2(_03685_),
    .B(_03346_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27727_ (.A1(_03684_),
    .A2(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27728_ (.A1(_03319_),
    .A2(_03305_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27729_ (.A1(_03688_),
    .A2(_03353_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27730_ (.A1(_03689_),
    .A2(_03247_),
    .A3(_03124_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27731_ (.A1(_03687_),
    .A2(_03690_),
    .A3(_03315_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27732_ (.A1(_03683_),
    .A2(_03691_),
    .A3(_03258_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27733_ (.A1(_03674_),
    .A2(_03692_),
    .B(_03264_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27734_ (.A1(_03332_),
    .A2(_03528_),
    .B(_03536_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27735_ (.A1(_03694_),
    .A2(_03289_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27736_ (.A1(_03454_),
    .A2(_03295_),
    .B(_03211_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27737_ (.A1(_03695_),
    .A2(_03696_),
    .B(_03257_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27738_ (.A1(net702),
    .A2(_16023_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27739_ (.A1(_03698_),
    .A2(_03143_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27740_ (.A1(_03699_),
    .A2(_03654_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27741_ (.A1(_03634_),
    .A2(_03453_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27742_ (.A1(_03392_),
    .A2(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27743_ (.A1(_03700_),
    .A2(_03702_),
    .B(_03315_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27744_ (.A1(_03703_),
    .A2(_03697_),
    .B(_03325_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27745_ (.A1(_03357_),
    .A2(_03239_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27746_ (.A1(_03192_),
    .A2(_03453_),
    .A3(_03340_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27747_ (.A1(_03705_),
    .A2(_03706_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27748_ (.A1(_03707_),
    .A2(_03289_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27749_ (.A1(_03236_),
    .A2(_03164_),
    .A3(_03619_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27750_ (.A1(_03706_),
    .A2(_03709_),
    .A3(_03295_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27751_ (.A1(_03708_),
    .A2(_03710_),
    .A3(_03315_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27752_ (.A1(_03233_),
    .A2(_03284_),
    .B(_03331_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27753_ (.A1(_03712_),
    .A2(_03289_),
    .B(_03211_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27754_ (.I(_03367_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27755_ (.A1(_03714_),
    .A2(_03164_),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27756_ (.A1(_03524_),
    .A2(_03715_),
    .B(_03295_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27757_ (.A1(_03713_),
    .A2(_03716_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27758_ (.A1(_03711_),
    .A2(_03717_),
    .A3(_03258_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27759_ (.A1(_03718_),
    .A2(_03704_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27760_ (.A1(_03693_),
    .A2(_03719_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27761_ (.I(_03386_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27762_ (.A1(_03405_),
    .A2(_03453_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27763_ (.A1(_03720_),
    .A2(_03721_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27764_ (.A1(_03722_),
    .A2(_03189_),
    .A3(_03303_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27765_ (.A1(_03283_),
    .A2(_03714_),
    .A3(_03164_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27766_ (.A1(_03303_),
    .A2(_03201_),
    .A3(_03292_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27767_ (.A1(_03724_),
    .A2(_03725_),
    .B(_03369_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27768_ (.A1(_03723_),
    .A2(_03726_),
    .B(_03278_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27769_ (.A1(_16010_),
    .A2(_03333_),
    .B(_03211_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27770_ (.A1(_03728_),
    .A2(_03684_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27771_ (.A1(_03203_),
    .A2(_03286_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27772_ (.A1(_03730_),
    .A2(_03530_),
    .A3(_03211_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27773_ (.A1(_03729_),
    .A2(_03731_),
    .A3(_03361_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27774_ (.A1(_03727_),
    .A2(_03258_),
    .A3(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27775_ (.A1(_03598_),
    .A2(_03395_),
    .A3(_03165_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27776_ (.A1(_03373_),
    .A2(_03207_),
    .B(net645),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27777_ (.A1(_03735_),
    .A2(_03306_),
    .B(_03369_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27778_ (.A1(_03734_),
    .A2(_03736_),
    .B(_03257_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27779_ (.A1(_03380_),
    .A2(_03236_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27780_ (.A1(_03327_),
    .A2(net881),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27781_ (.A1(_03738_),
    .A2(_03361_),
    .A3(_03739_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27782_ (.A1(_03319_),
    .A2(_03169_),
    .B(_03453_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27783_ (.A1(_03228_),
    .A2(_16031_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27784_ (.A1(_03741_),
    .A2(_03346_),
    .A3(_03742_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27785_ (.A1(_03740_),
    .A2(_03743_),
    .A3(_03280_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27786_ (.A1(_03737_),
    .A2(_03744_),
    .B(_03264_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27787_ (.A1(_03733_),
    .A2(_03745_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27788_ (.A1(net44),
    .A2(_03678_),
    .B(_03453_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27789_ (.A1(_03747_),
    .A2(_03274_),
    .B(_03346_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27790_ (.A1(_03493_),
    .A2(_03608_),
    .A3(_03452_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27791_ (.A1(_03748_),
    .A2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27792_ (.A1(_03750_),
    .A2(_03190_),
    .B(_03257_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27793_ (.A1(net640),
    .A2(_03164_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27794_ (.A1(_03554_),
    .A2(_03346_),
    .A3(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27795_ (.A1(_03203_),
    .A2(_03236_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27796_ (.A1(_03433_),
    .A2(_03754_),
    .B(_03289_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27797_ (.A1(_03753_),
    .A2(_03755_),
    .B(_03212_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27798_ (.A1(_03751_),
    .A2(_03756_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27799_ (.A1(_03380_),
    .A2(_03273_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27800_ (.A1(_03366_),
    .A2(_03303_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27801_ (.A1(_03758_),
    .A2(_03176_),
    .A3(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27802_ (.A1(_03292_),
    .A2(_03239_),
    .B(_03175_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27803_ (.A1(_03761_),
    .A2(_03599_),
    .B(_03369_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27804_ (.A1(_03760_),
    .A2(_03762_),
    .B(_03220_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27805_ (.A1(_03441_),
    .A2(_03278_),
    .A3(_03681_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27806_ (.A1(_03328_),
    .A2(_03545_),
    .A3(_03247_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27807_ (.A1(_03764_),
    .A2(_03765_),
    .A3(_03280_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27808_ (.A1(_03766_),
    .A2(_03763_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27809_ (.A1(_03757_),
    .A2(_03767_),
    .A3(_03264_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27810_ (.A1(_03768_),
    .A2(_03746_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27811_ (.A1(\sa03_sr[1] ),
    .A2(net734),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27812_ (.A1(_03769_),
    .A2(_00811_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27813_ (.A1(_12833_),
    .A2(_00807_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27814_ (.A1(_03770_),
    .A2(_03771_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27815_ (.I(\sa32_sub[7] ),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27816_ (.A1(_12811_),
    .A2(_03773_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27817_ (.A1(\sa32_sub[0] ),
    .A2(_13067_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27818_ (.A1(_03774_),
    .A2(_03775_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27819_ (.A1(_03776_),
    .A2(_12766_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27820_ (.A1(_03773_),
    .A2(\sa32_sub[0] ),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27821_ (.A1(_12811_),
    .A2(_13067_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27822_ (.A1(_03778_),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27823_ (.A1(_03780_),
    .A2(net911),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27824_ (.A1(_03777_),
    .A2(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27825_ (.A1(_03782_),
    .A2(_03772_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27826_ (.A1(_03769_),
    .A2(_00807_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27827_ (.A1(_12833_),
    .A2(_00811_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27828_ (.A1(_03784_),
    .A2(_03785_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27829_ (.A1(_03780_),
    .A2(_12766_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27830_ (.A1(_03776_),
    .A2(\sa32_sub[1] ),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27831_ (.A1(_03787_),
    .A2(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27832_ (.A1(_03789_),
    .A2(_03786_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27833_ (.A1(net756),
    .A2(_03790_),
    .B(_12193_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27834_ (.I(\text_in_r[9] ),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27835_ (.A1(_03792_),
    .A2(_10410_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27836_ (.A1(_03791_),
    .A2(_03793_),
    .B(\u0.tmp_w[9] ),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27837_ (.A1(_03783_),
    .A2(_03790_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27838_ (.A1(_10403_),
    .A2(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27839_ (.I(\u0.tmp_w[9] ),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27840_ (.I(_03793_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27841_ (.A1(_03796_),
    .A2(_03797_),
    .A3(_03798_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27842_ (.A1(_03799_),
    .A2(_03794_),
    .ZN(_16043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27843_ (.A1(_12762_),
    .A2(_12780_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27844_ (.A1(net717),
    .A2(net491),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27845_ (.A1(_03800_),
    .A2(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27846_ (.A1(_00804_),
    .A2(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27847_ (.A1(_03800_),
    .A2(net744),
    .A3(_03801_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27848_ (.A1(_03804_),
    .A2(_03803_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27849_ (.A1(_03805_),
    .A2(_03776_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27850_ (.A1(_03803_),
    .A2(_03804_),
    .A3(_03780_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27851_ (.A1(_03807_),
    .A2(_03806_),
    .B(_10525_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27852_ (.I(\text_in_r[8] ),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27853_ (.A1(_03809_),
    .A2(_10431_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27854_ (.A1(_03808_),
    .A2(_03810_),
    .B(\u0.tmp_w[8] ),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27855_ (.A1(_03806_),
    .A2(_03807_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27856_ (.A1(_10405_),
    .A2(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27857_ (.I(\u0.tmp_w[8] ),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27858_ (.I(_03810_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27859_ (.A1(net749),
    .A2(_03814_),
    .A3(_03815_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27860_ (.A1(_03816_),
    .A2(_03811_),
    .ZN(_16048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27861_ (.A1(_12842_),
    .A2(_12840_),
    .A3(\sa03_sr[2] ),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27862_ (.A1(_12839_),
    .A2(_12841_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27863_ (.A1(\sa10_sub[2] ),
    .A2(\sa32_sub[2] ),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27864_ (.A1(_03819_),
    .A2(_12864_),
    .A3(_03818_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27865_ (.A1(_03817_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27866_ (.A1(_12770_),
    .A2(_03821_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27867_ (.A1(_03817_),
    .A2(_12777_),
    .A3(_03820_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27868_ (.A1(_03822_),
    .A2(_03823_),
    .B(_11202_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27869_ (.I(\text_in_r[10] ),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27870_ (.A1(_03825_),
    .A2(net475),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27871_ (.A1(_03824_),
    .A2(_03826_),
    .B(\u0.tmp_w[10] ),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27872_ (.A1(_03822_),
    .A2(_03823_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27873_ (.A1(net811),
    .A2(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27874_ (.I(_03826_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27875_ (.A1(_03829_),
    .A2(_07615_),
    .A3(_03830_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27876_ (.A1(_03827_),
    .A2(_03831_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _27877_ (.I(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27878_ (.I(_03833_),
    .Z(_16064_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27879_ (.A1(_03793_),
    .A2(_03791_),
    .B(_03797_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27880_ (.A1(_03796_),
    .A2(\u0.tmp_w[9] ),
    .A3(_03798_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27881_ (.A1(_03835_),
    .A2(_03834_),
    .ZN(_16038_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27882_ (.I(_03832_),
    .Z(_16057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27883_ (.I(_16039_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27884_ (.A1(_16057_),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27885_ (.A1(_12882_),
    .A2(_00890_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27886_ (.A1(\sa10_sub[3] ),
    .A2(\sa03_sr[3] ),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27887_ (.A1(_03838_),
    .A2(_03839_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27888_ (.I(_03840_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27889_ (.A1(_12839_),
    .A2(_03773_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27890_ (.A1(\sa32_sub[2] ),
    .A2(_13067_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27891_ (.A1(_03842_),
    .A2(_03843_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27892_ (.A1(_03841_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27893_ (.I(_03844_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27894_ (.A1(_03846_),
    .A2(_03840_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27895_ (.A1(_03845_),
    .A2(_03847_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27896_ (.A1(\sa32_sub[3] ),
    .A2(_00881_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27897_ (.A1(_03848_),
    .A2(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27898_ (.A1(_12868_),
    .A2(_00881_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27899_ (.A1(_03845_),
    .A2(_03847_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27900_ (.A1(_03851_),
    .A2(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27901_ (.A1(_03850_),
    .A2(_03853_),
    .A3(_14333_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27902_ (.A1(_11203_),
    .A2(\text_in_r[11] ),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27903_ (.A1(_03854_),
    .A2(_03855_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27904_ (.I(\u0.tmp_w[11] ),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27905_ (.A1(_03856_),
    .A2(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27906_ (.A1(_03854_),
    .A2(\u0.tmp_w[11] ),
    .A3(_03855_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27907_ (.A1(_03858_),
    .A2(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27908_ (.I(_03860_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27909_ (.A1(_03837_),
    .A2(_03861_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27910_ (.A1(_00918_),
    .A2(_00916_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27911_ (.I(_12955_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27912_ (.A1(\sa32_sub[3] ),
    .A2(_13067_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27913_ (.A1(_03864_),
    .A2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _27914_ (.A1(\sa32_sub[3] ),
    .A2(net54),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27915_ (.A1(_03867_),
    .A2(_12955_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27916_ (.A1(_03866_),
    .A2(_03868_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27917_ (.A1(_03863_),
    .A2(_03869_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27918_ (.A1(_03863_),
    .A2(_03869_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27919_ (.A1(_03870_),
    .A2(_13010_),
    .A3(_03871_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27920_ (.A1(_11385_),
    .A2(\text_in_r[12] ),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27921_ (.A1(_03872_),
    .A2(_03873_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27922_ (.A1(_03874_),
    .A2(\u0.tmp_w[12] ),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27923_ (.I(\u0.tmp_w[12] ),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27924_ (.A1(_03872_),
    .A2(_03876_),
    .A3(_03873_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27925_ (.A1(_03877_),
    .A2(_03875_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27926_ (.A1(_03862_),
    .A2(net64),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _27927_ (.I(_16040_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27928_ (.A1(_03832_),
    .A2(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27929_ (.A1(_03861_),
    .A2(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _27930_ (.I(_03882_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27931_ (.A1(_16064_),
    .A2(_16039_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27932_ (.A1(_03883_),
    .A2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27933_ (.I(_16049_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27934_ (.A1(_16064_),
    .A2(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27935_ (.I(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27936_ (.A1(_03856_),
    .A2(\u0.tmp_w[11] ),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27937_ (.A1(_03854_),
    .A2(_03857_),
    .A3(_03855_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27938_ (.A1(_03890_),
    .A2(_03889_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27939_ (.I(net753),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27940_ (.I(_03892_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27941_ (.A1(_03888_),
    .A2(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27942_ (.A1(_03879_),
    .A2(_03885_),
    .A3(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27943_ (.A1(net9),
    .A2(_03833_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27944_ (.I(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27945_ (.I(net753),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27946_ (.A1(_03897_),
    .A2(_03898_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27947_ (.I(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27948_ (.I(_03881_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27949_ (.A1(_03898_),
    .A2(_03901_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27950_ (.A1(net52),
    .A2(net53),
    .A3(_03880_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27951_ (.A1(_03903_),
    .A2(_03861_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27952_ (.A1(_03902_),
    .A2(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27953_ (.A1(_03874_),
    .A2(_03876_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27954_ (.A1(_03872_),
    .A2(\u0.tmp_w[12] ),
    .A3(_03873_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27955_ (.A1(_03906_),
    .A2(_03907_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27956_ (.I(_03908_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27957_ (.I(_03909_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27958_ (.A1(_03900_),
    .A2(_03905_),
    .B(_03910_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27959_ (.A1(\sa32_sub[5] ),
    .A2(_00921_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27960_ (.A1(_03912_),
    .A2(_13004_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27961_ (.A1(_03912_),
    .A2(_13004_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27962_ (.A1(_03913_),
    .A2(_03914_),
    .A3(_11279_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27963_ (.A1(_10411_),
    .A2(\text_in_r[13] ),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27964_ (.A1(_03915_),
    .A2(_03916_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27965_ (.A1(_03917_),
    .A2(\u0.tmp_w[13] ),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27966_ (.I(\u0.tmp_w[13] ),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27967_ (.A1(_03915_),
    .A2(_03919_),
    .A3(_03916_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27968_ (.A1(_03918_),
    .A2(_03920_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27969_ (.I(_03921_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27970_ (.A1(_03895_),
    .A2(_03911_),
    .A3(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27971_ (.A1(_03810_),
    .A2(_03808_),
    .B(_03814_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27972_ (.A1(_03815_),
    .A2(\u0.tmp_w[8] ),
    .A3(_03813_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27973_ (.A1(_03925_),
    .A2(_03924_),
    .ZN(_16037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27974_ (.A1(net9),
    .A2(net724),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _27975_ (.I(_03832_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27976_ (.A1(net59),
    .A2(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27977_ (.A1(_03926_),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27978_ (.I(_03861_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27979_ (.A1(_03929_),
    .A2(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27980_ (.A1(_03928_),
    .A2(_03891_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27981_ (.I(_03932_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27982_ (.A1(_03933_),
    .A2(_03926_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27983_ (.I(_03909_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27984_ (.A1(_03931_),
    .A2(_03934_),
    .A3(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27985_ (.A1(_03881_),
    .A2(net753),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27986_ (.A1(_03833_),
    .A2(_16053_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27987_ (.A1(_03937_),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27988_ (.I(_03878_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27989_ (.I(_03860_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27990_ (.I(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27991_ (.A1(_16057_),
    .A2(_16049_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27992_ (.A1(_03884_),
    .A2(_03942_),
    .A3(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27993_ (.A1(_03939_),
    .A2(_03940_),
    .A3(_03944_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _27994_ (.I(_03921_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _27995_ (.I(_03946_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27996_ (.A1(_03936_),
    .A2(_03945_),
    .A3(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27997_ (.A1(\sa10_sub[6] ),
    .A2(\sa32_sub[6] ),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27998_ (.A1(_03949_),
    .A2(_01000_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27999_ (.A1(_03949_),
    .A2(_01000_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28000_ (.A1(_03950_),
    .A2(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28001_ (.A1(_12958_),
    .A2(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28002_ (.A1(_03953_),
    .A2(_13010_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28003_ (.A1(_10585_),
    .A2(\text_in_r[14] ),
    .B(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28004_ (.I(\u0.tmp_w[14] ),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28005_ (.A1(_03955_),
    .A2(_03956_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28006_ (.A1(_03955_),
    .A2(_03956_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28007_ (.A1(_03957_),
    .A2(_03958_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28008_ (.I(_03959_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28009_ (.A1(_03923_),
    .A2(_03948_),
    .A3(_03960_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28010_ (.I(_16055_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28011_ (.A1(net52),
    .A2(net53),
    .A3(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28012_ (.A1(_03883_),
    .A2(net1052),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28013_ (.A1(net742),
    .A2(net729),
    .A3(_16044_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28014_ (.A1(_03898_),
    .A2(_03965_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28015_ (.A1(net713),
    .A2(net91),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28016_ (.I(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28017_ (.A1(_03966_),
    .A2(_03968_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28018_ (.A1(_03964_),
    .A2(_03969_),
    .A3(_03935_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28019_ (.A1(_03860_),
    .A2(_03965_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28020_ (.I(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28021_ (.I(_16046_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28022_ (.A1(net91),
    .A2(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28023_ (.A1(_03972_),
    .A2(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28024_ (.A1(net714),
    .A2(_03833_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28025_ (.A1(net751),
    .A2(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28026_ (.A1(_03975_),
    .A2(_03940_),
    .A3(_03977_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28027_ (.A1(_03970_),
    .A2(_03978_),
    .A3(_03947_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28028_ (.A1(_16057_),
    .A2(_16041_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28029_ (.A1(_03980_),
    .A2(_03892_),
    .B(_03908_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28030_ (.A1(_16053_),
    .A2(_03927_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28031_ (.A1(_03976_),
    .A2(_03930_),
    .A3(net1057),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28032_ (.A1(_03981_),
    .A2(_03983_),
    .A3(_03899_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28033_ (.A1(_16038_),
    .A2(_03927_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28034_ (.I(_03898_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28035_ (.A1(_03985_),
    .A2(_03986_),
    .A3(_03965_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28036_ (.A1(_03962_),
    .A2(_03927_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28037_ (.A1(_03976_),
    .A2(_03942_),
    .A3(_03988_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28038_ (.I(_03909_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28039_ (.A1(_03987_),
    .A2(_03989_),
    .A3(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28040_ (.A1(_03984_),
    .A2(_03991_),
    .A3(_03922_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28041_ (.I(_03959_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28042_ (.I(_03993_),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28043_ (.A1(_03979_),
    .A2(_03992_),
    .A3(_03994_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _28044_ (.A1(net54),
    .A2(net975),
    .A3(_13007_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28045_ (.A1(_11385_),
    .A2(\text_in_r[15] ),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28046_ (.A1(_03996_),
    .A2(_10585_),
    .B(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28047_ (.A1(\u0.tmp_w[15] ),
    .A2(_03998_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28048_ (.I(_03999_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28049_ (.A1(_03961_),
    .A2(_03995_),
    .A3(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28050_ (.I(_03878_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28051_ (.A1(_03833_),
    .A2(_16046_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28052_ (.I(_16044_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28053_ (.A1(_16057_),
    .A2(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28054_ (.A1(_04003_),
    .A2(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28055_ (.A1(_04006_),
    .A2(_03892_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _28056_ (.I(_03861_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28057_ (.A1(_16057_),
    .A2(_16039_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28058_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04009_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28059_ (.A1(net90),
    .A2(_16041_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28060_ (.A1(_04011_),
    .A2(_03930_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _28061_ (.A1(_04002_),
    .A2(_04007_),
    .A3(_04010_),
    .A4(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28062_ (.I(_03898_),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28063_ (.A1(net742),
    .A2(net732),
    .A3(net729),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28064_ (.A1(_03898_),
    .A2(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28065_ (.A1(_16062_),
    .A2(_04014_),
    .B(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28066_ (.I(_03946_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28067_ (.A1(_04017_),
    .A2(_03935_),
    .B(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28068_ (.A1(_04013_),
    .A2(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28069_ (.A1(net91),
    .A2(_16044_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28070_ (.A1(_04021_),
    .A2(_03861_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28071_ (.I(_16051_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28072_ (.A1(net742),
    .A2(_04023_),
    .A3(net728),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28073_ (.A1(_04022_),
    .A2(net730),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28074_ (.I(_03878_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28075_ (.A1(_03980_),
    .A2(_04014_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28076_ (.A1(_04025_),
    .A2(_04026_),
    .A3(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28077_ (.A1(_04005_),
    .A2(_03861_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28078_ (.A1(_03980_),
    .A2(_04008_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28079_ (.A1(_04029_),
    .A2(_04030_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _28080_ (.I(_03898_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28081_ (.A1(_03888_),
    .A2(_04032_),
    .B(net64),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28082_ (.A1(_04031_),
    .A2(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28083_ (.I(_03946_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28084_ (.A1(_04028_),
    .A2(_04034_),
    .A3(_04035_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28085_ (.A1(_04020_),
    .A2(_03960_),
    .A3(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28086_ (.I(_04003_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28087_ (.I(_03908_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28088_ (.A1(_04038_),
    .A2(_03986_),
    .B(_04039_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28089_ (.A1(_04040_),
    .A2(_03983_),
    .B(_04018_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28090_ (.A1(net91),
    .A2(_16051_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28091_ (.A1(_04003_),
    .A2(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28092_ (.A1(_04043_),
    .A2(_04032_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28093_ (.A1(_04044_),
    .A2(_03882_),
    .A3(_03990_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28094_ (.A1(_04041_),
    .A2(_04045_),
    .B(_03959_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28095_ (.A1(net742),
    .A2(net728),
    .A3(_16049_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28096_ (.A1(net59),
    .A2(net90),
    .B(_03942_),
    .C(_04047_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28097_ (.A1(net60),
    .A2(_03927_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28098_ (.I(_03891_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28099_ (.A1(_04049_),
    .A2(_04050_),
    .A3(_04015_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28100_ (.A1(_04048_),
    .A2(_03940_),
    .A3(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28101_ (.I(_03980_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28102_ (.A1(net90),
    .A2(_03836_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28103_ (.A1(_04053_),
    .A2(_04054_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28104_ (.A1(_04055_),
    .A2(_03986_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28105_ (.I(_03941_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28106_ (.A1(_03974_),
    .A2(_04057_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28107_ (.A1(_04056_),
    .A2(_03910_),
    .A3(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28108_ (.A1(_04052_),
    .A2(_04059_),
    .A3(_04035_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28109_ (.A1(_04046_),
    .A2(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _28110_ (.I(_04000_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28111_ (.A1(_04037_),
    .A2(_04061_),
    .A3(_04062_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28112_ (.A1(_04001_),
    .A2(_04063_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28113_ (.I(_03878_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28114_ (.A1(_03980_),
    .A2(_04014_),
    .B(_04064_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28115_ (.I(_03904_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28116_ (.A1(_04066_),
    .A2(_04009_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28117_ (.A1(_03833_),
    .A2(net750),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28118_ (.I(_04068_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28119_ (.A1(_04069_),
    .A2(_04032_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28120_ (.A1(_04065_),
    .A2(_04067_),
    .A3(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28121_ (.A1(_03896_),
    .A2(_03930_),
    .A3(_03974_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28122_ (.A1(_03884_),
    .A2(_03928_),
    .A3(_04032_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28123_ (.A1(_04072_),
    .A2(_04073_),
    .A3(_04026_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28124_ (.A1(_04071_),
    .A2(_04074_),
    .A3(_04035_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28125_ (.A1(_03882_),
    .A2(_04064_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28126_ (.A1(_03976_),
    .A2(_03986_),
    .A3(net1058),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28127_ (.A1(_04076_),
    .A2(_04077_),
    .B(_04018_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28128_ (.I(_16053_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28129_ (.A1(_16064_),
    .A2(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28130_ (.A1(_04080_),
    .A2(_03881_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28131_ (.A1(_04081_),
    .A2(_03942_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28132_ (.I(_16041_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28133_ (.A1(net52),
    .A2(net53),
    .A3(_04083_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28134_ (.A1(_04084_),
    .A2(_03891_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28135_ (.I(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28136_ (.A1(_04086_),
    .A2(_03988_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28137_ (.A1(_04082_),
    .A2(_04087_),
    .A3(_03910_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28138_ (.A1(_04078_),
    .A2(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28139_ (.A1(_04075_),
    .A2(_04089_),
    .B(_03960_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28140_ (.A1(_03982_),
    .A2(_04047_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28141_ (.A1(_04091_),
    .A2(_03861_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28142_ (.I(_16065_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28143_ (.A1(_03921_),
    .A2(_03942_),
    .A3(_04093_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28144_ (.A1(_04092_),
    .A2(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28145_ (.A1(_04095_),
    .A2(_03935_),
    .B(_03959_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28146_ (.A1(_04072_),
    .A2(_03990_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28147_ (.A1(_16043_),
    .A2(_03833_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28148_ (.A1(_03933_),
    .A2(_04098_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _28149_ (.A1(_04097_),
    .A2(_04099_),
    .A3(_04035_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28150_ (.A1(_03972_),
    .A2(net1059),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28151_ (.A1(_03884_),
    .A2(_03967_),
    .A3(_04032_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28152_ (.A1(_03946_),
    .A2(_03909_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28153_ (.A1(_04101_),
    .A2(_04102_),
    .A3(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _28154_ (.A1(_04096_),
    .A2(_04100_),
    .A3(_04104_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28155_ (.A1(_04090_),
    .A2(_04105_),
    .B(_04000_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28156_ (.A1(_04038_),
    .A2(_04032_),
    .B(_04064_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28157_ (.A1(_04050_),
    .A2(_16069_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28158_ (.I(_03985_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28159_ (.A1(_04109_),
    .A2(_03893_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28160_ (.A1(_04107_),
    .A2(_04108_),
    .A3(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28161_ (.A1(_04066_),
    .A2(_03988_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28162_ (.A1(_04007_),
    .A2(_04112_),
    .A3(_04026_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28163_ (.A1(_04111_),
    .A2(_04113_),
    .A3(_03922_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28164_ (.A1(_03941_),
    .A2(net90),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28165_ (.A1(_04115_),
    .A2(_04004_),
    .B(_04039_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28166_ (.A1(_04049_),
    .A2(_03891_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28167_ (.A1(_04117_),
    .A2(_03926_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28168_ (.A1(_04116_),
    .A2(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28169_ (.A1(_04068_),
    .A2(_03986_),
    .A3(_03974_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28170_ (.A1(_03976_),
    .A2(net51),
    .A3(_03942_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28171_ (.A1(_04120_),
    .A2(_04121_),
    .A3(_03990_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28172_ (.A1(_04119_),
    .A2(_04122_),
    .A3(_04035_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28173_ (.A1(_04114_),
    .A2(_04123_),
    .A3(_03960_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28174_ (.A1(_16057_),
    .A2(_16046_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28175_ (.A1(_04125_),
    .A2(_04032_),
    .B(_04039_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28176_ (.I(_03921_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28177_ (.A1(_04126_),
    .A2(_04082_),
    .B(_04127_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28178_ (.A1(_03941_),
    .A2(net1052),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28179_ (.A1(_04109_),
    .A2(_04129_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28180_ (.A1(_16057_),
    .A2(_04079_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28181_ (.A1(_04131_),
    .A2(_03986_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28182_ (.A1(_04130_),
    .A2(_03990_),
    .A3(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28183_ (.A1(_04128_),
    .A2(_04133_),
    .B(_03959_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28184_ (.A1(_03883_),
    .A2(_04003_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28185_ (.A1(_04068_),
    .A2(_04050_),
    .A3(_03837_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28186_ (.A1(_04135_),
    .A2(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28187_ (.A1(_04137_),
    .A2(_03935_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28188_ (.A1(net60),
    .A2(net59),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28189_ (.A1(_04139_),
    .A2(_03967_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28190_ (.A1(_04140_),
    .A2(_04057_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28191_ (.A1(_04016_),
    .A2(_03968_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28192_ (.A1(_04141_),
    .A2(_04142_),
    .A3(_04026_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28193_ (.A1(_04138_),
    .A2(_04143_),
    .A3(_04127_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28194_ (.A1(_04134_),
    .A2(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28195_ (.A1(_04124_),
    .A2(_04062_),
    .A3(_04145_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28196_ (.A1(_04106_),
    .A2(_04146_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28197_ (.A1(_03974_),
    .A2(_03898_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28198_ (.I(_03963_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28199_ (.A1(_04147_),
    .A2(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _28200_ (.A1(net9),
    .A2(net90),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28201_ (.A1(_03971_),
    .A2(_04150_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28202_ (.I(_03908_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28203_ (.A1(_04149_),
    .A2(_04151_),
    .B(_04152_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28204_ (.A1(_04003_),
    .A2(_03930_),
    .A3(_04005_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28205_ (.I(_03878_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28206_ (.A1(_04051_),
    .A2(_04154_),
    .A3(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28207_ (.A1(_04153_),
    .A2(_04156_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28208_ (.A1(_04157_),
    .A2(_03922_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28209_ (.A1(_04011_),
    .A2(_03928_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28210_ (.A1(_04159_),
    .A2(_04057_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28211_ (.A1(_04098_),
    .A2(net51),
    .A3(_04014_),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28212_ (.A1(_04160_),
    .A2(_04161_),
    .A3(_03910_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28213_ (.A1(_03938_),
    .A2(_03941_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28214_ (.I(_03988_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28215_ (.A1(_04163_),
    .A2(_04164_),
    .B(_04026_),
    .C(_03966_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28216_ (.A1(_04162_),
    .A2(_04165_),
    .A3(_03947_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28217_ (.A1(_04158_),
    .A2(_04166_),
    .A3(_03960_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28218_ (.A1(net52),
    .A2(net53),
    .A3(_16055_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28219_ (.I(_04168_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28220_ (.A1(_03932_),
    .A2(_04169_),
    .B(_03908_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28221_ (.A1(_03896_),
    .A2(_03930_),
    .A3(_04042_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28222_ (.A1(_04170_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28223_ (.A1(_03967_),
    .A2(_03892_),
    .A3(net730),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28224_ (.A1(net51),
    .A2(_03942_),
    .A3(_04015_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28225_ (.A1(_04173_),
    .A2(_04174_),
    .B(_04152_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28226_ (.A1(_04172_),
    .A2(_04175_),
    .B(_03947_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28227_ (.A1(net52),
    .A2(net53),
    .A3(net1056),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28228_ (.A1(_03941_),
    .A2(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28229_ (.A1(_04178_),
    .A2(_03985_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28230_ (.A1(_04044_),
    .A2(_04179_),
    .A3(_03940_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28231_ (.A1(_04178_),
    .A2(_03967_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28232_ (.A1(_04042_),
    .A2(_04168_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28233_ (.A1(_04182_),
    .A2(_04014_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28234_ (.A1(_04181_),
    .A2(_04183_),
    .A3(_03990_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28235_ (.A1(_04180_),
    .A2(_04184_),
    .A3(_04127_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28236_ (.A1(_04176_),
    .A2(_04185_),
    .A3(_03994_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28237_ (.A1(_04167_),
    .A2(_04186_),
    .A3(_04000_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28238_ (.I(_04151_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28239_ (.A1(_16071_),
    .A2(_04032_),
    .B(_04064_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28240_ (.A1(_04188_),
    .A2(_04189_),
    .B(_04018_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28241_ (.A1(_04050_),
    .A2(_16060_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28242_ (.A1(_04191_),
    .A2(_03940_),
    .A3(_03966_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28243_ (.I(_03993_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28244_ (.A1(_04190_),
    .A2(_04192_),
    .B(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28245_ (.A1(_03883_),
    .A2(_04177_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28246_ (.A1(_04195_),
    .A2(_03879_),
    .B(_04127_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28247_ (.I(_04163_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28248_ (.A1(_04083_),
    .A2(_03973_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28249_ (.A1(_04198_),
    .A2(net91),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28250_ (.A1(_04197_),
    .A2(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28251_ (.A1(_04200_),
    .A2(_03935_),
    .A3(_04092_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28252_ (.A1(_04201_),
    .A2(_04196_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28253_ (.A1(_04202_),
    .A2(_04194_),
    .B(_04000_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28254_ (.A1(_03926_),
    .A2(_04049_),
    .A3(_03941_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28255_ (.A1(_04204_),
    .A2(_04064_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28256_ (.A1(_03893_),
    .A2(_04093_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28257_ (.A1(_04205_),
    .A2(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28258_ (.A1(_04049_),
    .A2(_04054_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28259_ (.A1(_04208_),
    .A2(_03893_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28260_ (.A1(_16057_),
    .A2(_03886_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28261_ (.A1(_04210_),
    .A2(_04015_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28262_ (.A1(_04211_),
    .A2(_04057_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28263_ (.A1(_04209_),
    .A2(_04212_),
    .A3(_03910_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28264_ (.A1(_04207_),
    .A2(_03922_),
    .A3(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28265_ (.A1(_03896_),
    .A2(_03941_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28266_ (.A1(_04215_),
    .A2(_03967_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28267_ (.A1(_04216_),
    .A2(_03910_),
    .A3(_04051_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28268_ (.A1(_03892_),
    .A2(_16062_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28269_ (.A1(_03903_),
    .A2(_04022_),
    .B(_04218_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28270_ (.A1(_04219_),
    .A2(_04002_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28271_ (.A1(_04217_),
    .A2(_04220_),
    .A3(_04035_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28272_ (.A1(_04214_),
    .A2(_04221_),
    .A3(_03994_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28273_ (.A1(_04222_),
    .A2(_04203_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28274_ (.A1(_04187_),
    .A2(_04223_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28275_ (.A1(_03972_),
    .A2(_03943_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28276_ (.A1(net1057),
    .A2(_03892_),
    .A3(net712),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28277_ (.A1(_04224_),
    .A2(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28278_ (.A1(_04226_),
    .A2(_04155_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28279_ (.A1(_03937_),
    .A2(_03887_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28280_ (.A1(_03931_),
    .A2(_04228_),
    .A3(_04152_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28281_ (.A1(_04227_),
    .A2(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28282_ (.A1(_04230_),
    .A2(_03994_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28283_ (.A1(_04178_),
    .A2(_03988_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28284_ (.A1(net743),
    .A2(_16057_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28285_ (.A1(_03896_),
    .A2(_04014_),
    .A3(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28286_ (.A1(_04232_),
    .A2(_04234_),
    .A3(_03940_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28287_ (.A1(_04068_),
    .A2(_04050_),
    .A3(_04210_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28288_ (.A1(_03837_),
    .A2(_03930_),
    .A3(net712),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28289_ (.A1(_04236_),
    .A2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28290_ (.A1(_04238_),
    .A2(_03935_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28291_ (.A1(_04235_),
    .A2(_04239_),
    .A3(_03960_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28292_ (.A1(_04231_),
    .A2(_03947_),
    .A3(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28293_ (.A1(_03904_),
    .A2(_04039_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28294_ (.A1(_03896_),
    .A2(_04014_),
    .A3(_03967_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28295_ (.A1(_04242_),
    .A2(_04243_),
    .B(_03993_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _28296_ (.A1(net9),
    .A2(net59),
    .B(_03928_),
    .C(_04050_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28297_ (.A1(_03896_),
    .A2(net51),
    .A3(_04057_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28298_ (.A1(_04245_),
    .A2(_04246_),
    .A3(_03940_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28299_ (.A1(_04244_),
    .A2(_04247_),
    .B(_04035_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28300_ (.A1(_04245_),
    .A2(_04002_),
    .A3(_03971_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28301_ (.A1(net752),
    .A2(net730),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28302_ (.I(_04250_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28303_ (.A1(_04251_),
    .A2(_04233_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28304_ (.A1(_04130_),
    .A2(_04252_),
    .A3(_03910_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28305_ (.A1(_04249_),
    .A2(_04193_),
    .A3(_04253_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28306_ (.A1(_04248_),
    .A2(_04254_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28307_ (.A1(_04241_),
    .A2(_04255_),
    .A3(_04062_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28308_ (.A1(_04118_),
    .A2(_04010_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28309_ (.A1(_04257_),
    .A2(_04155_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28310_ (.A1(_03937_),
    .A2(_03963_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28311_ (.A1(_03976_),
    .A2(_04042_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28312_ (.A1(_04260_),
    .A2(_04008_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28313_ (.A1(_04259_),
    .A2(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28314_ (.A1(_04262_),
    .A2(_04152_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28315_ (.A1(_04263_),
    .A2(_04035_),
    .A3(_04258_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28316_ (.A1(_04170_),
    .A2(_03921_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28317_ (.A1(_03860_),
    .A2(_04024_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28318_ (.I(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28319_ (.A1(_04267_),
    .A2(_04199_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28320_ (.A1(_04092_),
    .A2(_04268_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28321_ (.A1(_04269_),
    .A2(_04155_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28322_ (.A1(_04265_),
    .A2(_04270_),
    .B(_03959_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28323_ (.A1(_04264_),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28324_ (.A1(_04199_),
    .A2(_03861_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28325_ (.A1(_04273_),
    .A2(_04148_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28326_ (.A1(_03976_),
    .A2(_03881_),
    .A3(_03898_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28327_ (.A1(_04274_),
    .A2(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28328_ (.A1(_04276_),
    .A2(_04018_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28329_ (.I(_04042_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28330_ (.A1(_04278_),
    .A2(_03941_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28331_ (.A1(_04173_),
    .A2(_03946_),
    .A3(_04279_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28332_ (.A1(_04277_),
    .A2(_04280_),
    .B(_04002_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28333_ (.A1(_03898_),
    .A2(_04047_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _28334_ (.A1(_04282_),
    .A2(_04150_),
    .A3(_03946_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28335_ (.A1(_03902_),
    .A2(_03921_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28336_ (.A1(_04283_),
    .A2(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28337_ (.I(_03903_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28338_ (.A1(_03921_),
    .A2(_04008_),
    .A3(_04286_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28339_ (.A1(_04030_),
    .A2(_03909_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28340_ (.A1(_04287_),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28341_ (.A1(_04285_),
    .A2(_04289_),
    .B(_04193_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28342_ (.A1(_04290_),
    .A2(_04281_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28343_ (.A1(_04291_),
    .A2(_04272_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28344_ (.A1(_04292_),
    .A2(_04000_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28345_ (.A1(_04256_),
    .A2(_04293_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28346_ (.A1(_04056_),
    .A2(_03931_),
    .B(_03990_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28347_ (.A1(_03985_),
    .A2(_04139_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28348_ (.A1(_04295_),
    .A2(_04050_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28349_ (.A1(_04267_),
    .A2(_03928_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28350_ (.A1(_04296_),
    .A2(_04297_),
    .B(_04026_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28351_ (.A1(_04294_),
    .A2(_04298_),
    .B(_03960_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28352_ (.A1(_03933_),
    .A2(net1055),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28353_ (.A1(_04115_),
    .A2(_04039_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28354_ (.A1(_04300_),
    .A2(_04301_),
    .B(_03959_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28355_ (.A1(_04098_),
    .A2(_03986_),
    .A3(_04009_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28356_ (.A1(_04072_),
    .A2(_04303_),
    .A3(_03910_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28357_ (.A1(_04302_),
    .A2(_04304_),
    .B(_04062_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28358_ (.A1(_04299_),
    .A2(_04305_),
    .B(_03947_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28359_ (.A1(_04007_),
    .A2(_04064_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28360_ (.A1(_04215_),
    .A2(_04009_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28361_ (.A1(_04307_),
    .A2(_04308_),
    .B(_04193_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28362_ (.A1(_04022_),
    .A2(_03896_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _28363_ (.A1(_04310_),
    .A2(_04155_),
    .A3(_04149_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28364_ (.A1(_04309_),
    .A2(_04311_),
    .B(_04000_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28365_ (.A1(_03893_),
    .A2(_04208_),
    .B(_04296_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28366_ (.A1(_04313_),
    .A2(_03935_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28367_ (.I(_04099_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28368_ (.A1(_04205_),
    .A2(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28369_ (.A1(_04314_),
    .A2(_03994_),
    .A3(_04316_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28370_ (.A1(_04312_),
    .A2(_04317_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28371_ (.A1(_04306_),
    .A2(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28372_ (.A1(_03892_),
    .A2(_04079_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28373_ (.A1(_04015_),
    .A2(_04008_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28374_ (.A1(_04320_),
    .A2(_04321_),
    .A3(net64),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28375_ (.A1(_04322_),
    .A2(_04193_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28376_ (.A1(_04029_),
    .A2(_03909_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28377_ (.A1(_04267_),
    .A2(_03985_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28378_ (.A1(_04324_),
    .A2(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28379_ (.A1(_04323_),
    .A2(_04326_),
    .B(_04062_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28380_ (.I(_04015_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28381_ (.A1(_04328_),
    .A2(_04147_),
    .B(_03983_),
    .C(_04026_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28382_ (.A1(_04163_),
    .A2(_03909_),
    .A3(_04085_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28383_ (.A1(_04330_),
    .A2(_03959_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28384_ (.A1(_04329_),
    .A2(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28385_ (.A1(_04327_),
    .A2(_04332_),
    .B(_03922_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28386_ (.A1(_04098_),
    .A2(_03930_),
    .A3(_03967_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28387_ (.A1(_04334_),
    .A2(_04102_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28388_ (.A1(_04266_),
    .A2(_04053_),
    .B(_04064_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _28389_ (.A1(_04002_),
    .A2(_04335_),
    .B(_04336_),
    .C(_03959_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28390_ (.A1(_04279_),
    .A2(_03909_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28391_ (.A1(_04328_),
    .A2(_03941_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28392_ (.I(_04339_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28393_ (.A1(_04340_),
    .A2(_04044_),
    .A3(_04338_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28394_ (.A1(_03988_),
    .A2(_03891_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28395_ (.A1(_04342_),
    .A2(net712),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28396_ (.A1(_04025_),
    .A2(_04343_),
    .A3(_04026_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28397_ (.A1(_04344_),
    .A2(_04341_),
    .B(_04193_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28398_ (.A1(_04345_),
    .A2(_04337_),
    .B(_04062_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28399_ (.A1(_04346_),
    .A2(_04333_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28400_ (.A1(_04347_),
    .A2(_04319_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28401_ (.A1(_03974_),
    .A2(_04008_),
    .A3(_03963_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28402_ (.A1(_03981_),
    .A2(_03899_),
    .A3(_04348_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28403_ (.A1(_04021_),
    .A2(_03892_),
    .A3(net731),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28404_ (.I(_04198_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28405_ (.A1(_04008_),
    .A2(_04177_),
    .A3(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28406_ (.A1(_04350_),
    .A2(_04352_),
    .A3(_04039_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28407_ (.A1(_04349_),
    .A2(_04018_),
    .A3(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28408_ (.I(_03937_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28409_ (.A1(_04355_),
    .A2(_04064_),
    .A3(_04261_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28410_ (.A1(net90),
    .A2(_04004_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28411_ (.A1(_04147_),
    .A2(_04039_),
    .A3(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28412_ (.A1(_04356_),
    .A2(_03921_),
    .A3(_04358_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28413_ (.A1(_04359_),
    .A2(_04354_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28414_ (.A1(_04360_),
    .A2(_03994_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28415_ (.A1(_04085_),
    .A2(_04150_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28416_ (.A1(_04362_),
    .A2(_04339_),
    .B(_04152_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28417_ (.A1(_03883_),
    .A2(_04054_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28418_ (.A1(_04050_),
    .A2(_04168_),
    .B(_03909_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28419_ (.A1(_04364_),
    .A2(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28420_ (.A1(_04363_),
    .A2(_04127_),
    .A3(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28421_ (.A1(_04091_),
    .A2(_03930_),
    .B(net64),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28422_ (.I(_03977_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28423_ (.A1(_04369_),
    .A2(_04139_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28424_ (.A1(_04368_),
    .A2(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28425_ (.A1(net9),
    .A2(_03930_),
    .B(_03909_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28426_ (.A1(_04296_),
    .A2(_04372_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28427_ (.A1(_04371_),
    .A2(_04373_),
    .A3(_04018_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28428_ (.A1(_04367_),
    .A2(_04374_),
    .A3(_03960_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28429_ (.A1(_04375_),
    .A2(_04361_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28430_ (.A1(_04376_),
    .A2(_04062_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28431_ (.A1(_04107_),
    .A2(_04129_),
    .B(_03993_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28432_ (.A1(net1057),
    .A2(_04014_),
    .A3(_03965_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28433_ (.A1(_04379_),
    .A2(_03940_),
    .A3(_04273_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28434_ (.A1(_04378_),
    .A2(_04380_),
    .B(_04127_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28435_ (.A1(_03972_),
    .A2(net51),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28436_ (.A1(_04251_),
    .A2(_03985_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28437_ (.A1(_04382_),
    .A2(_04383_),
    .B(_04152_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28438_ (.A1(_04008_),
    .A2(net59),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28439_ (.A1(_03934_),
    .A2(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28440_ (.A1(_04386_),
    .A2(_04155_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28441_ (.A1(_04384_),
    .A2(_04387_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28442_ (.A1(_04388_),
    .A2(_04193_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28443_ (.A1(_04381_),
    .A2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28444_ (.A1(_03883_),
    .A2(_04047_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28445_ (.A1(_04233_),
    .A2(_03986_),
    .A3(net1053),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28446_ (.A1(_04391_),
    .A2(_03910_),
    .A3(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28447_ (.A1(net1057),
    .A2(_03892_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28448_ (.A1(_16049_),
    .A2(_03893_),
    .B(_04394_),
    .C(_04155_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28449_ (.A1(_04393_),
    .A2(_04395_),
    .A3(_03959_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28450_ (.A1(_03888_),
    .A2(_04057_),
    .B(_04064_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28451_ (.A1(_04394_),
    .A2(_04148_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28452_ (.A1(_04397_),
    .A2(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28453_ (.A1(_03967_),
    .A2(_04032_),
    .A3(_04177_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28454_ (.A1(_03983_),
    .A2(_04400_),
    .A3(_04026_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28455_ (.A1(_04399_),
    .A2(_04401_),
    .A3(_04193_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28456_ (.A1(_04396_),
    .A2(_04402_),
    .A3(_03922_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28457_ (.A1(_04390_),
    .A2(_04403_),
    .A3(_04000_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28458_ (.A1(_04377_),
    .A2(_04404_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28459_ (.A1(_03933_),
    .A2(_04015_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28460_ (.A1(_04115_),
    .A2(_04351_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28461_ (.A1(_04338_),
    .A2(_04405_),
    .A3(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28462_ (.A1(_04053_),
    .A2(_04080_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28463_ (.A1(_04408_),
    .A2(_04057_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28464_ (.A1(_04251_),
    .A2(_03988_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28465_ (.A1(_04409_),
    .A2(_04410_),
    .A3(_04002_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28466_ (.A1(_04407_),
    .A2(_04411_),
    .A3(_03922_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28467_ (.A1(_04115_),
    .A2(_16041_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28468_ (.A1(_04338_),
    .A2(_03862_),
    .A3(_04413_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28469_ (.A1(_04295_),
    .A2(_04057_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28470_ (.A1(_16058_),
    .A2(_16067_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28471_ (.A1(_04416_),
    .A2(_04014_),
    .B(_04039_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28472_ (.A1(_04415_),
    .A2(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28473_ (.A1(_04414_),
    .A2(_03947_),
    .A3(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28474_ (.A1(_04412_),
    .A2(_04419_),
    .A3(_03994_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28475_ (.A1(_04086_),
    .A2(_04233_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28476_ (.A1(_03972_),
    .A2(_03985_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28477_ (.A1(_04421_),
    .A2(_04422_),
    .A3(_04002_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28478_ (.A1(_04357_),
    .A2(net747),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28479_ (.A1(_04424_),
    .A2(_03893_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28480_ (.A1(_04425_),
    .A2(_03910_),
    .A3(_04191_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28481_ (.A1(_04423_),
    .A2(_04426_),
    .A3(_03947_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28482_ (.A1(_04022_),
    .A2(_04068_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28483_ (.A1(_04199_),
    .A2(_03986_),
    .A3(_04015_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28484_ (.A1(_04428_),
    .A2(_03940_),
    .A3(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28485_ (.A1(_04098_),
    .A2(_03861_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28486_ (.A1(_04431_),
    .A2(_04021_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28487_ (.A1(_04432_),
    .A2(_04033_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28488_ (.A1(_04430_),
    .A2(_04433_),
    .A3(_04127_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28489_ (.A1(_04427_),
    .A2(_04434_),
    .A3(_03960_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28490_ (.A1(_04062_),
    .A2(_04435_),
    .A3(_04420_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28491_ (.A1(_04342_),
    .A2(_04068_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28492_ (.A1(_03926_),
    .A2(_04068_),
    .A3(_04008_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28493_ (.A1(_04437_),
    .A2(_04438_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28494_ (.A1(_04439_),
    .A2(_04152_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28495_ (.A1(_03985_),
    .A2(_04357_),
    .A3(_04050_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28496_ (.A1(_04441_),
    .A2(_04438_),
    .A3(_04155_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28497_ (.A1(_04440_),
    .A2(_04442_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28498_ (.A1(_04443_),
    .A2(_03947_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28499_ (.A1(_03969_),
    .A2(_03990_),
    .A3(_04108_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28500_ (.I(_04233_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28501_ (.A1(_04446_),
    .A2(_03986_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28502_ (.A1(_04261_),
    .A2(_04026_),
    .A3(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28503_ (.A1(_04445_),
    .A2(_04448_),
    .A3(_04127_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28504_ (.A1(_04449_),
    .A2(_03994_),
    .A3(_04444_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28505_ (.A1(_04109_),
    .A2(_04266_),
    .B(_04282_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28506_ (.A1(_04451_),
    .A2(_04152_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28507_ (.A1(_04154_),
    .A2(_04155_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28508_ (.A1(_04452_),
    .A2(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28509_ (.A1(_04454_),
    .A2(_03922_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28510_ (.I(_16059_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28511_ (.A1(_03942_),
    .A2(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28512_ (.A1(_04109_),
    .A2(_04250_),
    .B(_04457_),
    .C(_04155_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28513_ (.A1(_04233_),
    .A2(_03942_),
    .A3(net1054),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28514_ (.A1(_04459_),
    .A2(_04070_),
    .A3(_04152_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28515_ (.A1(_04458_),
    .A2(_04460_),
    .A3(_04035_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28516_ (.A1(_04455_),
    .A2(_04461_),
    .A3(_03960_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28517_ (.A1(_04450_),
    .A2(_04000_),
    .A3(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28518_ (.A1(_04436_),
    .A2(_04463_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _28519_ (.A1(_04109_),
    .A2(_03977_),
    .B1(_03904_),
    .B2(_04446_),
    .C(_03990_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28520_ (.A1(_04278_),
    .A2(_03892_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28521_ (.A1(_04008_),
    .A2(_16067_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28522_ (.A1(_04465_),
    .A2(net64),
    .A3(_04466_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28523_ (.A1(_04286_),
    .A2(_03893_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28524_ (.A1(_04467_),
    .A2(_04468_),
    .B(_04018_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28525_ (.A1(_04464_),
    .A2(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28526_ (.A1(_04324_),
    .A2(_03899_),
    .A3(_04072_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28527_ (.A1(_04079_),
    .A2(_03942_),
    .B(_04039_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28528_ (.A1(_04472_),
    .A2(_04012_),
    .B(_04127_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28529_ (.A1(_04471_),
    .A2(_04473_),
    .B(_04193_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28530_ (.A1(_04474_),
    .A2(_04470_),
    .B(_04000_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28531_ (.A1(_04431_),
    .A2(_04086_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28532_ (.A1(_03921_),
    .A2(_04009_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28533_ (.A1(_04476_),
    .A2(_04477_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28534_ (.A1(_03938_),
    .A2(_04014_),
    .A3(_04009_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28535_ (.A1(_04233_),
    .A2(_04057_),
    .A3(_04047_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28536_ (.A1(_04479_),
    .A2(_04480_),
    .B(_04127_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28537_ (.A1(_04478_),
    .A2(_04481_),
    .B(_04002_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28538_ (.A1(net1060),
    .A2(_03893_),
    .B(_03946_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28539_ (.A1(_04483_),
    .A2(_04415_),
    .B(_03940_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28540_ (.A1(_04117_),
    .A2(_03938_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28541_ (.A1(_04485_),
    .A2(_04018_),
    .A3(_04268_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28542_ (.A1(_04484_),
    .A2(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28543_ (.A1(_04482_),
    .A2(_03994_),
    .A3(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28544_ (.A1(_04475_),
    .A2(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28545_ (.A1(_03902_),
    .A2(_04064_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28546_ (.A1(_04131_),
    .A2(_04057_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28547_ (.A1(_04490_),
    .A2(_04491_),
    .B(_04018_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28548_ (.A1(_03893_),
    .A2(_04081_),
    .B(_04022_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28549_ (.A1(_04493_),
    .A2(_03935_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28550_ (.A1(_04494_),
    .A2(_04492_),
    .B(_04193_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28551_ (.A1(_04050_),
    .A2(net718),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28552_ (.A1(_04334_),
    .A2(_04039_),
    .A3(_04496_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28553_ (.A1(_03985_),
    .A2(_03938_),
    .A3(_04032_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28554_ (.A1(_04204_),
    .A2(_04498_),
    .B(_04152_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28555_ (.A1(_04497_),
    .A2(_04499_),
    .B(_04035_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28556_ (.A1(_04500_),
    .A2(_04495_),
    .B(_04062_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28557_ (.A1(_04369_),
    .A2(_04021_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28558_ (.A1(_04197_),
    .A2(_04009_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28559_ (.A1(_04502_),
    .A2(_04503_),
    .A3(_03935_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28560_ (.I(_04342_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28561_ (.A1(_04325_),
    .A2(_04002_),
    .A3(_04505_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28562_ (.A1(_04504_),
    .A2(_04506_),
    .A3(_03947_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28563_ (.A1(_04216_),
    .A2(_04002_),
    .A3(_04410_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28564_ (.A1(_04112_),
    .A2(_04275_),
    .A3(_03990_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28565_ (.A1(_04508_),
    .A2(_03922_),
    .A3(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28566_ (.A1(_04507_),
    .A2(_04510_),
    .A3(_03994_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28567_ (.A1(_04511_),
    .A2(_04501_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28568_ (.A1(_04512_),
    .A2(_04489_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28569_ (.A1(_01564_),
    .A2(_01588_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28570_ (.A1(net1117),
    .A2(_01560_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28571_ (.A1(_04513_),
    .A2(_04514_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28572_ (.A1(_10351_),
    .A2(net615),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28573_ (.A1(net876),
    .A2(_10342_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28574_ (.A1(_04516_),
    .A2(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28575_ (.A1(_04518_),
    .A2(_04515_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28576_ (.A1(_04517_),
    .A2(_04516_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28577_ (.A1(_04514_),
    .A2(_04513_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28578_ (.A1(_04520_),
    .A2(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28579_ (.A1(_04522_),
    .A2(_04519_),
    .A3(_10549_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28580_ (.I(\u0.w[0][1] ),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28581_ (.A1(_11989_),
    .A2(\text_in_r[97] ),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28582_ (.A1(_04524_),
    .A2(_04523_),
    .A3(_04525_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28583_ (.A1(_04520_),
    .A2(_04515_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28584_ (.A1(_04518_),
    .A2(_04521_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28585_ (.A1(_04528_),
    .A2(_04527_),
    .A3(_10549_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28586_ (.A1(_12193_),
    .A2(\text_in_r[97] ),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28587_ (.A1(_04530_),
    .A2(\u0.w[0][1] ),
    .A3(_04529_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28588_ (.A1(_04526_),
    .A2(_04531_),
    .ZN(_16079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28589_ (.A1(_10394_),
    .A2(net679),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28590_ (.A1(_10357_),
    .A2(net574),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28591_ (.A1(_04533_),
    .A2(_04532_),
    .A3(_01557_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28592_ (.A1(_10396_),
    .A2(_10635_),
    .A3(_10395_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28593_ (.A1(_04535_),
    .A2(_04534_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28594_ (.A1(_10342_),
    .A2(_04536_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28595_ (.A1(net1069),
    .A2(_04535_),
    .A3(_10351_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28596_ (.A1(_04538_),
    .A2(_04537_),
    .B(_10410_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28597_ (.I(\text_in_r[96] ),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28598_ (.A1(_04540_),
    .A2(_11202_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28599_ (.A1(_04539_),
    .A2(_04541_),
    .B(\u0.w[0][0] ),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28600_ (.A1(_04537_),
    .A2(_04538_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28601_ (.A1(_04543_),
    .A2(_14333_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28602_ (.I(\u0.w[0][0] ),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28603_ (.I(_04541_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28604_ (.A1(_04544_),
    .A2(_04545_),
    .A3(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28605_ (.A1(_04542_),
    .A2(_04547_),
    .ZN(_16082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28606_ (.A1(net606),
    .A2(\sa20_sr[2] ),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28607_ (.A1(\sa30_sr[1] ),
    .A2(\sa20_sr[2] ),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28608_ (.A1(_04549_),
    .A2(_04548_),
    .B(\sa00_sr[2] ),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28609_ (.A1(_10343_),
    .A2(_10417_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28610_ (.A1(net607),
    .A2(\sa20_sr[2] ),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28611_ (.A1(_04551_),
    .A2(_10450_),
    .A3(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28612_ (.A1(_04550_),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _28613_ (.A1(net619),
    .A2(net860),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28614_ (.I(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28615_ (.A1(_04556_),
    .A2(_04554_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28616_ (.A1(_04555_),
    .A2(_04553_),
    .A3(_04550_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _28617_ (.A1(_04558_),
    .A2(_04557_),
    .B(_10381_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28618_ (.I(\text_in_r[98] ),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28619_ (.A1(_04560_),
    .A2(net595),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28620_ (.I(\u0.w[0][2] ),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _28621_ (.A1(_04559_),
    .A2(_04561_),
    .B(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28622_ (.A1(_04558_),
    .A2(_04557_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28623_ (.A1(_10402_),
    .A2(_04564_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28624_ (.I(_04561_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28625_ (.A1(_04565_),
    .A2(\u0.w[0][2] ),
    .A3(_04566_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28626_ (.A1(_04567_),
    .A2(_04563_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28627_ (.I(_04568_),
    .Z(_16098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28628_ (.A1(_04539_),
    .A2(_04541_),
    .B(_04545_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28629_ (.A1(_04546_),
    .A2(\u0.w[0][0] ),
    .A3(_04544_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28630_ (.A1(_04570_),
    .A2(_04569_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _28631_ (.I(_04571_),
    .Z(_16073_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28632_ (.A1(_04559_),
    .A2(_04561_),
    .B(\u0.w[0][2] ),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28633_ (.A1(_04565_),
    .A2(_04562_),
    .A3(_04566_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28634_ (.A1(_04573_),
    .A2(_04572_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _28635_ (.I(_04574_),
    .Z(_16091_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _28636_ (.I(_04568_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28637_ (.A1(net1075),
    .A2(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28638_ (.A1(_10453_),
    .A2(\sa20_sr[3] ),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28639_ (.A1(_10457_),
    .A2(_10458_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28640_ (.A1(_04577_),
    .A2(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28641_ (.A1(_01634_),
    .A2(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28642_ (.I(_04579_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28643_ (.A1(_01638_),
    .A2(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28644_ (.A1(_04580_),
    .A2(_04582_),
    .A3(_10549_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28645_ (.I(\u0.w[0][3] ),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28646_ (.A1(_11989_),
    .A2(\text_in_r[99] ),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28647_ (.A1(_04583_),
    .A2(_04584_),
    .A3(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28648_ (.A1(_01634_),
    .A2(_04581_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28649_ (.A1(_01638_),
    .A2(_04579_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28650_ (.A1(_04587_),
    .A2(_04588_),
    .A3(_10549_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28651_ (.A1(_12193_),
    .A2(\text_in_r[99] ),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28652_ (.A1(_04589_),
    .A2(\u0.w[0][3] ),
    .A3(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28653_ (.A1(_04586_),
    .A2(_04591_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28654_ (.A1(_04576_),
    .A2(_04592_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28655_ (.A1(_04523_),
    .A2(\u0.w[0][1] ),
    .A3(_04525_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28656_ (.A1(_04529_),
    .A2(_04524_),
    .A3(_04530_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28657_ (.A1(_04594_),
    .A2(_04595_),
    .ZN(_16074_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _28658_ (.A1(net1068),
    .A2(net1065),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28659_ (.A1(_04596_),
    .A2(net1076),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28660_ (.A1(_04593_),
    .A2(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28661_ (.A1(_16074_),
    .A2(net1080),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _28662_ (.I(_04574_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28663_ (.A1(net1074),
    .A2(_16077_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28664_ (.A1(_04599_),
    .A2(_04601_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28665_ (.A1(_04589_),
    .A2(_04584_),
    .A3(_04590_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28666_ (.A1(_04583_),
    .A2(\u0.w[0][3] ),
    .A3(_04585_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28667_ (.A1(_04603_),
    .A2(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28668_ (.I(_04605_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28669_ (.I(_04606_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28670_ (.A1(_04602_),
    .A2(_04607_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28671_ (.A1(_04598_),
    .A2(_04608_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28672_ (.A1(_10515_),
    .A2(_01654_),
    .B(_13010_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28673_ (.A1(_10515_),
    .A2(_01654_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28674_ (.I(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28675_ (.A1(_12115_),
    .A2(\text_in_r[100] ),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28676_ (.A1(_04610_),
    .A2(_04612_),
    .B(_04613_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28677_ (.I(\u0.w[0][4] ),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28678_ (.A1(_04614_),
    .A2(_04615_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28679_ (.A1(_10515_),
    .A2(_01654_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28680_ (.A1(_04617_),
    .A2(_10585_),
    .A3(_04611_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28681_ (.A1(_04618_),
    .A2(\u0.w[0][4] ),
    .A3(_04613_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28682_ (.A1(_04616_),
    .A2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28683_ (.I(_04620_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28684_ (.A1(_04609_),
    .A2(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28685_ (.I(_04592_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28686_ (.I(_04623_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28687_ (.I(_16089_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28688_ (.A1(_04563_),
    .A2(_04625_),
    .A3(_04567_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28689_ (.A1(_04576_),
    .A2(_04624_),
    .A3(_04626_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28690_ (.I(_04620_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28691_ (.A1(_04627_),
    .A2(_04628_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28692_ (.A1(net1143),
    .A2(net74),
    .A3(_04575_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28693_ (.I(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28694_ (.A1(net73),
    .A2(_04600_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28695_ (.I(_04605_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28696_ (.A1(_04632_),
    .A2(_04633_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28697_ (.A1(_04631_),
    .A2(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _28698_ (.A1(\sa30_sr[4] ),
    .A2(\sa20_sr[5] ),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28699_ (.A1(_04636_),
    .A2(\sa00_sr[5] ),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28700_ (.A1(_04636_),
    .A2(\sa00_sr[5] ),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28701_ (.A1(_04637_),
    .A2(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28702_ (.A1(\sa00_sr[4] ),
    .A2(\sa10_sr[5] ),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28703_ (.A1(_04639_),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28704_ (.I(_04640_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28705_ (.A1(_04637_),
    .A2(_04642_),
    .A3(_04638_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28706_ (.A1(_04641_),
    .A2(_04643_),
    .A3(_13010_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28707_ (.A1(_11385_),
    .A2(\text_in_r[101] ),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28708_ (.A1(_04644_),
    .A2(_04645_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28709_ (.I(\u0.w[0][5] ),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28710_ (.A1(_04646_),
    .A2(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28711_ (.A1(_04644_),
    .A2(\u0.w[0][5] ),
    .A3(_04645_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28712_ (.A1(_04648_),
    .A2(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _28713_ (.I(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28714_ (.I(_04651_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28715_ (.A1(_04629_),
    .A2(_04635_),
    .B(_04652_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28716_ (.A1(_04622_),
    .A2(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28717_ (.A1(net1066),
    .A2(_04600_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28718_ (.A1(_04606_),
    .A2(_04655_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28719_ (.A1(_04656_),
    .A2(net1084),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28720_ (.A1(_04657_),
    .A2(_04628_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28721_ (.I(_16076_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28722_ (.A1(_04659_),
    .A2(_04574_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28723_ (.A1(_04660_),
    .A2(_04592_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _28724_ (.I(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28725_ (.A1(_04575_),
    .A2(_04625_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28726_ (.A1(_04662_),
    .A2(_04663_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28727_ (.A1(_04658_),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _28728_ (.I(_16080_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28729_ (.A1(_16091_),
    .A2(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28730_ (.I(_04592_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28731_ (.A1(_04667_),
    .A2(_04668_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28732_ (.A1(_04631_),
    .A2(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28733_ (.A1(_04576_),
    .A2(_04606_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28734_ (.A1(_04614_),
    .A2(\u0.w[0][4] ),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28735_ (.A1(_04618_),
    .A2(_04615_),
    .A3(_04613_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28736_ (.A1(_04672_),
    .A2(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28737_ (.I(_04674_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28738_ (.A1(_04671_),
    .A2(_04675_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28739_ (.I(_04650_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28740_ (.I(_04677_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28741_ (.A1(_04670_),
    .A2(_04676_),
    .B(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28742_ (.A1(_04679_),
    .A2(_04665_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28743_ (.A1(\sa30_sr[5] ),
    .A2(\sa20_sr[6] ),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28744_ (.A1(\sa00_sr[6] ),
    .A2(_04681_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28745_ (.A1(\sa00_sr[5] ),
    .A2(\sa10_sr[6] ),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28746_ (.A1(_04682_),
    .A2(_04683_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28747_ (.A1(_04682_),
    .A2(_04683_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28748_ (.A1(_10587_),
    .A2(\text_in_r[102] ),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _28749_ (.A1(_04684_),
    .A2(_10639_),
    .A3(_04685_),
    .B(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28750_ (.A1(_04687_),
    .A2(\u0.w[0][6] ),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28751_ (.A1(_04687_),
    .A2(\u0.w[0][6] ),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28752_ (.A1(_04688_),
    .A2(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28753_ (.I(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28754_ (.I(_04691_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28755_ (.A1(_04680_),
    .A2(_04654_),
    .B(_04692_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28756_ (.I(_16075_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28757_ (.A1(_16098_),
    .A2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28758_ (.I(_16083_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28759_ (.A1(_16091_),
    .A2(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28760_ (.A1(_04695_),
    .A2(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28761_ (.A1(_04698_),
    .A2(_04624_),
    .B(_04620_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28762_ (.A1(_04596_),
    .A2(_16098_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28763_ (.A1(_04660_),
    .A2(_04606_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28764_ (.A1(_04700_),
    .A2(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28765_ (.A1(_04702_),
    .A2(_04699_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28766_ (.A1(net73),
    .A2(net74),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28767_ (.A1(_04600_),
    .A2(_16082_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28768_ (.A1(_04704_),
    .A2(_04705_),
    .A3(_04607_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28769_ (.A1(net1143),
    .A2(net1065),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28770_ (.A1(_16082_),
    .A2(_04575_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28771_ (.A1(_04707_),
    .A2(_04668_),
    .A3(_04708_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28772_ (.A1(_04706_),
    .A2(_04709_),
    .A3(_04628_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28773_ (.A1(_04710_),
    .A2(_04703_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28774_ (.I(_04677_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28775_ (.A1(_04712_),
    .A2(_04711_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28776_ (.A1(_16098_),
    .A2(_16075_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28777_ (.A1(_04660_),
    .A2(_04714_),
    .A3(_04624_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28778_ (.A1(_16091_),
    .A2(_16075_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28779_ (.A1(_04575_),
    .A2(_16083_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28780_ (.A1(_04716_),
    .A2(_04717_),
    .A3(_04607_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28781_ (.A1(_04715_),
    .A2(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28782_ (.I(_04674_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28783_ (.A1(_04719_),
    .A2(_04720_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28784_ (.I(_04651_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28785_ (.A1(net1143),
    .A2(_04575_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28786_ (.A1(net578),
    .A2(_04600_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28787_ (.I(_04606_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28788_ (.A1(_04723_),
    .A2(_04724_),
    .A3(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28789_ (.I(_04620_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28790_ (.A1(_04659_),
    .A2(_04575_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28791_ (.A1(_04728_),
    .A2(_04592_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28792_ (.A1(_04726_),
    .A2(_04727_),
    .A3(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28793_ (.A1(_04721_),
    .A2(_04722_),
    .A3(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28794_ (.I(_04690_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28795_ (.A1(_04732_),
    .A2(_04731_),
    .A3(_04713_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28796_ (.A1(_04733_),
    .A2(_04693_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28797_ (.A1(\sa30_sr[6] ),
    .A2(_10389_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _28798_ (.A1(_13742_),
    .A2(net47),
    .A3(_04735_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28799_ (.A1(_12961_),
    .A2(\text_in_r[103] ),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28800_ (.A1(_04736_),
    .A2(_12965_),
    .B(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28801_ (.A1(\u0.w[0][7] ),
    .A2(_04738_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28802_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28803_ (.A1(_04740_),
    .A2(_04734_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28804_ (.A1(_16098_),
    .A2(_16080_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28805_ (.A1(_04742_),
    .A2(_04668_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28806_ (.A1(_04743_),
    .A2(_04675_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28807_ (.A1(_04744_),
    .A2(_04598_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28808_ (.A1(net1074),
    .A2(_16085_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28809_ (.A1(_04742_),
    .A2(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28810_ (.A1(_04747_),
    .A2(_04607_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28811_ (.A1(_04748_),
    .A2(_04621_),
    .A3(_04661_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28812_ (.I(_04651_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28813_ (.A1(_04745_),
    .A2(_04749_),
    .A3(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28814_ (.A1(net1142),
    .A2(net1074),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28815_ (.A1(_04575_),
    .A2(net578),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28816_ (.A1(_04752_),
    .A2(_04753_),
    .A3(_04633_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28817_ (.A1(_04754_),
    .A2(_04675_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28818_ (.A1(_04655_),
    .A2(_04717_),
    .A3(_04624_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28819_ (.A1(_04755_),
    .A2(_04756_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28820_ (.I(_04620_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28821_ (.A1(_04669_),
    .A2(_04758_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28822_ (.A1(_04695_),
    .A2(_04601_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28823_ (.I(_04633_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28824_ (.A1(_04760_),
    .A2(_04761_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28825_ (.A1(_04759_),
    .A2(_04762_),
    .B(_04652_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28826_ (.A1(_04757_),
    .A2(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28827_ (.A1(_04751_),
    .A2(_04764_),
    .B(_04732_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28828_ (.I(_16085_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28829_ (.A1(_04766_),
    .A2(_04575_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28830_ (.A1(_04767_),
    .A2(_04623_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28831_ (.A1(net22),
    .A2(_04600_),
    .A3(net74),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28832_ (.A1(_04768_),
    .A2(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _28833_ (.I(_04601_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28834_ (.A1(_04771_),
    .A2(_04761_),
    .B(_04628_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28835_ (.A1(_04770_),
    .A2(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28836_ (.A1(_04717_),
    .A2(_04606_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28837_ (.I(_04774_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28838_ (.A1(_04775_),
    .A2(_04769_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28839_ (.A1(_04771_),
    .A2(_04624_),
    .B(_04674_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28840_ (.A1(_04776_),
    .A2(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28841_ (.I(_04677_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28842_ (.A1(_04773_),
    .A2(_04778_),
    .A3(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28843_ (.A1(_04575_),
    .A2(_04666_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28844_ (.A1(_04769_),
    .A2(_04607_),
    .A3(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28845_ (.A1(_04593_),
    .A2(_04716_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28846_ (.A1(_16098_),
    .A2(_16077_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28847_ (.I(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28848_ (.A1(_04785_),
    .A2(_04725_),
    .B(_04758_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28849_ (.A1(_04782_),
    .A2(_04783_),
    .A3(_04786_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28850_ (.A1(_04607_),
    .A2(_16096_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28851_ (.A1(_04753_),
    .A2(_04606_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28852_ (.A1(_04788_),
    .A2(_04789_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28853_ (.A1(_04790_),
    .A2(_04621_),
    .B(_04678_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28854_ (.A1(_04787_),
    .A2(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28855_ (.A1(_04780_),
    .A2(_04792_),
    .B(_04692_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _28856_ (.I(_04739_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28857_ (.A1(_04765_),
    .A2(_04793_),
    .B(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28858_ (.A1(_04795_),
    .A2(_04741_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28859_ (.A1(_04708_),
    .A2(_04633_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28860_ (.A1(net1074),
    .A2(_04694_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28861_ (.A1(_04796_),
    .A2(_04797_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28862_ (.A1(net1083),
    .A2(_04742_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28863_ (.A1(_04798_),
    .A2(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28864_ (.I(_04758_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28865_ (.A1(_04800_),
    .A2(_04801_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28866_ (.I(_04789_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28867_ (.A1(_04803_),
    .A2(_04655_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28868_ (.A1(net22),
    .A2(_16082_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28869_ (.A1(_04805_),
    .A2(_04655_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28870_ (.I(_04624_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28871_ (.A1(_04806_),
    .A2(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28872_ (.I(_04675_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28873_ (.A1(_04804_),
    .A2(_04808_),
    .A3(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28874_ (.A1(_04802_),
    .A2(_04810_),
    .A3(_04750_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _28875_ (.I(_04623_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28876_ (.A1(_04700_),
    .A2(_04812_),
    .A3(_04724_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28877_ (.A1(_04607_),
    .A2(_16080_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28878_ (.A1(_04814_),
    .A2(net1076),
    .B(_04727_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28879_ (.A1(_04813_),
    .A2(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28880_ (.A1(_04632_),
    .A2(net579),
    .A3(_04668_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28881_ (.A1(_04805_),
    .A2(net1076),
    .A3(_04761_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28882_ (.I(_04758_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28883_ (.A1(_04817_),
    .A2(_04818_),
    .A3(_04819_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28884_ (.A1(_04816_),
    .A2(_04820_),
    .A3(_04779_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28885_ (.A1(_04811_),
    .A2(_04821_),
    .A3(_04692_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28886_ (.A1(_04752_),
    .A2(_04606_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28887_ (.A1(_04823_),
    .A2(_04704_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28888_ (.A1(_04623_),
    .A2(_16098_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28889_ (.A1(_04825_),
    .A2(_04707_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28890_ (.A1(_04824_),
    .A2(_04809_),
    .A3(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28891_ (.A1(_04593_),
    .A2(_04660_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28892_ (.A1(_04708_),
    .A2(_04667_),
    .A3(_04761_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28893_ (.A1(_04828_),
    .A2(_04819_),
    .A3(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28894_ (.A1(_04827_),
    .A2(_04830_),
    .A3(_04779_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28895_ (.A1(_04743_),
    .A2(_04758_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28896_ (.A1(_04723_),
    .A2(_04623_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28897_ (.A1(_04833_),
    .A2(_04632_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28898_ (.A1(_04832_),
    .A2(_04834_),
    .B(_04712_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28899_ (.I(_04729_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28900_ (.A1(_04836_),
    .A2(_04626_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28901_ (.A1(_04782_),
    .A2(_04837_),
    .A3(_04809_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28902_ (.A1(_04835_),
    .A2(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28903_ (.A1(_04831_),
    .A2(_04839_),
    .A3(_04732_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28904_ (.A1(_04822_),
    .A2(_04840_),
    .A3(_04794_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28905_ (.A1(_04708_),
    .A2(_04601_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28906_ (.I(_04633_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28907_ (.A1(_04842_),
    .A2(_04843_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28908_ (.A1(_04716_),
    .A2(_04728_),
    .A3(_04812_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28909_ (.A1(_04844_),
    .A2(_04845_),
    .A3(_04819_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28910_ (.A1(_04599_),
    .A2(_04667_),
    .A3(_04812_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28911_ (.A1(_04705_),
    .A2(_04714_),
    .A3(_04761_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28912_ (.I(_04674_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28913_ (.A1(_04847_),
    .A2(_04848_),
    .A3(_04849_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28914_ (.A1(_04846_),
    .A2(_04850_),
    .A3(_04779_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _28915_ (.I(_04671_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28916_ (.A1(_04852_),
    .A2(_04597_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28917_ (.A1(_04661_),
    .A2(_04675_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28918_ (.A1(_04853_),
    .A2(_04854_),
    .B(_04678_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28919_ (.A1(_04626_),
    .A2(_04633_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28920_ (.I(_16077_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28921_ (.A1(_16098_),
    .A2(_04857_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28922_ (.A1(_04856_),
    .A2(_04858_),
    .B(_04675_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28923_ (.A1(_04813_),
    .A2(_04859_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28924_ (.A1(_04855_),
    .A2(_04860_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28925_ (.A1(_04861_),
    .A2(_04851_),
    .B(_04732_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28926_ (.A1(_04623_),
    .A2(net1076),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28927_ (.A1(_04863_),
    .A2(net74),
    .B(_04652_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28928_ (.A1(_04707_),
    .A2(_04752_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28929_ (.A1(_04865_),
    .A2(_04812_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28930_ (.A1(_04656_),
    .A2(_04714_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28931_ (.A1(_04864_),
    .A2(_04866_),
    .A3(_04867_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28932_ (.A1(_04705_),
    .A2(_04606_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28933_ (.I(_04869_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28934_ (.A1(_04870_),
    .A2(_04723_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28935_ (.A1(_04871_),
    .A2(_04722_),
    .A3(_04847_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28936_ (.A1(_04868_),
    .A2(_04872_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _28937_ (.A1(_04677_),
    .A2(_16099_),
    .A3(_04725_),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28938_ (.A1(_04597_),
    .A2(_04775_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28939_ (.A1(_04874_),
    .A2(_04875_),
    .A3(_04720_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28940_ (.I(_04690_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28941_ (.A1(_04876_),
    .A2(_04877_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28942_ (.A1(_04873_),
    .A2(_04801_),
    .B(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28943_ (.A1(_04862_),
    .A2(_04879_),
    .B(_04740_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28944_ (.A1(_04841_),
    .A2(_04880_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28945_ (.A1(_04781_),
    .A2(_04623_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28946_ (.A1(_04881_),
    .A2(_04632_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28947_ (.A1(_04882_),
    .A2(_04675_),
    .A3(_04748_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28948_ (.A1(_04746_),
    .A2(_04668_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28949_ (.A1(_04884_),
    .A2(_04674_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28950_ (.A1(net1070),
    .A2(_04781_),
    .A3(_04624_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28951_ (.A1(_16098_),
    .A2(_16089_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28952_ (.A1(_04887_),
    .A2(_04607_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28953_ (.A1(_04885_),
    .A2(_04886_),
    .A3(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28954_ (.A1(_04883_),
    .A2(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28955_ (.A1(_04890_),
    .A2(_04750_),
    .B(_04877_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28956_ (.A1(_04656_),
    .A2(net1072),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28957_ (.A1(net1083),
    .A2(_04753_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28958_ (.A1(_04892_),
    .A2(_04893_),
    .A3(_04677_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28959_ (.A1(_04677_),
    .A2(_04620_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28960_ (.A1(_04599_),
    .A2(_04623_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28961_ (.A1(_04896_),
    .A2(_04746_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28962_ (.A1(_04869_),
    .A2(_04887_),
    .B(_04620_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28963_ (.A1(_04897_),
    .A2(_04898_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28964_ (.A1(_04894_),
    .A2(_04895_),
    .B(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28965_ (.A1(_04891_),
    .A2(_04900_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28966_ (.A1(_04724_),
    .A2(_04606_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28967_ (.A1(_04902_),
    .A2(_04599_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28968_ (.A1(_04705_),
    .A2(_04784_),
    .A3(_04812_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28969_ (.A1(_04903_),
    .A2(_04904_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28970_ (.A1(_04905_),
    .A2(_04809_),
    .B(_04712_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _28971_ (.I(_04668_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28972_ (.A1(_04700_),
    .A2(_04907_),
    .A3(_04626_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28973_ (.A1(_04630_),
    .A2(_04607_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28974_ (.A1(_04908_),
    .A2(_04909_),
    .B(_04621_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28975_ (.A1(_04906_),
    .A2(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28976_ (.A1(_04865_),
    .A2(_04727_),
    .A3(_04907_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28977_ (.A1(_04620_),
    .A2(net579),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28978_ (.A1(_04667_),
    .A2(_04633_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28979_ (.A1(_04913_),
    .A2(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28980_ (.A1(_04915_),
    .A2(_04678_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28981_ (.A1(_04912_),
    .A2(_04916_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28982_ (.A1(_04769_),
    .A2(_04781_),
    .B(_04725_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28983_ (.A1(_04755_),
    .A2(_04918_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28984_ (.A1(_04917_),
    .A2(_04919_),
    .B(_04732_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28985_ (.A1(_04911_),
    .A2(_04920_),
    .B(_04740_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28986_ (.A1(_04901_),
    .A2(_04921_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28987_ (.A1(_16103_),
    .A2(_04843_),
    .B(_04677_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28988_ (.A1(_04866_),
    .A2(_04923_),
    .B(_04849_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28989_ (.A1(_04857_),
    .A2(_04666_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28990_ (.I(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28991_ (.A1(_04863_),
    .A2(_04926_),
    .B(_04652_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28992_ (.A1(_04599_),
    .A2(_04576_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28993_ (.A1(_04928_),
    .A2(_04907_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28994_ (.A1(_04927_),
    .A2(_04875_),
    .A3(_04929_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28995_ (.A1(_04924_),
    .A2(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28996_ (.A1(_04843_),
    .A2(_04797_),
    .B(_04651_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28997_ (.A1(net1083),
    .A2(_04781_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28998_ (.A1(_04932_),
    .A2(_04933_),
    .B(_04621_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28999_ (.A1(_04633_),
    .A2(_16094_),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29000_ (.A1(_04909_),
    .A2(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29001_ (.A1(_04936_),
    .A2(_04678_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29002_ (.A1(_04934_),
    .A2(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29003_ (.A1(_04931_),
    .A2(_04938_),
    .A3(_04732_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29004_ (.A1(_04896_),
    .A2(net1070),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29005_ (.A1(_04940_),
    .A2(_04819_),
    .A3(_04754_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29006_ (.A1(_04836_),
    .A2(_04769_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29007_ (.A1(_16096_),
    .A2(_04761_),
    .B(_04628_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29008_ (.A1(_04942_),
    .A2(_04943_),
    .B(_04722_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29009_ (.A1(_04941_),
    .A2(_04944_),
    .B(_04877_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29010_ (.A1(_04823_),
    .A2(_04695_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29011_ (.A1(_04753_),
    .A2(_04697_),
    .A3(_04812_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29012_ (.A1(_04946_),
    .A2(_04947_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29013_ (.A1(_04948_),
    .A2(_04801_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29014_ (.A1(_04704_),
    .A2(_04752_),
    .A3(_04668_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29015_ (.A1(_04812_),
    .A2(_16099_),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29016_ (.A1(_04950_),
    .A2(_04849_),
    .A3(_04951_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29017_ (.A1(_04949_),
    .A2(_04952_),
    .A3(_04750_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29018_ (.A1(_04945_),
    .A2(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29019_ (.A1(_04939_),
    .A2(_04954_),
    .B(_04740_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29020_ (.A1(_04922_),
    .A2(_04955_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29021_ (.A1(_04881_),
    .A2(_04626_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29022_ (.A1(_04677_),
    .A2(_04674_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29023_ (.A1(_04903_),
    .A2(_04956_),
    .A3(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29024_ (.A1(_04958_),
    .A2(_04690_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29025_ (.I(_04797_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29026_ (.A1(_04836_),
    .A2(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29027_ (.A1(_04708_),
    .A2(_04633_),
    .A3(_04697_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29028_ (.A1(_04961_),
    .A2(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29029_ (.A1(_04963_),
    .A2(_04895_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29030_ (.A1(_04959_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29031_ (.A1(_04704_),
    .A2(_04708_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29032_ (.A1(_04966_),
    .A2(_04725_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29033_ (.A1(_04599_),
    .A2(_04660_),
    .A3(_04624_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29034_ (.A1(_04967_),
    .A2(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29035_ (.A1(_04969_),
    .A2(_04720_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29036_ (.I(_04728_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29037_ (.A1(_04971_),
    .A2(_04668_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29038_ (.I(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29039_ (.A1(_04871_),
    .A2(_04973_),
    .A3(_04727_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29040_ (.A1(_04970_),
    .A2(_04974_),
    .A3(_04750_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29041_ (.A1(_04965_),
    .A2(_04975_),
    .B(_04740_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _29042_ (.A1(_04599_),
    .A2(_04708_),
    .A3(_04697_),
    .A4(_04812_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29043_ (.A1(_04805_),
    .A2(net1076),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29044_ (.A1(_04803_),
    .A2(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29045_ (.A1(_04979_),
    .A2(_04720_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29046_ (.A1(_16098_),
    .A2(_04696_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29047_ (.I(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29048_ (.A1(_04701_),
    .A2(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29049_ (.A1(_04983_),
    .A2(_04727_),
    .A3(_04709_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29050_ (.A1(_04977_),
    .A2(_04980_),
    .B(_04984_),
    .C(_04712_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29051_ (.A1(_04902_),
    .A2(_04767_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29052_ (.A1(_04986_),
    .A2(_04628_),
    .A3(_04817_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _29053_ (.A1(_04966_),
    .A2(_04620_),
    .A3(_04863_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29054_ (.A1(_04987_),
    .A2(_04988_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29055_ (.A1(_04989_),
    .A2(_04750_),
    .B(_04877_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29056_ (.A1(_04985_),
    .A2(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29057_ (.A1(_04976_),
    .A2(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29058_ (.A1(_04925_),
    .A2(net1074),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29059_ (.A1(_04993_),
    .A2(_04623_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29060_ (.A1(_04994_),
    .A2(net1071),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29061_ (.A1(_04875_),
    .A2(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29062_ (.A1(_04996_),
    .A2(_04720_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29063_ (.A1(_04898_),
    .A2(_04652_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29064_ (.A1(_04997_),
    .A2(_04998_),
    .B(_04877_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29065_ (.A1(_04824_),
    .A2(_04783_),
    .A3(_04675_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29066_ (.A1(_04701_),
    .A2(_04663_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29067_ (.I(_04746_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29068_ (.A1(_05002_),
    .A2(_04624_),
    .B(_04674_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29069_ (.A1(_04825_),
    .A2(net74),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29070_ (.A1(_05001_),
    .A2(_05003_),
    .A3(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29071_ (.A1(_05000_),
    .A2(_05005_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29072_ (.A1(_05006_),
    .A2(_04779_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29073_ (.A1(_04999_),
    .A2(_05007_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29074_ (.A1(_04852_),
    .A2(_04660_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29075_ (.A1(_04994_),
    .A2(_04663_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29076_ (.A1(_05009_),
    .A2(_05010_),
    .A3(_04652_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29077_ (.A1(_05002_),
    .A2(_04668_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29078_ (.A1(_04892_),
    .A2(_04677_),
    .A3(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29079_ (.A1(_05011_),
    .A2(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29080_ (.A1(_05014_),
    .A2(_04809_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29081_ (.I(_04752_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29082_ (.A1(_04774_),
    .A2(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29083_ (.A1(_05017_),
    .A2(_04972_),
    .B(_04652_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29084_ (.I(_04777_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29085_ (.A1(_04660_),
    .A2(_04623_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29086_ (.A1(_05020_),
    .A2(_04651_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29087_ (.A1(_05019_),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29088_ (.A1(_05018_),
    .A2(_05022_),
    .B(_04691_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29089_ (.A1(_05015_),
    .A2(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29090_ (.A1(_05008_),
    .A2(_05024_),
    .A3(_04740_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29091_ (.A1(_04992_),
    .A2(_05025_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29092_ (.A1(_04871_),
    .A2(_04950_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29093_ (.A1(_05026_),
    .A2(_04720_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29094_ (.A1(_04599_),
    .A2(_04707_),
    .A3(_04725_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29095_ (.A1(_04752_),
    .A2(_04695_),
    .A3(_04812_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29096_ (.A1(_05028_),
    .A2(_05029_),
    .A3(_04621_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29097_ (.A1(_05027_),
    .A2(_04691_),
    .A3(_05030_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29098_ (.A1(_04769_),
    .A2(_04758_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29099_ (.A1(_04674_),
    .A2(_04716_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29100_ (.A1(_05032_),
    .A2(_05033_),
    .B(_04896_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29101_ (.A1(_04782_),
    .A2(_04727_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29102_ (.A1(_04915_),
    .A2(_04691_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29103_ (.A1(_05034_),
    .A2(_05035_),
    .A3(_05036_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29104_ (.A1(_05031_),
    .A2(_05037_),
    .B(_04750_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29105_ (.A1(_04768_),
    .A2(_04720_),
    .A3(_04771_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29106_ (.A1(_05039_),
    .A2(_04877_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29107_ (.I(_04833_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29108_ (.A1(_05041_),
    .A2(_04655_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29109_ (.A1(_05042_),
    .A2(_04867_),
    .A3(_04849_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29110_ (.A1(_05040_),
    .A2(_05043_),
    .B(_04750_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29111_ (.A1(_04856_),
    .A2(_04728_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29112_ (.A1(_04770_),
    .A2(_05045_),
    .A3(_04809_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29113_ (.I(_04753_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29114_ (.A1(_05047_),
    .A2(_04668_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29115_ (.A1(_05003_),
    .A2(_04748_),
    .A3(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29116_ (.A1(_05046_),
    .A2(_05049_),
    .A3(_04732_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29117_ (.A1(_05044_),
    .A2(_05050_),
    .B(_04740_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29118_ (.A1(_05038_),
    .A2(_05051_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29119_ (.I(_16087_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29120_ (.A1(_05053_),
    .A2(_04807_),
    .B(_05048_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29121_ (.A1(_05054_),
    .A2(_04712_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29122_ (.A1(_04762_),
    .A2(_04709_),
    .A3(_04722_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29123_ (.A1(_05055_),
    .A2(_04809_),
    .A3(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29124_ (.A1(_04768_),
    .A2(_04705_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29125_ (.A1(_05058_),
    .A2(_05028_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29126_ (.A1(_04651_),
    .A2(_04620_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29127_ (.A1(_05059_),
    .A2(_05060_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29128_ (.A1(_04768_),
    .A2(_04632_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29129_ (.A1(_04707_),
    .A2(net1076),
    .A3(_04761_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29130_ (.A1(_05062_),
    .A2(_05063_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29131_ (.A1(_05064_),
    .A2(_04895_),
    .B(_04691_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29132_ (.A1(_05057_),
    .A2(_05061_),
    .A3(_05065_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29133_ (.A1(_04700_),
    .A2(_04807_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29134_ (.A1(_04858_),
    .A2(_04633_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29135_ (.A1(_05068_),
    .A2(_04628_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29136_ (.A1(_05067_),
    .A2(_05069_),
    .B(_04722_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29137_ (.A1(_04914_),
    .A2(_05047_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29138_ (.A1(_04598_),
    .A2(_05071_),
    .A3(_04849_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29139_ (.A1(_05070_),
    .A2(_05072_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29140_ (.A1(_04870_),
    .A2(_04663_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29141_ (.A1(_04825_),
    .A2(_04727_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29142_ (.A1(_05074_),
    .A2(_05075_),
    .B(_04712_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29143_ (.A1(_04723_),
    .A2(_04607_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29144_ (.A1(_05077_),
    .A2(_04716_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29145_ (.A1(_05078_),
    .A2(_04819_),
    .A3(_04847_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29146_ (.A1(_05076_),
    .A2(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29147_ (.A1(_05073_),
    .A2(_05080_),
    .A3(_04692_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29148_ (.A1(_05066_),
    .A2(_05081_),
    .A3(_04740_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29149_ (.A1(_05052_),
    .A2(_05082_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29150_ (.A1(_04826_),
    .A2(_04628_),
    .A3(_04914_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29151_ (.A1(_04576_),
    .A2(_04746_),
    .B(_04725_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29152_ (.A1(_05084_),
    .A2(_04727_),
    .A3(_04701_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _29153_ (.A1(_05083_),
    .A2(_05085_),
    .A3(_04877_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29154_ (.A1(_05048_),
    .A2(_04628_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29155_ (.I(_05068_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29156_ (.A1(_05088_),
    .A2(_04752_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29157_ (.A1(_05087_),
    .A2(_05089_),
    .B(_04691_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29158_ (.A1(_04660_),
    .A2(_04695_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29159_ (.A1(_04843_),
    .A2(_05091_),
    .B(_04888_),
    .C(_04720_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29160_ (.A1(_05090_),
    .A2(_05092_),
    .B(_04779_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29161_ (.A1(_05086_),
    .A2(_05093_),
    .B(_04740_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29162_ (.A1(_04597_),
    .A2(_04717_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29163_ (.A1(_04671_),
    .A2(_04596_),
    .B(_04727_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29164_ (.A1(_05095_),
    .A2(_04807_),
    .B(_05096_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29165_ (.A1(_04812_),
    .A2(net73),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29166_ (.A1(_05028_),
    .A2(_04720_),
    .A3(_05098_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29167_ (.A1(_05099_),
    .A2(_04877_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29168_ (.A1(_05097_),
    .A2(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29169_ (.A1(_04769_),
    .A2(_04843_),
    .A3(net1071),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29170_ (.A1(_04881_),
    .A2(_04926_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29171_ (.A1(_05102_),
    .A2(_05103_),
    .A3(_04819_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29172_ (.I(_04663_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29173_ (.A1(_04669_),
    .A2(_05105_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29174_ (.A1(_05106_),
    .A2(_04608_),
    .A3(_04849_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29175_ (.A1(_05104_),
    .A2(_05107_),
    .B(_04732_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29176_ (.A1(_05101_),
    .A2(_05108_),
    .B(_04779_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29177_ (.A1(_05094_),
    .A2(_05109_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29178_ (.A1(_04724_),
    .A2(_04663_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29179_ (.A1(_05111_),
    .A2(_04725_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29180_ (.A1(_04662_),
    .A2(_04717_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29181_ (.A1(_05113_),
    .A2(_05112_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29182_ (.A1(_05060_),
    .A2(_05114_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29183_ (.A1(_04877_),
    .A2(_05115_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29184_ (.A1(_04597_),
    .A2(_04761_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29185_ (.A1(_04907_),
    .A2(_04696_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _29186_ (.A1(_05117_),
    .A2(_05118_),
    .B(_04678_),
    .C(_04621_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29187_ (.A1(_05119_),
    .A2(_05116_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29188_ (.I(_04994_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29189_ (.A1(_05117_),
    .A2(_04631_),
    .B(_04849_),
    .C(_05121_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29190_ (.A1(_04663_),
    .A2(_04807_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29191_ (.A1(_04832_),
    .A2(_05123_),
    .B(_04722_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29192_ (.A1(_05122_),
    .A2(_05124_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29193_ (.A1(_05120_),
    .A2(_05125_),
    .B(_04794_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29194_ (.A1(net1077),
    .A2(_04781_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _29195_ (.A1(_04722_),
    .A2(_04598_),
    .A3(_05127_),
    .A4(_04849_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29196_ (.A1(_04981_),
    .A2(_04907_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29197_ (.A1(_05117_),
    .A2(_05105_),
    .B(_05060_),
    .C(_05129_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29198_ (.A1(_05128_),
    .A2(_05130_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29199_ (.I(_04634_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29200_ (.A1(_05132_),
    .A2(net1071),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29201_ (.A1(_04662_),
    .A2(_04630_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29202_ (.A1(_05133_),
    .A2(_05134_),
    .A3(_04819_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29203_ (.A1(_04907_),
    .A2(_16082_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29204_ (.A1(_04706_),
    .A2(_04849_),
    .A3(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29205_ (.A1(_05135_),
    .A2(_05137_),
    .B(_04750_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29206_ (.A1(_05131_),
    .A2(_05138_),
    .B(_04692_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29207_ (.A1(_05139_),
    .A2(_05126_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29208_ (.A1(_05140_),
    .A2(_05110_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29209_ (.A1(_05004_),
    .A2(_04675_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29210_ (.A1(_04803_),
    .A2(_04993_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29211_ (.A1(_05141_),
    .A2(_04709_),
    .A3(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29212_ (.A1(_05041_),
    .A2(_04707_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29213_ (.A1(_04981_),
    .A2(_04843_),
    .B(_04675_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29214_ (.A1(_05144_),
    .A2(_05145_),
    .B(_04712_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29215_ (.A1(_05143_),
    .A2(_05146_),
    .B(_04692_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29216_ (.A1(_04630_),
    .A2(_04907_),
    .A3(_04632_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29217_ (.A1(_05088_),
    .A2(_04724_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29218_ (.A1(_05148_),
    .A2(_05149_),
    .B(_04819_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29219_ (.A1(_05020_),
    .A2(_04758_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29220_ (.A1(_04936_),
    .A2(_05151_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29221_ (.A1(_05150_),
    .A2(_05152_),
    .B(_04779_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29222_ (.A1(_05147_),
    .A2(_05153_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29223_ (.A1(_04797_),
    .A2(_04725_),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29224_ (.I(_05012_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29225_ (.A1(_05155_),
    .A2(_05156_),
    .B(_04678_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29226_ (.A1(_04785_),
    .A2(_04807_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29227_ (.A1(_05157_),
    .A2(_05158_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29228_ (.A1(_05159_),
    .A2(_04801_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29229_ (.A1(_16092_),
    .A2(_16101_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29230_ (.A1(_04843_),
    .A2(_05161_),
    .B(_04652_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29231_ (.A1(_04896_),
    .A2(_04707_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29232_ (.A1(_05162_),
    .A2(_05163_),
    .B(_04819_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29233_ (.A1(_04771_),
    .A2(_04907_),
    .B(_04677_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29234_ (.A1(_04856_),
    .A2(net1072),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29235_ (.A1(_05165_),
    .A2(_04929_),
    .A3(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29236_ (.A1(_05164_),
    .A2(_05167_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29237_ (.A1(_04803_),
    .A2(_04705_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29238_ (.A1(_04747_),
    .A2(_04807_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29239_ (.A1(_05169_),
    .A2(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29240_ (.A1(_05171_),
    .A2(_05060_),
    .B(_04877_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29241_ (.A1(_05160_),
    .A2(_05168_),
    .A3(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29242_ (.A1(_05154_),
    .A2(_05173_),
    .A3(_04794_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29243_ (.A1(_04807_),
    .A2(net1144),
    .B(_05004_),
    .C(_05012_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29244_ (.A1(_04833_),
    .A2(_04758_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29245_ (.A1(_05176_),
    .A2(_04657_),
    .B(_04678_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29246_ (.A1(_05175_),
    .A2(_04801_),
    .B(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29247_ (.A1(_04966_),
    .A2(_04725_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29248_ (.A1(_05179_),
    .A2(_04865_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29249_ (.A1(_05180_),
    .A2(_04809_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29250_ (.A1(_04856_),
    .A2(_04708_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29251_ (.A1(_05179_),
    .A2(_04801_),
    .A3(_05182_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29252_ (.A1(_05181_),
    .A2(_05183_),
    .A3(_04779_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29253_ (.A1(_05178_),
    .A2(_05184_),
    .A3(_04692_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29254_ (.A1(_04774_),
    .A2(_04758_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29255_ (.A1(_05062_),
    .A2(_05186_),
    .B(_04678_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29256_ (.A1(_04918_),
    .A2(_04809_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29257_ (.A1(_05187_),
    .A2(_05188_),
    .B(_04692_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29258_ (.I(_16093_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29259_ (.A1(_05190_),
    .A2(_04907_),
    .B(_04628_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29260_ (.A1(_05133_),
    .A2(_05191_),
    .B(_04722_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29261_ (.A1(_05111_),
    .A2(_04843_),
    .B(_04796_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29262_ (.A1(_05193_),
    .A2(_04801_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29263_ (.A1(_05192_),
    .A2(_05194_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29264_ (.A1(_05189_),
    .A2(_05195_),
    .B(_04794_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29265_ (.A1(_05185_),
    .A2(_05196_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29266_ (.A1(_05174_),
    .A2(_05197_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29267_ (.A1(_04700_),
    .A2(_04807_),
    .A3(_04716_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29268_ (.A1(_04852_),
    .A2(_04769_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29269_ (.A1(_05198_),
    .A2(_05199_),
    .A3(_04712_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29270_ (.A1(_05009_),
    .A2(_04837_),
    .A3(_04722_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29271_ (.A1(_05200_),
    .A2(_04801_),
    .A3(_05201_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29272_ (.A1(_04940_),
    .A2(_05166_),
    .A3(_04722_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29273_ (.A1(_04856_),
    .A2(_04652_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29274_ (.A1(_05062_),
    .A2(_05204_),
    .B(_04621_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29275_ (.A1(_05203_),
    .A2(_05205_),
    .B(_04732_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29276_ (.A1(_05202_),
    .A2(_05206_),
    .B(_04794_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29277_ (.A1(_04761_),
    .A2(net74),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29278_ (.A1(_05042_),
    .A2(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29279_ (.A1(_05209_),
    .A2(_04801_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29280_ (.A1(_05132_),
    .A2(_04700_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29281_ (.A1(_05211_),
    .A2(_04809_),
    .A3(_04950_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29282_ (.A1(_05210_),
    .A2(_05212_),
    .A3(_04779_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29283_ (.A1(_04843_),
    .A2(_04978_),
    .B(_05020_),
    .C(_04849_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29284_ (.A1(_04769_),
    .A2(_04807_),
    .B(_04720_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29285_ (.A1(_04700_),
    .A2(_04902_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29286_ (.A1(_05215_),
    .A2(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29287_ (.A1(_05214_),
    .A2(_04750_),
    .A3(_05217_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29288_ (.A1(_05213_),
    .A2(_05218_),
    .A3(_04732_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29289_ (.A1(_05207_),
    .A2(_05219_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _29290_ (.A1(_04852_),
    .A2(_04632_),
    .B1(_04836_),
    .B2(_04724_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29291_ (.A1(_05221_),
    .A2(_04801_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29292_ (.A1(_04624_),
    .A2(_16101_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29293_ (.A1(_04884_),
    .A2(_05223_),
    .A3(_04727_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29294_ (.A1(_04971_),
    .A2(_04843_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29295_ (.A1(_05224_),
    .A2(_05225_),
    .B(_04712_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29296_ (.A1(_05222_),
    .A2(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29297_ (.A1(_05077_),
    .A2(_04707_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29298_ (.A1(_05228_),
    .A2(_04819_),
    .A3(_04847_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29299_ (.A1(_04907_),
    .A2(_05053_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29300_ (.A1(_04786_),
    .A2(_05230_),
    .B(_04652_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29301_ (.A1(_05229_),
    .A2(_05231_),
    .B(_04692_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29302_ (.A1(_05227_),
    .A2(_05232_),
    .B(_04740_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29303_ (.A1(_04823_),
    .A2(_04805_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29304_ (.A1(_05234_),
    .A2(_04995_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29305_ (.A1(_05235_),
    .A2(_04621_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29306_ (.A1(_04700_),
    .A2(_04716_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29307_ (.A1(_05237_),
    .A2(_04761_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29308_ (.A1(_04662_),
    .A2(_04982_),
    .B(_04758_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29309_ (.A1(_05239_),
    .A2(_05238_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29310_ (.A1(_05236_),
    .A2(_05240_),
    .A3(_04712_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29311_ (.I(_05163_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29312_ (.A1(_05242_),
    .A2(_04814_),
    .B(_04621_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29313_ (.A1(_04833_),
    .A2(_05068_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29314_ (.A1(_05244_),
    .A2(_05033_),
    .B(_04678_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29315_ (.A1(_05243_),
    .A2(_05245_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29316_ (.A1(_05241_),
    .A2(_05246_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29317_ (.A1(_05247_),
    .A2(_04692_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29318_ (.A1(_05233_),
    .A2(_05248_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29319_ (.A1(_05220_),
    .A2(_05249_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29320_ (.A1(_02288_),
    .A2(_02281_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29321_ (.A1(_11215_),
    .A2(_02285_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29322_ (.A1(_05251_),
    .A2(_05250_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _29323_ (.I(_05252_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29324_ (.A1(_11156_),
    .A2(net946),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29325_ (.A1(_11152_),
    .A2(_11157_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29326_ (.A1(_05254_),
    .A2(_05255_),
    .Z(_05256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29327_ (.A1(_05253_),
    .A2(_05256_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29328_ (.A1(_05254_),
    .A2(_05255_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29329_ (.A1(_05252_),
    .A2(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29330_ (.A1(_05257_),
    .A2(_10403_),
    .A3(_05259_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29331_ (.A1(_10411_),
    .A2(\text_in_r[65] ),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29332_ (.A1(_05260_),
    .A2(\u0.w[1][1] ),
    .A3(_05261_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29333_ (.A1(_05253_),
    .A2(_05258_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29334_ (.A1(_05256_),
    .A2(_05252_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29335_ (.A1(_05263_),
    .A2(_05264_),
    .A3(_11279_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29336_ (.A1(_10489_),
    .A2(\text_in_r[65] ),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29337_ (.A1(_05265_),
    .A2(_07791_),
    .A3(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29338_ (.A1(_05267_),
    .A2(_05262_),
    .ZN(_16111_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29339_ (.A1(_11193_),
    .A2(_11195_),
    .A3(net817),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29340_ (.A1(_11166_),
    .A2(_11194_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29341_ (.A1(net796),
    .A2(net814),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29342_ (.A1(_05269_),
    .A2(_02278_),
    .A3(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29343_ (.A1(_05268_),
    .A2(_05271_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29344_ (.A1(_05272_),
    .A2(_11156_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29345_ (.A1(_05268_),
    .A2(_05271_),
    .A3(_11152_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29346_ (.A1(_05273_),
    .A2(_05274_),
    .B(_10410_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29347_ (.I(\text_in_r[64] ),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29348_ (.A1(_05276_),
    .A2(_11202_),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29349_ (.A1(_05275_),
    .A2(_05277_),
    .B(\u0.w[1][0] ),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29350_ (.A1(_05273_),
    .A2(_05274_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29351_ (.A1(_05279_),
    .A2(_14333_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29352_ (.I(_05277_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29353_ (.A1(_05280_),
    .A2(_07782_),
    .A3(_05281_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29354_ (.A1(_05278_),
    .A2(_05282_),
    .ZN(_16114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29355_ (.A1(\sa30_sub[1] ),
    .A2(_11218_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29356_ (.A1(\sa30_sub[1] ),
    .A2(_11218_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29357_ (.A1(_05283_),
    .A2(_05284_),
    .B(\sa01_sr[2] ),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29358_ (.A1(_11158_),
    .A2(_11216_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29359_ (.A1(\sa30_sub[1] ),
    .A2(_11218_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29360_ (.A1(_05286_),
    .A2(_11250_),
    .A3(_05287_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29361_ (.A1(_05285_),
    .A2(_05288_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _29362_ (.A1(\sa01_sr[1] ),
    .A2(\sa11_sr[2] ),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29363_ (.I(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29364_ (.A1(_05289_),
    .A2(_05291_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29365_ (.A1(_05285_),
    .A2(_05288_),
    .A3(_05290_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29366_ (.A1(_05292_),
    .A2(_05293_),
    .B(net594),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _29367_ (.I(\text_in_r[66] ),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29368_ (.A1(_05295_),
    .A2(net478),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _29369_ (.A1(_05296_),
    .A2(_05294_),
    .B(\u0.w[1][2] ),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29370_ (.A1(_05292_),
    .A2(_05293_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29371_ (.A1(_05298_),
    .A2(_10378_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _29372_ (.I(_05296_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29373_ (.A1(_05299_),
    .A2(_07796_),
    .A3(_05300_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29374_ (.A1(_05301_),
    .A2(_05297_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _29375_ (.I(_05302_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 _29376_ (.I(_05303_),
    .Z(_16130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29377_ (.A1(_05275_),
    .A2(_05277_),
    .B(_07782_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29378_ (.A1(_05280_),
    .A2(\u0.w[1][0] ),
    .A3(_05281_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29379_ (.A1(_05304_),
    .A2(_05305_),
    .ZN(_16105_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _29380_ (.I(_05302_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _29381_ (.I(_05306_),
    .Z(_16123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29382_ (.A1(_05303_),
    .A2(net1121),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29383_ (.A1(_11257_),
    .A2(\sa21_sr[3] ),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29384_ (.A1(_11253_),
    .A2(_11258_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29385_ (.A1(_05308_),
    .A2(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29386_ (.A1(_02356_),
    .A2(_05310_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29387_ (.I(_05310_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29388_ (.A1(_02360_),
    .A2(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29389_ (.A1(_05311_),
    .A2(_05313_),
    .A3(_10403_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29390_ (.A1(_10411_),
    .A2(\text_in_r[67] ),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29391_ (.A1(_05314_),
    .A2(_07801_),
    .A3(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29392_ (.A1(_02356_),
    .A2(_05312_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29393_ (.A1(_02360_),
    .A2(_05310_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29394_ (.A1(_05317_),
    .A2(_10403_),
    .A3(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29395_ (.A1(_10405_),
    .A2(\text_in_r[67] ),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29396_ (.A1(_05319_),
    .A2(\u0.w[1][3] ),
    .A3(_05320_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29397_ (.A1(_05316_),
    .A2(_05321_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29398_ (.I(_05322_),
    .Z(_05323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29399_ (.A1(_05307_),
    .A2(_05323_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29400_ (.A1(\sa21_sr[4] ),
    .A2(_11301_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29401_ (.A1(_05325_),
    .A2(_02374_),
    .B(_13010_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29402_ (.A1(_05325_),
    .A2(_02374_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29403_ (.I(_05327_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29404_ (.A1(_12115_),
    .A2(\text_in_r[68] ),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29405_ (.A1(_05326_),
    .A2(_05328_),
    .B(_05329_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29406_ (.A1(_05330_),
    .A2(\u0.w[1][4] ),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29407_ (.A1(_05325_),
    .A2(_02374_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29408_ (.A1(_05332_),
    .A2(_11348_),
    .A3(_05327_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29409_ (.A1(_05333_),
    .A2(_07808_),
    .A3(_05329_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29410_ (.A1(_05331_),
    .A2(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29411_ (.I(_05335_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29412_ (.A1(_05324_),
    .A2(_05336_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _29413_ (.I(_16112_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29414_ (.A1(_16123_),
    .A2(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29415_ (.A1(_05314_),
    .A2(\u0.w[1][3] ),
    .A3(_05315_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29416_ (.A1(_05319_),
    .A2(_07801_),
    .A3(_05320_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29417_ (.A1(_05340_),
    .A2(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29418_ (.I(_05342_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29419_ (.A1(_05339_),
    .A2(_05343_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29420_ (.A1(net3),
    .A2(_16130_),
    .A3(net1122),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29421_ (.A1(_05344_),
    .A2(_05345_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _29422_ (.A1(\sa30_sub[4] ),
    .A2(\sa21_sr[5] ),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29423_ (.A1(_05347_),
    .A2(\sa01_sr[5] ),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29424_ (.A1(_05347_),
    .A2(\sa01_sr[5] ),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29425_ (.A1(_05348_),
    .A2(_05349_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29426_ (.A1(\sa01_sr[4] ),
    .A2(\sa11_sr[5] ),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29427_ (.A1(_05350_),
    .A2(_05351_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29428_ (.A1(_05350_),
    .A2(_05351_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29429_ (.A1(_10411_),
    .A2(\text_in_r[69] ),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _29430_ (.A1(_05352_),
    .A2(_10526_),
    .A3(_05353_),
    .B(_05354_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29431_ (.A1(_05355_),
    .A2(\u0.w[1][5] ),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29432_ (.A1(_05355_),
    .A2(\u0.w[1][5] ),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29433_ (.A1(_05356_),
    .A2(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29434_ (.I(_05358_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29435_ (.A1(_05337_),
    .A2(_05346_),
    .B(_05359_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29436_ (.A1(_05302_),
    .A2(net1121),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29437_ (.A1(_05361_),
    .A2(_05323_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29438_ (.A1(_16111_),
    .A2(_16105_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29439_ (.A1(_05362_),
    .A2(_05363_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29440_ (.A1(_05330_),
    .A2(_07808_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29441_ (.A1(_05333_),
    .A2(\u0.w[1][4] ),
    .A3(_05329_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29442_ (.A1(_05365_),
    .A2(_05366_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29443_ (.I(_05367_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29444_ (.I(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29445_ (.I(_16121_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29446_ (.A1(_05370_),
    .A2(_05303_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29447_ (.I(_05343_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _29448_ (.I(_16108_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29449_ (.A1(net1098),
    .A2(_05373_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29450_ (.A1(_05371_),
    .A2(_05372_),
    .A3(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29451_ (.A1(_05364_),
    .A2(_05369_),
    .A3(_05375_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29452_ (.A1(\sa30_sub[5] ),
    .A2(\sa21_sr[6] ),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29453_ (.A1(\sa01_sr[6] ),
    .A2(_05377_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29454_ (.A1(\sa01_sr[5] ),
    .A2(\sa11_sr[6] ),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29455_ (.A1(_05378_),
    .A2(_05379_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29456_ (.A1(_05378_),
    .A2(_05379_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29457_ (.A1(_12115_),
    .A2(\text_in_r[70] ),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _29458_ (.A1(_05380_),
    .A2(_11385_),
    .A3(_05381_),
    .B(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29459_ (.A1(_05383_),
    .A2(\u0.w[1][6] ),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29460_ (.A1(_05383_),
    .A2(\u0.w[1][6] ),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29461_ (.A1(_05384_),
    .A2(_05385_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29462_ (.I(_05386_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29463_ (.A1(_05360_),
    .A2(_05376_),
    .B(_05387_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29464_ (.A1(_05266_),
    .A2(\u0.w[1][1] ),
    .A3(_05265_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29465_ (.A1(_07791_),
    .A2(_05260_),
    .A3(_05261_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29466_ (.A1(_05389_),
    .A2(_05390_),
    .ZN(_16106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29467_ (.A1(_16106_),
    .A2(_05303_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29468_ (.A1(_05303_),
    .A2(_16114_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29469_ (.A1(_05391_),
    .A2(_05392_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29470_ (.A1(_16111_),
    .A2(_05306_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29471_ (.I(_05323_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29472_ (.A1(_05394_),
    .A2(_05395_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29473_ (.A1(_05393_),
    .A2(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29474_ (.A1(_05306_),
    .A2(_05370_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29475_ (.I(_05322_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29476_ (.I(_05399_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29477_ (.A1(_05307_),
    .A2(_05398_),
    .B(_05400_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29478_ (.A1(_05397_),
    .A2(_05401_),
    .B(_05369_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29479_ (.A1(net3),
    .A2(_16114_),
    .A3(_05306_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29480_ (.I(_05342_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29481_ (.A1(_05403_),
    .A2(_05404_),
    .A3(_05307_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29482_ (.A1(_05302_),
    .A2(_16109_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29483_ (.A1(_05391_),
    .A2(_05406_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29484_ (.A1(_05407_),
    .A2(_05400_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29485_ (.I(_05336_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29486_ (.A1(_05405_),
    .A2(_05408_),
    .A3(_05409_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29487_ (.I(_05358_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29488_ (.I(_05411_),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29489_ (.A1(_05402_),
    .A2(_05410_),
    .A3(_05412_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29490_ (.A1(\sa30_sub[6] ),
    .A2(_11189_),
    .Z(_05414_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _29491_ (.A1(_14478_),
    .A2(net26),
    .A3(_05414_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29492_ (.A1(_12961_),
    .A2(\text_in_r[71] ),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29493_ (.A1(_05415_),
    .A2(_12965_),
    .B(_05416_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _29494_ (.A1(\u0.w[1][7] ),
    .A2(_05417_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _29495_ (.I(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29496_ (.A1(_05388_),
    .A2(_05413_),
    .B(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29497_ (.A1(net3),
    .A2(_16130_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29498_ (.A1(_16123_),
    .A2(_16108_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29499_ (.A1(_05421_),
    .A2(_05395_),
    .A3(_05422_),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29500_ (.A1(_05303_),
    .A2(_05373_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29501_ (.A1(_05424_),
    .A2(_05404_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29502_ (.A1(_05423_),
    .A2(_05409_),
    .A3(_05425_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29503_ (.A1(_05343_),
    .A2(_05374_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _29504_ (.I(_05427_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29505_ (.A1(_16130_),
    .A2(_16107_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29506_ (.A1(_05428_),
    .A2(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29507_ (.I(_16115_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29508_ (.A1(_05306_),
    .A2(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29509_ (.A1(_05432_),
    .A2(_05342_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29510_ (.A1(_16123_),
    .A2(_16107_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29511_ (.A1(_05433_),
    .A2(_05434_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29512_ (.I(_05368_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29513_ (.A1(_05430_),
    .A2(_05435_),
    .B(_05436_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29514_ (.A1(_05426_),
    .A2(_05437_),
    .B(_05412_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29515_ (.A1(_05374_),
    .A2(_05323_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29516_ (.A1(_16111_),
    .A2(_05303_),
    .A3(_16114_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29517_ (.A1(_05439_),
    .A2(_05440_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29518_ (.I(_16107_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29519_ (.A1(_16130_),
    .A2(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29520_ (.A1(_16123_),
    .A2(_05431_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29521_ (.A1(_05443_),
    .A2(_05444_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29522_ (.I(_05404_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29523_ (.A1(_05445_),
    .A2(_05446_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29524_ (.I(_05336_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29525_ (.A1(_05441_),
    .A2(_05447_),
    .A3(_05448_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29526_ (.A1(_05306_),
    .A2(_16114_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29527_ (.A1(_05450_),
    .A2(_05323_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29528_ (.A1(net7),
    .A2(_16105_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29529_ (.A1(_05451_),
    .A2(_05452_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29530_ (.I(_05343_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29531_ (.A1(_05363_),
    .A2(_05392_),
    .A3(_05454_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29532_ (.A1(_05453_),
    .A2(_05455_),
    .A3(_05369_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _29533_ (.I(_05358_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29534_ (.I(_05457_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29535_ (.A1(_05449_),
    .A2(_05456_),
    .A3(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29536_ (.A1(_05438_),
    .A2(_05459_),
    .A3(_05387_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29537_ (.A1(_05420_),
    .A2(_05460_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29538_ (.A1(_05307_),
    .A2(_05404_),
    .A3(_05434_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29539_ (.A1(_05462_),
    .A2(_05336_),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29540_ (.A1(_16130_),
    .A2(_16109_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29541_ (.A1(_05464_),
    .A2(_05454_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29542_ (.I(_05361_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29543_ (.A1(_05466_),
    .A2(net3),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29544_ (.A1(net1240),
    .A2(_05301_),
    .A3(_05338_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29545_ (.A1(_05467_),
    .A2(_05395_),
    .A3(_05468_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29546_ (.A1(_05463_),
    .A2(_05465_),
    .A3(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29547_ (.A1(net1240),
    .A2(_05301_),
    .A3(net1123),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29548_ (.A1(_05471_),
    .A2(_05323_),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29549_ (.I(_05323_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29550_ (.A1(_05473_),
    .A2(_16128_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29551_ (.A1(_05472_),
    .A2(_05474_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29552_ (.I(_05457_),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29553_ (.A1(_05475_),
    .A2(_05369_),
    .B(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29554_ (.A1(_05470_),
    .A2(_05477_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29555_ (.A1(_05306_),
    .A2(_16117_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29556_ (.A1(_05479_),
    .A2(_05323_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29557_ (.A1(_05467_),
    .A2(_05480_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29558_ (.I(_05406_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29559_ (.A1(_05482_),
    .A2(_05400_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29560_ (.A1(_05481_),
    .A2(_05409_),
    .A3(_05483_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29561_ (.A1(_05482_),
    .A2(_05343_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29562_ (.A1(_05485_),
    .A2(_05368_),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29563_ (.A1(_05467_),
    .A2(_05433_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29564_ (.A1(_05486_),
    .A2(_05487_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29565_ (.I(_05457_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29566_ (.A1(_05484_),
    .A2(_05488_),
    .A3(_05489_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29567_ (.A1(_05478_),
    .A2(_05490_),
    .A3(_05387_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _29568_ (.I(_05443_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _29569_ (.A1(_05492_),
    .A2(_05482_),
    .B(_05400_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29570_ (.I(_05335_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29571_ (.A1(_05344_),
    .A2(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29572_ (.A1(_05493_),
    .A2(_05495_),
    .B(_05359_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29573_ (.A1(_05394_),
    .A2(_05399_),
    .A3(_05471_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29574_ (.A1(_05497_),
    .A2(_05336_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29575_ (.I(_05432_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29576_ (.A1(_05499_),
    .A2(_05454_),
    .A3(_05361_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29577_ (.A1(_05498_),
    .A2(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29578_ (.A1(_05496_),
    .A2(_05501_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29579_ (.A1(_05297_),
    .A2(_05301_),
    .A3(_16112_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29580_ (.I(_05503_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29581_ (.A1(_05504_),
    .A2(_05473_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29582_ (.A1(_05405_),
    .A2(_05505_),
    .A3(_05409_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29583_ (.I(_05367_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29584_ (.A1(_05427_),
    .A2(_05507_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29585_ (.A1(_05306_),
    .A2(_16117_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29586_ (.A1(_05509_),
    .A2(_05503_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29587_ (.A1(_05510_),
    .A2(_05395_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29588_ (.A1(_05508_),
    .A2(_05511_),
    .B(_05476_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29589_ (.A1(_05506_),
    .A2(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29590_ (.I(_05386_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29591_ (.I(_05514_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29592_ (.A1(_05502_),
    .A2(_05513_),
    .A3(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29593_ (.A1(_05491_),
    .A2(_05516_),
    .A3(_05419_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29594_ (.A1(_05461_),
    .A2(_05517_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29595_ (.A1(_05343_),
    .A2(_16130_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29596_ (.I(_05368_),
    .Z(_05519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29597_ (.A1(_05518_),
    .A2(_05363_),
    .B(_05519_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29598_ (.A1(_05394_),
    .A2(_05452_),
    .A3(_05399_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29599_ (.A1(_05520_),
    .A2(_05521_),
    .B(_05359_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29600_ (.A1(_05339_),
    .A2(_05399_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29601_ (.A1(_05523_),
    .A2(_05392_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29602_ (.A1(_05428_),
    .A2(_05307_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29603_ (.A1(_05524_),
    .A2(_05525_),
    .A3(_05369_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29604_ (.A1(_05522_),
    .A2(_05526_),
    .B(_05515_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29605_ (.A1(_05421_),
    .A2(_05404_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29606_ (.A1(net7),
    .A2(_05306_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29607_ (.A1(_05528_),
    .A2(_05529_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29608_ (.A1(_05505_),
    .A2(_05507_),
    .Z(_05531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29609_ (.A1(_05530_),
    .A2(_05531_),
    .B(_05489_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29610_ (.A1(_05425_),
    .A2(_05398_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29611_ (.A1(_05469_),
    .A2(_05533_),
    .A3(_05448_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29612_ (.A1(_05532_),
    .A2(_05534_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29613_ (.I(_05418_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29614_ (.A1(_05527_),
    .A2(_05535_),
    .B(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29615_ (.A1(_05392_),
    .A2(_05395_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29616_ (.A1(_16123_),
    .A2(_05442_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29617_ (.I(_05539_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _29618_ (.A1(_05538_),
    .A2(_05540_),
    .B1(_05427_),
    .B2(_05504_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29619_ (.I(_05507_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29620_ (.A1(_05541_),
    .A2(_05542_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29621_ (.A1(net3),
    .A2(_16114_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29622_ (.I(_05404_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29623_ (.A1(_05544_),
    .A2(_05466_),
    .B(_05545_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29624_ (.A1(_05472_),
    .A2(_05361_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29625_ (.A1(_05546_),
    .A2(_05448_),
    .A3(_05547_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29626_ (.A1(_05543_),
    .A2(_05412_),
    .A3(_05548_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29627_ (.A1(_05440_),
    .A2(_05404_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29628_ (.I(_05422_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29629_ (.A1(_05550_),
    .A2(_05551_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29630_ (.A1(_16123_),
    .A2(_16112_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29631_ (.I(_05553_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29632_ (.I(_05473_),
    .Z(_05555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29633_ (.A1(_05554_),
    .A2(_05555_),
    .B(_05519_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29634_ (.A1(_05552_),
    .A2(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29635_ (.A1(_05371_),
    .A2(_05343_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29636_ (.I(_05558_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29637_ (.A1(_05559_),
    .A2(_05529_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29638_ (.A1(_05529_),
    .A2(_05361_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29639_ (.I(_05399_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29640_ (.A1(_05561_),
    .A2(_05562_),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29641_ (.I(_05368_),
    .Z(_05564_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29642_ (.A1(_05560_),
    .A2(_05563_),
    .A3(_05564_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29643_ (.A1(_05557_),
    .A2(_05565_),
    .A3(_05458_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29644_ (.A1(_05549_),
    .A2(_05515_),
    .A3(_05566_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29645_ (.A1(_05537_),
    .A2(_05567_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29646_ (.A1(_05398_),
    .A2(_05399_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29647_ (.I(_16109_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29648_ (.A1(_16130_),
    .A2(_05570_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29649_ (.A1(_05569_),
    .A2(_05571_),
    .B(_05494_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29650_ (.A1(_05552_),
    .A2(_05572_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _29651_ (.I(_05324_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29652_ (.A1(_05574_),
    .A2(_05403_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29653_ (.A1(_05427_),
    .A2(_05336_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29654_ (.A1(_05575_),
    .A2(_05576_),
    .B(_05476_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29655_ (.A1(_05573_),
    .A2(_05577_),
    .B(_05387_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29656_ (.A1(_05425_),
    .A2(_05434_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29657_ (.A1(_05399_),
    .A2(_16130_),
    .A3(_16114_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29658_ (.A1(_05580_),
    .A2(_05368_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29659_ (.I(_05581_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29660_ (.A1(_05579_),
    .A2(_05582_),
    .A3(_05483_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29661_ (.A1(_05451_),
    .A2(_05429_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29662_ (.A1(_05344_),
    .A2(_05391_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29663_ (.A1(_05584_),
    .A2(_05585_),
    .A3(_05409_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29664_ (.A1(_05583_),
    .A2(_05586_),
    .A3(_05458_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29665_ (.A1(_05578_),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29666_ (.A1(_05362_),
    .A2(_05429_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29667_ (.A1(_05589_),
    .A2(_05457_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29668_ (.A1(_05393_),
    .A2(_05561_),
    .B(_05545_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29669_ (.A1(_05590_),
    .A2(_05591_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29670_ (.A1(_05451_),
    .A2(_05421_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29671_ (.A1(_05593_),
    .A2(_05585_),
    .A3(_05359_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29672_ (.A1(_05592_),
    .A2(_05542_),
    .A3(_05594_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29673_ (.I(_16131_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29674_ (.A1(_05545_),
    .A2(_05596_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29675_ (.A1(_05433_),
    .A2(_05403_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29676_ (.A1(_05489_),
    .A2(_05597_),
    .B(_05598_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _29677_ (.I(_05514_),
    .Z(_05600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29678_ (.A1(_05599_),
    .A2(_05448_),
    .B(_05600_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29679_ (.A1(_05595_),
    .A2(_05601_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29680_ (.A1(_05588_),
    .A2(_05602_),
    .A3(_05536_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29681_ (.A1(_05568_),
    .A2(_05603_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29682_ (.A1(_05467_),
    .A2(_05468_),
    .B(_05395_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29683_ (.A1(_05604_),
    .A2(_05498_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29684_ (.A1(_05523_),
    .A2(_05371_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29685_ (.A1(_05394_),
    .A2(_05363_),
    .A3(_05372_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _29686_ (.I(_05335_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29687_ (.A1(_05606_),
    .A2(_05607_),
    .B(_05608_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29688_ (.A1(_05605_),
    .A2(_05609_),
    .B(_05412_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29689_ (.A1(_05345_),
    .A2(_05555_),
    .B(_05519_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29690_ (.A1(_05440_),
    .A2(_05446_),
    .A3(_05398_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29691_ (.A1(_05611_),
    .A2(_05612_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29692_ (.A1(_05464_),
    .A2(_05450_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29693_ (.A1(_05614_),
    .A2(_05446_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29694_ (.A1(_05421_),
    .A2(_05400_),
    .A3(_05374_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29695_ (.A1(_05615_),
    .A2(_05616_),
    .A3(_05564_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29696_ (.A1(_05613_),
    .A2(_05617_),
    .A3(_05458_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29697_ (.A1(_05610_),
    .A2(_05387_),
    .A3(_05618_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29698_ (.A1(_05479_),
    .A2(_05343_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29699_ (.A1(_05620_),
    .A2(_05361_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29700_ (.A1(_05471_),
    .A2(_05343_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29701_ (.A1(_05622_),
    .A2(_05374_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29702_ (.A1(_05621_),
    .A2(_05623_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29703_ (.A1(_05624_),
    .A2(_05608_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29704_ (.A1(_05391_),
    .A2(_05372_),
    .A3(_05509_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29705_ (.A1(net1241),
    .A2(_05301_),
    .A3(_16121_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29706_ (.A1(_05450_),
    .A2(_05473_),
    .A3(_05627_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29707_ (.A1(_05626_),
    .A2(_05436_),
    .A3(_05628_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29708_ (.A1(_05625_),
    .A2(_05629_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29709_ (.A1(_05630_),
    .A2(_05458_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29710_ (.A1(_05450_),
    .A2(_05503_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29711_ (.A1(_05627_),
    .A2(_05473_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29712_ (.A1(_05632_),
    .A2(_05562_),
    .B(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _29713_ (.I(_05509_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29714_ (.A1(_05635_),
    .A2(_05562_),
    .B(_05494_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29715_ (.A1(_05634_),
    .A2(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29716_ (.A1(_05529_),
    .A2(_05372_),
    .A3(_05468_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29717_ (.A1(_05638_),
    .A2(_05511_),
    .A3(_05608_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29718_ (.A1(_05637_),
    .A2(_05639_),
    .A3(_05359_),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29719_ (.A1(_05631_),
    .A2(_05515_),
    .A3(_05640_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29720_ (.A1(_05619_),
    .A2(_05641_),
    .A3(_05536_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29721_ (.A1(_05425_),
    .A2(_05467_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29722_ (.A1(_16128_),
    .A2(_05400_),
    .B(_05519_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29723_ (.A1(_05643_),
    .A2(_05644_),
    .B(_05411_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _29724_ (.A1(_16106_),
    .A2(_05303_),
    .B(_05323_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29725_ (.A1(_05646_),
    .A2(_05361_),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29726_ (.A1(_05647_),
    .A2(_05369_),
    .A3(_05497_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29727_ (.A1(_05645_),
    .A2(_05648_),
    .B(_05386_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29728_ (.A1(_05622_),
    .A2(_05444_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29729_ (.A1(_05396_),
    .A2(_05492_),
    .B(_05650_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29730_ (.A1(_05651_),
    .A2(_05542_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29731_ (.A1(_05394_),
    .A2(_05452_),
    .A3(_05404_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29732_ (.A1(_05653_),
    .A2(_05336_),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29733_ (.A1(_05555_),
    .A2(_05596_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29734_ (.A1(_05654_),
    .A2(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29735_ (.A1(_05652_),
    .A2(_05656_),
    .A3(_05412_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29736_ (.A1(_05649_),
    .A2(_05657_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29737_ (.A1(_05598_),
    .A2(_05507_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29738_ (.A1(_05391_),
    .A2(_05307_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29739_ (.A1(_05406_),
    .A2(_05553_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29740_ (.A1(_05660_),
    .A2(_05661_),
    .B(_05545_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29741_ (.A1(_05659_),
    .A2(_05662_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29742_ (.A1(_05540_),
    .A2(_05400_),
    .B(_05507_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29743_ (.A1(_05428_),
    .A2(_05468_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29744_ (.A1(_05665_),
    .A2(_05664_),
    .B(_05411_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29745_ (.A1(_05663_),
    .A2(_05666_),
    .B(_05600_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29746_ (.A1(_05345_),
    .A2(_05473_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29747_ (.A1(_05399_),
    .A2(_16126_),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29748_ (.A1(_05668_),
    .A2(_05669_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29749_ (.A1(_05670_),
    .A2(_05436_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29750_ (.A1(_05562_),
    .A2(_16135_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29751_ (.A1(_05607_),
    .A2(_05564_),
    .A3(_05672_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29752_ (.A1(_05671_),
    .A2(_05412_),
    .A3(_05673_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29753_ (.A1(_05667_),
    .A2(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29754_ (.A1(_05658_),
    .A2(_05675_),
    .A3(_05419_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29755_ (.A1(_05642_),
    .A2(_05676_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29756_ (.A1(_05646_),
    .A2(_05374_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29757_ (.A1(_05451_),
    .A2(_05363_),
    .ZN(_05678_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29758_ (.A1(_05677_),
    .A2(_05678_),
    .A3(_05448_),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29759_ (.I(_05424_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29760_ (.A1(_05680_),
    .A2(_05404_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29761_ (.A1(_05593_),
    .A2(_05681_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29762_ (.A1(_05682_),
    .A2(_05542_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29763_ (.A1(_05679_),
    .A2(_05683_),
    .A3(_05412_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29764_ (.A1(_05392_),
    .A2(_05395_),
    .A3(_05444_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29765_ (.A1(_05424_),
    .A2(_05454_),
    .A3(_05539_),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29766_ (.A1(_05685_),
    .A2(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29767_ (.A1(_05687_),
    .A2(_05542_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29768_ (.A1(_05422_),
    .A2(_05399_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29769_ (.A1(_05689_),
    .A2(_05391_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29770_ (.A1(_05398_),
    .A2(_05468_),
    .A3(_05372_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29771_ (.A1(_05690_),
    .A2(_05409_),
    .A3(_05691_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29772_ (.A1(_05688_),
    .A2(_05692_),
    .A3(_05489_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29773_ (.A1(_05684_),
    .A2(_05387_),
    .A3(_05693_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29774_ (.I(_05529_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29775_ (.A1(_05558_),
    .A2(_05695_),
    .B(_05507_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29776_ (.A1(_05620_),
    .A2(_05422_),
    .Z(_05697_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29777_ (.A1(_05696_),
    .A2(_05697_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29778_ (.A1(_05452_),
    .A2(_05392_),
    .A3(_05336_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29779_ (.A1(_05446_),
    .A2(_16123_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29780_ (.A1(_05699_),
    .A2(_05700_),
    .B(_05476_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29781_ (.A1(_05698_),
    .A2(_05701_),
    .B(_05387_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29782_ (.A1(_05392_),
    .A2(_05444_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29783_ (.A1(_05703_),
    .A2(_05646_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29784_ (.A1(net7),
    .A2(_16105_),
    .B(_16123_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29785_ (.A1(_05705_),
    .A2(_05472_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29786_ (.A1(_05704_),
    .A2(_05608_),
    .A3(_05706_),
    .ZN(_05707_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29787_ (.A1(_16130_),
    .A2(_05431_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29788_ (.I(_05708_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29789_ (.A1(_05439_),
    .A2(_05709_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29790_ (.A1(_05710_),
    .A2(_05455_),
    .A3(_05436_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29791_ (.A1(_05707_),
    .A2(_05711_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29792_ (.A1(_05712_),
    .A2(_05458_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29793_ (.A1(_05702_),
    .A2(_05713_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29794_ (.A1(_05694_),
    .A2(_05714_),
    .A3(_05419_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29795_ (.A1(_05433_),
    .A2(_05394_),
    .Z(_05716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29796_ (.I(_05681_),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29797_ (.A1(_05716_),
    .A2(_05717_),
    .B(_05411_),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29798_ (.I(_05374_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29799_ (.A1(_05719_),
    .A2(_05323_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29800_ (.A1(_05358_),
    .A2(_05720_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29801_ (.A1(_05721_),
    .A2(_05486_),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29802_ (.A1(_05718_),
    .A2(_05722_),
    .B(_05600_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29803_ (.A1(_05574_),
    .A2(_05374_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29804_ (.A1(_05570_),
    .A2(_05338_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29805_ (.A1(_05306_),
    .A2(_05725_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29806_ (.A1(_05726_),
    .A2(_05343_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29807_ (.A1(_05727_),
    .A2(_05371_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29808_ (.A1(_05724_),
    .A2(_05411_),
    .A3(_05728_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29809_ (.A1(_05635_),
    .A2(_05454_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29810_ (.A1(_05621_),
    .A2(_05457_),
    .A3(_05730_),
    .ZN(_05731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29811_ (.A1(_05729_),
    .A2(_05731_),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29812_ (.A1(_05732_),
    .A2(_05448_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29813_ (.A1(_05723_),
    .A2(_05733_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29814_ (.I(_05307_),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29815_ (.A1(_05735_),
    .A2(_05635_),
    .B(_05404_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29816_ (.A1(_05439_),
    .A2(_05371_),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29817_ (.A1(_05736_),
    .A2(_05737_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29818_ (.A1(_05738_),
    .A2(_05436_),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29819_ (.A1(_05521_),
    .A2(_05462_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29820_ (.A1(_05740_),
    .A2(_05608_),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29821_ (.A1(_05739_),
    .A2(_05489_),
    .A3(_05741_),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29822_ (.A1(_05480_),
    .A2(_05726_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29823_ (.A1(_05598_),
    .A2(_05743_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29824_ (.A1(_05744_),
    .A2(_05608_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29825_ (.A1(_05628_),
    .A2(_05436_),
    .B(_05457_),
    .ZN(_05746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29826_ (.A1(_05745_),
    .A2(_05746_),
    .B(_05386_),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29827_ (.A1(_05742_),
    .A2(_05747_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29828_ (.A1(_05734_),
    .A2(_05748_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29829_ (.A1(_05749_),
    .A2(_05536_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29830_ (.A1(_05715_),
    .A2(_05750_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29831_ (.A1(_05646_),
    .A2(_05434_),
    .B(_05436_),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29832_ (.A1(_05751_),
    .A2(_05469_),
    .ZN(_05752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29833_ (.A1(_05646_),
    .A2(_05467_),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29834_ (.A1(_05753_),
    .A2(_05369_),
    .A3(_05606_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29835_ (.A1(_05752_),
    .A2(_05754_),
    .A3(_05412_),
    .ZN(_05755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29836_ (.A1(_05569_),
    .A2(_05424_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29837_ (.A1(_05481_),
    .A2(_05756_),
    .A3(_05409_),
    .ZN(_05757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29838_ (.A1(_05635_),
    .A2(_05545_),
    .B(_05494_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29839_ (.A1(_05518_),
    .A2(_16108_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29840_ (.A1(_05758_),
    .A2(_05511_),
    .A3(_05759_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29841_ (.A1(_05757_),
    .A2(_05760_),
    .A3(_05458_),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29842_ (.A1(_05755_),
    .A2(_05761_),
    .A3(_05387_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29843_ (.A1(_05593_),
    .A2(_05653_),
    .A3(_05409_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29844_ (.A1(_05391_),
    .A2(_05363_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29845_ (.A1(_05764_),
    .A2(_05562_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29846_ (.A1(_05529_),
    .A2(_05429_),
    .A3(_05372_),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29847_ (.A1(_05765_),
    .A2(_05766_),
    .A3(_05564_),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29848_ (.A1(_05763_),
    .A2(_05767_),
    .A3(_05412_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29849_ (.A1(_05421_),
    .A2(_05454_),
    .A3(_05361_),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29850_ (.A1(_05589_),
    .A2(_05769_),
    .A3(_05608_),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _29851_ (.A1(_05480_),
    .A2(_05494_),
    .A3(_05482_),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29852_ (.A1(_05770_),
    .A2(_05489_),
    .A3(_05771_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29853_ (.A1(_05768_),
    .A2(_05515_),
    .A3(_05772_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29854_ (.A1(_05762_),
    .A2(_05773_),
    .A3(_05419_),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29855_ (.A1(_05405_),
    .A2(_05336_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29856_ (.A1(_05523_),
    .A2(_05471_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29857_ (.A1(_05775_),
    .A2(_05776_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29858_ (.A1(_05571_),
    .A2(_05399_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29859_ (.A1(_05778_),
    .A2(_05507_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29860_ (.A1(_05779_),
    .A2(_05550_),
    .B(_05359_),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29861_ (.A1(_05777_),
    .A2(_05780_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29862_ (.A1(_05451_),
    .A2(_05371_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29863_ (.A1(_05518_),
    .A2(_05519_),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29864_ (.A1(_05782_),
    .A2(_05783_),
    .B(_05476_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29865_ (.A1(_05421_),
    .A2(_05400_),
    .A3(_05434_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29866_ (.A1(_05585_),
    .A2(_05785_),
    .A3(_05564_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29867_ (.A1(_05784_),
    .A2(_05786_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29868_ (.A1(_05781_),
    .A2(_05515_),
    .A3(_05787_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29869_ (.A1(_05764_),
    .A2(_05454_),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29870_ (.A1(_05480_),
    .A2(_05450_),
    .ZN(_05790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29871_ (.A1(_05789_),
    .A2(_05369_),
    .A3(_05790_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29872_ (.A1(_05493_),
    .A2(_05455_),
    .A3(_05409_),
    .ZN(_05792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29873_ (.A1(_05791_),
    .A2(_05792_),
    .A3(_05359_),
    .ZN(_05793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29874_ (.I(_16119_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29875_ (.A1(_05794_),
    .A2(_05400_),
    .B(_05507_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29876_ (.I(_05622_),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29877_ (.A1(_05795_),
    .A2(_05796_),
    .B(_05411_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29878_ (.A1(_05529_),
    .A2(_05450_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29879_ (.A1(_05798_),
    .A2(_05473_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29880_ (.A1(_05480_),
    .A2(_05529_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29881_ (.A1(_05799_),
    .A2(_05800_),
    .A3(_05436_),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29882_ (.A1(_05797_),
    .A2(_05801_),
    .B(_05600_),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29883_ (.A1(_05793_),
    .A2(_05802_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29884_ (.A1(_05788_),
    .A2(_05536_),
    .A3(_05803_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29885_ (.A1(_05774_),
    .A2(_05804_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29886_ (.A1(net7),
    .A2(_05454_),
    .B(_05368_),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29887_ (.A1(_05789_),
    .A2(_05805_),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29888_ (.A1(_05806_),
    .A2(_05489_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29889_ (.A1(_05705_),
    .A2(_05709_),
    .A3(_05454_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29890_ (.A1(_05324_),
    .A2(_05544_),
    .B(_05519_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29891_ (.A1(_05808_),
    .A2(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29892_ (.A1(_05807_),
    .A2(_05810_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29893_ (.I(_05394_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29894_ (.A1(_05778_),
    .A2(_05812_),
    .Z(_05813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29895_ (.A1(_05813_),
    .A2(_05759_),
    .B(_05608_),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29896_ (.A1(_05427_),
    .A2(_05492_),
    .B(_05494_),
    .C(_05633_),
    .ZN(_05815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29897_ (.A1(_05815_),
    .A2(_05359_),
    .ZN(_05816_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29898_ (.A1(_05814_),
    .A2(_05816_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29899_ (.A1(_05811_),
    .A2(_05817_),
    .B(_05387_),
    .ZN(_05818_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29900_ (.A1(_05439_),
    .A2(_05436_),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29901_ (.A1(_05819_),
    .A2(_05736_),
    .B(_05476_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29902_ (.A1(_05393_),
    .A2(_05446_),
    .B(_05523_),
    .ZN(_05821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29903_ (.A1(_05821_),
    .A2(_05542_),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29904_ (.A1(_05820_),
    .A2(_05822_),
    .B(_05386_),
    .ZN(_05823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29905_ (.A1(_05446_),
    .A2(_16112_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29906_ (.A1(_05467_),
    .A2(_05620_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29907_ (.A1(_05486_),
    .A2(_05824_),
    .A3(_05825_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29908_ (.A1(_05559_),
    .A2(_05339_),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29909_ (.A1(_05827_),
    .A2(_05409_),
    .A3(_05408_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29910_ (.A1(_05826_),
    .A2(_05828_),
    .A3(_05458_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29911_ (.A1(_05823_),
    .A2(_05829_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29912_ (.A1(_05818_),
    .A2(_05419_),
    .A3(_05830_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29913_ (.A1(_16114_),
    .A2(_05545_),
    .B(_05519_),
    .ZN(_05832_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29914_ (.A1(_05832_),
    .A2(_05453_),
    .B(_05411_),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29915_ (.A1(_05428_),
    .A2(_05345_),
    .ZN(_05834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29916_ (.A1(_05620_),
    .A2(_05529_),
    .ZN(_05835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29917_ (.A1(_05834_),
    .A2(_05835_),
    .A3(_05564_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29918_ (.A1(_05833_),
    .A2(_05836_),
    .B(_05386_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29919_ (.A1(_05632_),
    .A2(_05555_),
    .ZN(_05838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29920_ (.A1(_05775_),
    .A2(_05838_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29921_ (.A1(_05403_),
    .A2(_05555_),
    .A3(_05371_),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29922_ (.A1(_05708_),
    .A2(_05545_),
    .B(_05494_),
    .ZN(_05841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29923_ (.A1(_05840_),
    .A2(_05841_),
    .B(_05489_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29924_ (.A1(_05839_),
    .A2(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29925_ (.A1(_05837_),
    .A2(_05843_),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29926_ (.A1(_05431_),
    .A2(_05372_),
    .B(_05507_),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29927_ (.A1(_05403_),
    .A2(_05562_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29928_ (.A1(_05845_),
    .A2(_05846_),
    .B(_05476_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29929_ (.A1(_05689_),
    .A2(_05371_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29930_ (.A1(_05428_),
    .A2(_05499_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29931_ (.A1(_05848_),
    .A2(_05849_),
    .A3(_05564_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29932_ (.A1(_05847_),
    .A2(_05850_),
    .B(_05600_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29933_ (.A1(_05393_),
    .A2(_05561_),
    .B(_05562_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29934_ (.I(_05727_),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29935_ (.A1(_05852_),
    .A2(_05448_),
    .A3(_05853_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29936_ (.A1(_05531_),
    .A2(_05558_),
    .B(_05411_),
    .ZN(_05855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29937_ (.A1(_05854_),
    .A2(_05855_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29938_ (.A1(_05851_),
    .A2(_05856_),
    .ZN(_05857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29939_ (.A1(_05844_),
    .A2(_05857_),
    .A3(_05536_),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29940_ (.A1(_05831_),
    .A2(_05858_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29941_ (.A1(_05467_),
    .A2(_05446_),
    .A3(_05392_),
    .ZN(_05859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29942_ (.A1(_05472_),
    .A2(_05726_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29943_ (.A1(_05859_),
    .A2(_05448_),
    .A3(_05860_),
    .ZN(_05861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29944_ (.A1(_05708_),
    .A2(_05562_),
    .B(_05494_),
    .ZN(_05862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29945_ (.A1(_05450_),
    .A2(net3),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29946_ (.A1(_05863_),
    .A2(_05545_),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29947_ (.A1(_05862_),
    .A2(_05864_),
    .B(_05600_),
    .ZN(_05865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29948_ (.A1(_05861_),
    .A2(_05865_),
    .B(_05489_),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29949_ (.A1(_05620_),
    .A2(_05398_),
    .B(_05507_),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29950_ (.A1(_05660_),
    .A2(_05446_),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29951_ (.A1(_05867_),
    .A2(_05485_),
    .A3(_05868_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29952_ (.A1(_05451_),
    .A2(_05471_),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29953_ (.A1(_16123_),
    .A2(_05725_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29954_ (.A1(_05635_),
    .A2(_05871_),
    .B(_05372_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29955_ (.A1(_05870_),
    .A2(_05872_),
    .A3(_05564_),
    .ZN(_05873_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29956_ (.A1(_05869_),
    .A2(_05515_),
    .A3(_05873_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29957_ (.A1(_05866_),
    .A2(_05874_),
    .B(_05536_),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29958_ (.A1(_05393_),
    .A2(_05812_),
    .ZN(_05876_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29959_ (.A1(_05876_),
    .A2(_05400_),
    .B(_05778_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29960_ (.A1(_05551_),
    .A2(_05395_),
    .B(_05368_),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29961_ (.A1(_05877_),
    .A2(_05878_),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29962_ (.A1(_05720_),
    .A2(_05368_),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29963_ (.A1(_05670_),
    .A2(_05880_),
    .B(_05514_),
    .ZN(_05881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29964_ (.A1(_05881_),
    .A2(_05879_),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29965_ (.A1(_05464_),
    .A2(_05509_),
    .B(_05473_),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29966_ (.A1(_05540_),
    .A2(_05473_),
    .Z(_05884_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29967_ (.A1(_05883_),
    .A2(_05494_),
    .A3(_05884_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29968_ (.A1(_05646_),
    .A2(_05363_),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29969_ (.A1(_16124_),
    .A2(_16133_),
    .Z(_05887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29970_ (.A1(_05473_),
    .A2(_05887_),
    .B(_05368_),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29971_ (.A1(_05886_),
    .A2(_05888_),
    .Z(_05889_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29972_ (.A1(_05885_),
    .A2(_05889_),
    .B(_05600_),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29973_ (.A1(_05882_),
    .A2(_05890_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29974_ (.A1(_05891_),
    .A2(_05458_),
    .ZN(_05892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29975_ (.A1(_05875_),
    .A2(_05892_),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29976_ (.A1(_05452_),
    .A2(_05454_),
    .Z(_05894_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29977_ (.A1(_05894_),
    .A2(_05569_),
    .B(_05392_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29978_ (.A1(_05895_),
    .A2(_05542_),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29979_ (.A1(_05555_),
    .A2(net7),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29980_ (.A1(_05699_),
    .A2(_05897_),
    .B(_05359_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29981_ (.A1(_05896_),
    .A2(_05898_),
    .ZN(_05899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29982_ (.A1(_05736_),
    .A2(_05878_),
    .B(_05476_),
    .ZN(_05900_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29983_ (.A1(_05364_),
    .A2(_05369_),
    .A3(_05528_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29984_ (.A1(_05900_),
    .A2(_05901_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29985_ (.A1(_05899_),
    .A2(_05902_),
    .A3(_05515_),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29986_ (.A1(_05551_),
    .A2(_05558_),
    .B(_05582_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29987_ (.I(_16125_),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29988_ (.A1(_05905_),
    .A2(_05372_),
    .B(_05519_),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29989_ (.A1(_05906_),
    .A2(_05835_),
    .B(_05411_),
    .ZN(_05907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29990_ (.A1(_05904_),
    .A2(_05907_),
    .ZN(_05908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29991_ (.A1(_05604_),
    .A2(_05448_),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29992_ (.A1(_05433_),
    .A2(_05494_),
    .ZN(_05910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29993_ (.A1(_05910_),
    .A2(_05800_),
    .B(_05476_),
    .ZN(_05911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29994_ (.A1(_05909_),
    .A2(_05911_),
    .ZN(_05912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29995_ (.A1(_05908_),
    .A2(_05912_),
    .A3(_05387_),
    .ZN(_05913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29996_ (.A1(_05903_),
    .A2(_05913_),
    .A3(_05536_),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29997_ (.A1(_05893_),
    .A2(_05914_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29998_ (.A1(_05440_),
    .A2(_05434_),
    .Z(_05915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29999_ (.A1(_05915_),
    .A2(_05555_),
    .ZN(_05916_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _30000_ (.A1(_05551_),
    .A2(_05395_),
    .A3(_05432_),
    .Z(_05917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30001_ (.A1(_05916_),
    .A2(_05448_),
    .A3(_05917_),
    .ZN(_05918_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30002_ (.A1(_05735_),
    .A2(net7),
    .B(_05555_),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30003_ (.A1(_05919_),
    .A2(_05542_),
    .A3(_05743_),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30004_ (.A1(_05918_),
    .A2(_05920_),
    .A3(_05458_),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30005_ (.A1(_05528_),
    .A2(_05778_),
    .ZN(_05922_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _30006_ (.A1(_05922_),
    .A2(_05608_),
    .A3(_05434_),
    .Z(_05923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30007_ (.A1(_05555_),
    .A2(_16112_),
    .ZN(_05924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30008_ (.A1(_05886_),
    .A2(_05924_),
    .B(_05608_),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30009_ (.A1(_05923_),
    .A2(_05925_),
    .B(_05412_),
    .ZN(_05926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30010_ (.A1(_05921_),
    .A2(_05926_),
    .A3(_05515_),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30011_ (.A1(_05794_),
    .A2(_05545_),
    .B(_05519_),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30012_ (.A1(_05928_),
    .A2(_05465_),
    .B(_05411_),
    .ZN(_05929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30013_ (.A1(_05863_),
    .A2(_05562_),
    .ZN(_05930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30014_ (.A1(_05585_),
    .A2(_05369_),
    .A3(_05930_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30015_ (.A1(_05929_),
    .A2(_05931_),
    .B(_05600_),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30016_ (.A1(_05425_),
    .A2(_05422_),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30017_ (.A1(_05574_),
    .A2(_05529_),
    .ZN(_05934_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30018_ (.A1(_05933_),
    .A2(_05934_),
    .A3(_05542_),
    .ZN(_05935_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30019_ (.A1(_05680_),
    .A2(_05635_),
    .B(_05562_),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30020_ (.A1(_16133_),
    .A2(_05372_),
    .B(_05519_),
    .ZN(_05937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30021_ (.A1(_05936_),
    .A2(_05937_),
    .B(_05476_),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30022_ (.A1(_05935_),
    .A2(_05938_),
    .ZN(_05939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30023_ (.A1(_05932_),
    .A2(_05939_),
    .B(_05536_),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30024_ (.A1(_05927_),
    .A2(_05940_),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30025_ (.I(_05799_),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30026_ (.A1(_05942_),
    .A2(_05581_),
    .ZN(_05943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30027_ (.A1(_05915_),
    .A2(_05446_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30028_ (.A1(_05943_),
    .A2(_05944_),
    .ZN(_05945_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30029_ (.A1(_05569_),
    .A2(_05436_),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30030_ (.A1(_05946_),
    .A2(_05800_),
    .B(_05386_),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30031_ (.A1(_05945_),
    .A2(_05947_),
    .B(_05359_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30032_ (.A1(_05812_),
    .A2(_05555_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30033_ (.A1(_05654_),
    .A2(_05765_),
    .A3(_05949_),
    .ZN(_05950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30034_ (.A1(_05395_),
    .A2(_16105_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30035_ (.A1(_05769_),
    .A2(_05951_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30036_ (.A1(_05952_),
    .A2(_05542_),
    .B(_05600_),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30037_ (.A1(_05950_),
    .A2(_05953_),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30038_ (.A1(_05948_),
    .A2(_05954_),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30039_ (.A1(_05720_),
    .A2(_05336_),
    .Z(_05956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30040_ (.A1(_05561_),
    .A2(_05545_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30041_ (.A1(_05956_),
    .A2(_05957_),
    .B(_05600_),
    .ZN(_05958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30042_ (.A1(_05467_),
    .A2(_05446_),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30043_ (.A1(_05689_),
    .A2(_05440_),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30044_ (.A1(_05959_),
    .A2(_05960_),
    .A3(_05564_),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30045_ (.A1(_05958_),
    .A2(_05961_),
    .B(_05489_),
    .ZN(_05962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30046_ (.A1(_05533_),
    .A2(_05724_),
    .A3(_05564_),
    .ZN(_05963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30047_ (.A1(_05867_),
    .A2(_05647_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30048_ (.A1(_05963_),
    .A2(_05964_),
    .A3(_05515_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30049_ (.A1(_05962_),
    .A2(_05965_),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30050_ (.A1(_05955_),
    .A2(_05966_),
    .A3(_05536_),
    .ZN(_05967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30051_ (.A1(_05941_),
    .A2(_05967_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30052_ (.A1(_03026_),
    .A2(_03018_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30053_ (.A1(_03022_),
    .A2(_12024_),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30054_ (.A1(_05969_),
    .A2(_05968_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30055_ (.I(_05970_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30056_ (.A1(_11973_),
    .A2(net1170),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30057_ (.A1(_11969_),
    .A2(_11959_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30058_ (.A1(_05973_),
    .A2(_05972_),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30059_ (.A1(_05971_),
    .A2(_05974_),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30060_ (.I(_05974_),
    .ZN(_05976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30061_ (.A1(_05976_),
    .A2(_05970_),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30062_ (.A1(_05975_),
    .A2(_05977_),
    .A3(_10479_),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30063_ (.I(\u0.w[2][1] ),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30064_ (.A1(_10489_),
    .A2(\text_in_r[33] ),
    .Z(_05980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30065_ (.A1(_05978_),
    .A2(_05979_),
    .A3(_05980_),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30066_ (.A1(_05971_),
    .A2(_05976_),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30067_ (.A1(_05970_),
    .A2(_05974_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30068_ (.A1(_05983_),
    .A2(_10479_),
    .A3(_05982_),
    .ZN(_05984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30069_ (.A1(_10483_),
    .A2(\text_in_r[33] ),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30070_ (.A1(_05985_),
    .A2(\u0.w[2][1] ),
    .A3(_05984_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30071_ (.A1(_05981_),
    .A2(_05986_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _30072_ (.I(_05987_),
    .Z(_16143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30073_ (.A1(_12005_),
    .A2(_12251_),
    .A3(_12007_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30074_ (.A1(_11981_),
    .A2(_12006_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30075_ (.A1(net1180),
    .A2(\sa20_sub[0] ),
    .ZN(_05990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30076_ (.A1(_05989_),
    .A2(_03015_),
    .A3(_05990_),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30077_ (.A1(_05988_),
    .A2(_05991_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30078_ (.A1(_11973_),
    .A2(_05992_),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30079_ (.A1(_05988_),
    .A2(_11969_),
    .A3(_05991_),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30080_ (.A1(_05993_),
    .A2(net1211),
    .B(_10586_),
    .ZN(_05995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30081_ (.I(\text_in_r[32] ),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30082_ (.A1(_05996_),
    .A2(_10381_),
    .Z(_05997_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30083_ (.A1(_05995_),
    .A2(_05997_),
    .B(\u0.w[2][0] ),
    .ZN(_05998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30084_ (.A1(_05993_),
    .A2(_05994_),
    .ZN(_05999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30085_ (.A1(_10549_),
    .A2(_05999_),
    .ZN(_06000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30086_ (.I(\u0.w[2][0] ),
    .ZN(_06001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30087_ (.I(_05997_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30088_ (.A1(net1194),
    .A2(_06001_),
    .A3(_06002_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30089_ (.A1(_06003_),
    .A2(_05998_),
    .ZN(_16146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30090_ (.A1(\sa31_sub[1] ),
    .A2(_12027_),
    .Z(_06004_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30091_ (.A1(\sa31_sub[1] ),
    .A2(_12027_),
    .ZN(_06005_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30092_ (.A1(_06005_),
    .A2(_06004_),
    .B(\sa02_sr[2] ),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30093_ (.A1(net1167),
    .A2(_12025_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30094_ (.A1(\sa31_sub[1] ),
    .A2(_12027_),
    .ZN(_06008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30095_ (.A1(_06007_),
    .A2(_12057_),
    .A3(_06008_),
    .ZN(_06009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30096_ (.A1(_06006_),
    .A2(_06009_),
    .ZN(_06010_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30097_ (.A1(\sa02_sr[1] ),
    .A2(\sa12_sr[2] ),
    .ZN(_06011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30098_ (.I(_06011_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30099_ (.A1(_06012_),
    .A2(_06010_),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30100_ (.A1(_06011_),
    .A2(_06009_),
    .A3(_06006_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30101_ (.A1(_06013_),
    .A2(_06014_),
    .B(_10482_),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30102_ (.I(\text_in_r[34] ),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30103_ (.A1(_06016_),
    .A2(_11202_),
    .Z(_06017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30104_ (.I(\u0.w[2][2] ),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _30105_ (.A1(_06017_),
    .A2(_06015_),
    .B(_06018_),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30106_ (.A1(_06013_),
    .A2(_06014_),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30107_ (.A1(_06020_),
    .A2(_14333_),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30108_ (.I(_06017_),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30109_ (.A1(_06021_),
    .A2(\u0.w[2][2] ),
    .A3(_06022_),
    .ZN(_06023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30110_ (.A1(_06019_),
    .A2(_06023_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _30111_ (.I(_06024_),
    .Z(_06025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _30112_ (.I(_06025_),
    .Z(_16162_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30113_ (.A1(_05995_),
    .A2(_05997_),
    .B(_06001_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30114_ (.A1(_06002_),
    .A2(\u0.w[2][0] ),
    .A3(_06000_),
    .ZN(_06027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30115_ (.A1(_06027_),
    .A2(_06026_),
    .ZN(_16137_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30116_ (.A1(_06015_),
    .A2(_06017_),
    .B(\u0.w[2][2] ),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30117_ (.A1(_06021_),
    .A2(_06018_),
    .A3(_06022_),
    .ZN(_06029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30118_ (.A1(_06028_),
    .A2(_06029_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _30119_ (.I(_06030_),
    .Z(_06031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _30120_ (.I(_06031_),
    .Z(_16155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30121_ (.A1(net1181),
    .A2(_16137_),
    .ZN(_06032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30122_ (.A1(_12064_),
    .A2(\sa20_sub[3] ),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30123_ (.A1(_12060_),
    .A2(_12065_),
    .ZN(_06034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30124_ (.A1(_06033_),
    .A2(_06034_),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30125_ (.A1(_03108_),
    .A2(_06035_),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30126_ (.A1(_12060_),
    .A2(\sa20_sub[3] ),
    .ZN(_06037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30127_ (.A1(_12064_),
    .A2(_12065_),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30128_ (.A1(_06037_),
    .A2(_06038_),
    .ZN(_06039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30129_ (.A1(_03116_),
    .A2(_06039_),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30130_ (.A1(_06036_),
    .A2(_06040_),
    .A3(_11279_),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30131_ (.I(\u0.w[2][3] ),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30132_ (.A1(_10411_),
    .A2(\text_in_r[35] ),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30133_ (.A1(_06041_),
    .A2(_06042_),
    .A3(_06043_),
    .ZN(_06044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30134_ (.A1(_03108_),
    .A2(_06039_),
    .ZN(_06045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30135_ (.A1(_03116_),
    .A2(_06035_),
    .ZN(_06046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30136_ (.A1(_06045_),
    .A2(_06046_),
    .A3(_11279_),
    .ZN(_06047_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30137_ (.A1(_10489_),
    .A2(\text_in_r[35] ),
    .Z(_06048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30138_ (.A1(_06047_),
    .A2(\u0.w[2][3] ),
    .A3(_06048_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30139_ (.A1(_06049_),
    .A2(_06044_),
    .ZN(_06050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30140_ (.A1(_06032_),
    .A2(net1199),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30141_ (.I(_16144_),
    .ZN(_06052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30142_ (.A1(_06019_),
    .A2(_06023_),
    .A3(_06052_),
    .ZN(_06053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30143_ (.A1(_06047_),
    .A2(_06042_),
    .A3(_06048_),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30144_ (.A1(_06041_),
    .A2(\u0.w[2][3] ),
    .A3(_06043_),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30145_ (.A1(_06054_),
    .A2(_06055_),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30146_ (.A1(_06053_),
    .A2(_06056_),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30147_ (.I(_06057_),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30148_ (.A1(_05978_),
    .A2(\u0.w[2][1] ),
    .A3(_05980_),
    .ZN(_06059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30149_ (.A1(_05984_),
    .A2(_05979_),
    .A3(_05985_),
    .ZN(_06060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30150_ (.A1(_06060_),
    .A2(_06059_),
    .ZN(_16138_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30151_ (.A1(_06032_),
    .A2(net24),
    .Z(_06061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30152_ (.A1(_06051_),
    .A2(_06058_),
    .B(_06061_),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30153_ (.A1(_03130_),
    .A2(_12112_),
    .ZN(_06063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30154_ (.A1(_12109_),
    .A2(_03135_),
    .ZN(_06064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30155_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_13010_),
    .ZN(_06065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30156_ (.A1(_11385_),
    .A2(\text_in_r[36] ),
    .ZN(_06066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30157_ (.A1(_06065_),
    .A2(_06066_),
    .ZN(_06067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30158_ (.A1(_06067_),
    .A2(\u0.w[2][4] ),
    .ZN(_06068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30159_ (.I(\u0.w[2][4] ),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30160_ (.A1(_06065_),
    .A2(_06069_),
    .A3(_06066_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30161_ (.A1(_06068_),
    .A2(_06070_),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30162_ (.I(_06071_),
    .Z(_06072_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30163_ (.I(_06072_),
    .Z(_06073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30164_ (.A1(_06062_),
    .A2(_06073_),
    .ZN(_06074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30165_ (.A1(net1206),
    .A2(net1184),
    .ZN(_06075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30166_ (.I(_06050_),
    .Z(_06076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30167_ (.A1(_06075_),
    .A2(_06076_),
    .Z(_06077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30168_ (.A1(_06061_),
    .A2(_06077_),
    .ZN(_06078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30169_ (.I(_16153_),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30170_ (.A1(_06025_),
    .A2(_06079_),
    .ZN(_06080_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30171_ (.I(_06056_),
    .Z(_06081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30172_ (.A1(_06080_),
    .A2(_06081_),
    .ZN(_06082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30173_ (.I(_06082_),
    .ZN(_06083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30174_ (.I(_16140_),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30175_ (.A1(_06084_),
    .A2(_06030_),
    .ZN(_06085_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30176_ (.I(_06085_),
    .Z(_06086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30177_ (.A1(_06083_),
    .A2(net23),
    .ZN(_06087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30178_ (.A1(_06067_),
    .A2(_06069_),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30179_ (.A1(_06065_),
    .A2(\u0.w[2][4] ),
    .A3(_06066_),
    .ZN(_06089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30180_ (.A1(_06088_),
    .A2(_06089_),
    .ZN(_06090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30181_ (.I(_06090_),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30182_ (.I(_06091_),
    .Z(_06092_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30183_ (.A1(_06078_),
    .A2(_06087_),
    .A3(_06092_),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30184_ (.A1(\sa31_sub[4] ),
    .A2(\sa20_sub[5] ),
    .Z(_06094_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30185_ (.A1(_06094_),
    .A2(_15180_),
    .Z(_06095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30186_ (.A1(_06094_),
    .A2(_15180_),
    .ZN(_06096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30187_ (.A1(_06095_),
    .A2(_06096_),
    .ZN(_06097_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30188_ (.A1(\sa02_sr[4] ),
    .A2(\sa12_sr[5] ),
    .ZN(_06098_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30189_ (.I(_06098_),
    .ZN(_06099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30190_ (.A1(_06097_),
    .A2(_06099_),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30191_ (.A1(_06095_),
    .A2(_06098_),
    .A3(_06096_),
    .ZN(_06101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30192_ (.A1(_06100_),
    .A2(_06101_),
    .A3(_10523_),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30193_ (.A1(_12115_),
    .A2(\text_in_r[37] ),
    .ZN(_06103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30194_ (.A1(_06102_),
    .A2(_06103_),
    .ZN(_06104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30195_ (.A1(_06104_),
    .A2(\u0.w[2][5] ),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30196_ (.I(\u0.w[2][5] ),
    .ZN(_06106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30197_ (.A1(_06102_),
    .A2(_06106_),
    .A3(_06103_),
    .ZN(_06107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30198_ (.A1(_06105_),
    .A2(_06107_),
    .ZN(_06108_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _30199_ (.I(_06108_),
    .ZN(_06109_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30200_ (.I(_06109_),
    .Z(_06110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30201_ (.A1(_06074_),
    .A2(_06093_),
    .A3(_06110_),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30202_ (.I(_06056_),
    .Z(_06112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30203_ (.A1(net24),
    .A2(_16155_),
    .B(_06112_),
    .ZN(_06113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30204_ (.A1(_06113_),
    .A2(_06061_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30205_ (.A1(_06032_),
    .A2(_06056_),
    .Z(_06115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30206_ (.A1(_06031_),
    .A2(_06079_),
    .ZN(_06116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30207_ (.A1(_06115_),
    .A2(net1195),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30208_ (.I(net1201),
    .Z(_06118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30209_ (.A1(_06114_),
    .A2(_06117_),
    .A3(_06118_),
    .ZN(_06119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30210_ (.A1(net1182),
    .A2(net1189),
    .A3(net1206),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30211_ (.A1(_06115_),
    .A2(_06120_),
    .ZN(_06121_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30212_ (.I(_16141_),
    .ZN(_06122_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _30213_ (.A1(_06122_),
    .A2(_06025_),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30214_ (.I(_06050_),
    .Z(_06124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30215_ (.A1(_06123_),
    .A2(_06124_),
    .B(net1201),
    .ZN(_06125_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _30216_ (.A1(net1202),
    .A2(_16155_),
    .ZN(_06126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30217_ (.I(_06050_),
    .Z(_06127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30218_ (.A1(_06126_),
    .A2(_06127_),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30219_ (.A1(_06121_),
    .A2(_06125_),
    .A3(_06128_),
    .ZN(_06129_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30220_ (.I(_06108_),
    .Z(_06130_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30221_ (.A1(_06119_),
    .A2(_06129_),
    .A3(_06130_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _30222_ (.A1(\sa31_sub[5] ),
    .A2(\sa20_sub[6] ),
    .A3(\sa02_sr[6] ),
    .Z(_06132_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30223_ (.A1(\sa02_sr[5] ),
    .A2(\sa12_sr[6] ),
    .Z(_06133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30224_ (.A1(_06132_),
    .A2(_06133_),
    .Z(_06134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30225_ (.A1(_06132_),
    .A2(_06133_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30226_ (.A1(_06134_),
    .A2(_12965_),
    .A3(_06135_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30227_ (.A1(_12961_),
    .A2(\text_in_r[38] ),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30228_ (.A1(_06136_),
    .A2(_06137_),
    .ZN(_06138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30229_ (.I(\u0.w[2][6] ),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30230_ (.A1(_06138_),
    .A2(_06139_),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30231_ (.A1(_06136_),
    .A2(\u0.w[2][6] ),
    .A3(_06137_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30232_ (.A1(_06140_),
    .A2(_06141_),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30233_ (.I(_06142_),
    .Z(_06143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30234_ (.A1(_06111_),
    .A2(_06131_),
    .A3(_06143_),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30235_ (.I(_16139_),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30236_ (.A1(_16162_),
    .A2(_06145_),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30237_ (.I(_06146_),
    .ZN(_06147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30238_ (.I(_16147_),
    .ZN(_06148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30239_ (.A1(_16155_),
    .A2(_06148_),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30240_ (.I(_06149_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30241_ (.I(_06081_),
    .Z(_06151_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30242_ (.A1(_06147_),
    .A2(_06150_),
    .B(_06151_),
    .ZN(_06152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30243_ (.A1(_06086_),
    .A2(_06076_),
    .Z(_06153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30244_ (.A1(_16143_),
    .A2(net1189),
    .A3(net1193),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30245_ (.A1(_06153_),
    .A2(_06154_),
    .ZN(_06155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30246_ (.A1(_06152_),
    .A2(_06155_),
    .A3(_06073_),
    .ZN(_06156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30247_ (.A1(_06031_),
    .A2(net1189),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30248_ (.A1(_06157_),
    .A2(_06076_),
    .Z(_06158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30249_ (.A1(net24),
    .A2(_16137_),
    .ZN(_06159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30250_ (.A1(_06158_),
    .A2(_06159_),
    .ZN(_06160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30251_ (.A1(net1183),
    .A2(net1185),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30252_ (.A1(net1193),
    .A2(net1189),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30253_ (.A1(_06161_),
    .A2(_06112_),
    .A3(_06162_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30254_ (.A1(_06160_),
    .A2(_06163_),
    .A3(_06118_),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30255_ (.A1(_06156_),
    .A2(_06164_),
    .A3(_06110_),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30256_ (.A1(net58),
    .A2(_16162_),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30257_ (.A1(_16155_),
    .A2(_16140_),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30258_ (.A1(_06166_),
    .A2(_06167_),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30259_ (.I(_06127_),
    .Z(_06169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30260_ (.A1(_06168_),
    .A2(_06169_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30261_ (.A1(_06084_),
    .A2(_06024_),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30262_ (.I(_06171_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30263_ (.A1(_06172_),
    .A2(_06056_),
    .Z(_06173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30264_ (.I(_06173_),
    .ZN(_06174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30265_ (.A1(_06170_),
    .A2(_06174_),
    .A3(_06118_),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30266_ (.A1(_06031_),
    .A2(_06145_),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30267_ (.A1(net1193),
    .A2(_06148_),
    .ZN(_06177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30268_ (.A1(_06176_),
    .A2(_06177_),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30269_ (.A1(_06178_),
    .A2(_06169_),
    .ZN(_06179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30270_ (.A1(_16162_),
    .A2(_16139_),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30271_ (.I(_06081_),
    .Z(_06181_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30272_ (.A1(net23),
    .A2(_06180_),
    .A3(_06181_),
    .ZN(_06182_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30273_ (.I(_06072_),
    .Z(_06183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30274_ (.A1(_06179_),
    .A2(_06182_),
    .A3(_06183_),
    .ZN(_06184_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30275_ (.I(_06108_),
    .Z(_06185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30276_ (.A1(_06175_),
    .A2(_06184_),
    .A3(_06185_),
    .ZN(_06186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30277_ (.I(_06142_),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30278_ (.I(_06187_),
    .Z(_06188_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30279_ (.A1(_06165_),
    .A2(_06186_),
    .A3(_06188_),
    .ZN(_06189_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30280_ (.A1(\sa31_sub[6] ),
    .A2(net1174),
    .Z(_06190_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _30281_ (.A1(_15233_),
    .A2(net49),
    .A3(_06190_),
    .Z(_06191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30282_ (.A1(_12961_),
    .A2(\text_in_r[39] ),
    .Z(_06192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30283_ (.A1(_06191_),
    .A2(_12965_),
    .B(_06192_),
    .ZN(_06193_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30284_ (.A1(\u0.w[2][7] ),
    .A2(_06193_),
    .Z(_06194_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30285_ (.I(_06194_),
    .Z(_06195_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30286_ (.A1(_06144_),
    .A2(_06189_),
    .A3(_06195_),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30287_ (.A1(net1193),
    .A2(net1205),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30288_ (.A1(_06157_),
    .A2(_06197_),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30289_ (.A1(_16138_),
    .A2(net1206),
    .ZN(_06199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30290_ (.I(_06199_),
    .ZN(_06200_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30291_ (.A1(_06198_),
    .A2(_06200_),
    .B(_06124_),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30292_ (.A1(_06025_),
    .A2(_16141_),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30293_ (.I(_06202_),
    .ZN(_06203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30294_ (.A1(_06203_),
    .A2(_06127_),
    .ZN(_06204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30295_ (.A1(_06162_),
    .A2(_06176_),
    .ZN(_06205_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30296_ (.I(_06056_),
    .Z(_06206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30297_ (.A1(_06205_),
    .A2(_06206_),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30298_ (.A1(_06201_),
    .A2(_06204_),
    .A3(_06207_),
    .ZN(_06208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30299_ (.A1(_16140_),
    .A2(_06025_),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30300_ (.A1(_06209_),
    .A2(_06076_),
    .Z(_06210_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30301_ (.I(_06050_),
    .Z(_06211_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30302_ (.A1(_06211_),
    .A2(_16160_),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30303_ (.A1(_06210_),
    .A2(_06212_),
    .Z(_06213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30304_ (.A1(_06213_),
    .A2(_06092_),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30305_ (.A1(_06208_),
    .A2(_06092_),
    .B(_06185_),
    .C(_06214_),
    .ZN(_06215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30306_ (.A1(net1181),
    .A2(_16147_),
    .ZN(_06216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30307_ (.A1(_06216_),
    .A2(net1199),
    .Z(_06217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30308_ (.A1(net1182),
    .A2(net1184),
    .A3(net1206),
    .ZN(_06218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30309_ (.A1(_06217_),
    .A2(_06218_),
    .Z(_06219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30310_ (.A1(_06123_),
    .A2(_06081_),
    .ZN(_06220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30311_ (.A1(_06220_),
    .A2(net1201),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30312_ (.A1(_06219_),
    .A2(_06221_),
    .Z(_06222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30313_ (.I(_16149_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30314_ (.A1(net1181),
    .A2(_06223_),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30315_ (.A1(_06224_),
    .A2(_06056_),
    .Z(_06225_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30316_ (.A1(_06225_),
    .A2(_06218_),
    .ZN(_06226_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30317_ (.I(_06108_),
    .Z(_06227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30318_ (.A1(_06226_),
    .A2(_06125_),
    .B(_06227_),
    .ZN(_06228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30319_ (.A1(_06222_),
    .A2(_06228_),
    .B(_06143_),
    .ZN(_06229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30320_ (.A1(_06215_),
    .A2(_06229_),
    .ZN(_06230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30321_ (.A1(_06085_),
    .A2(_06056_),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30322_ (.I(_06090_),
    .Z(_06232_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30323_ (.A1(_06231_),
    .A2(_06232_),
    .Z(_06233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30324_ (.A1(net1206),
    .A2(_16149_),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30325_ (.A1(_06197_),
    .A2(_06234_),
    .ZN(_06235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30326_ (.A1(_06235_),
    .A2(_06124_),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30327_ (.I(_06109_),
    .Z(_06237_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30328_ (.A1(_06233_),
    .A2(_06236_),
    .B(_06237_),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30329_ (.I(_06197_),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30330_ (.I(_06076_),
    .Z(_06240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30331_ (.A1(_06239_),
    .A2(_06240_),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30332_ (.A1(_06121_),
    .A2(_06183_),
    .A3(_06241_),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30333_ (.I(_06187_),
    .Z(_06243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30334_ (.A1(_06238_),
    .A2(_06242_),
    .B(_06243_),
    .ZN(_06244_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30335_ (.I(_06076_),
    .Z(_06245_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30336_ (.A1(_06147_),
    .A2(net1186),
    .B(_06245_),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30337_ (.I(_06091_),
    .Z(_06247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30338_ (.A1(_06246_),
    .A2(_06247_),
    .A3(_06057_),
    .ZN(_06248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30339_ (.A1(net58),
    .A2(net1206),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30340_ (.A1(_06249_),
    .A2(_06211_),
    .A3(_06209_),
    .ZN(_06250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30341_ (.A1(_06075_),
    .A2(_06216_),
    .A3(_06181_),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30342_ (.A1(_06250_),
    .A2(_06251_),
    .A3(_06183_),
    .ZN(_06252_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30343_ (.I(_06109_),
    .Z(_06253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30344_ (.A1(_06248_),
    .A2(_06252_),
    .A3(_06253_),
    .ZN(_06254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30345_ (.A1(_06244_),
    .A2(_06254_),
    .B(_06195_),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30346_ (.A1(_06230_),
    .A2(_06255_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30347_ (.A1(_06196_),
    .A2(_06256_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _30348_ (.I(_06086_),
    .ZN(_06257_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30349_ (.I(_06081_),
    .Z(_06258_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30350_ (.A1(_06257_),
    .A2(_06239_),
    .B(_06258_),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30351_ (.A1(_06205_),
    .A2(_06169_),
    .ZN(_06260_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30352_ (.A1(_06259_),
    .A2(_06092_),
    .A3(_06260_),
    .ZN(_06261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30353_ (.A1(net1202),
    .A2(net1189),
    .ZN(_06262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30354_ (.A1(_06262_),
    .A2(_06075_),
    .ZN(_06263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30355_ (.A1(_06263_),
    .A2(_06151_),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30356_ (.A1(_06075_),
    .A2(_06209_),
    .A3(_06245_),
    .ZN(_06265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30357_ (.A1(_06264_),
    .A2(_06073_),
    .A3(_06265_),
    .ZN(_06266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30358_ (.A1(_06261_),
    .A2(_06266_),
    .A3(_06130_),
    .ZN(_06267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30359_ (.A1(_06199_),
    .A2(_06075_),
    .ZN(_06268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30360_ (.A1(_06268_),
    .A2(_06169_),
    .ZN(_06269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30361_ (.A1(_06199_),
    .A2(_06181_),
    .A3(_06080_),
    .ZN(_06270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30362_ (.A1(_06269_),
    .A2(_06270_),
    .A3(_06247_),
    .ZN(_06271_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30363_ (.A1(_06154_),
    .A2(_06181_),
    .A3(_06167_),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30364_ (.A1(_16155_),
    .A2(net1208),
    .ZN(_06273_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30365_ (.I(_06273_),
    .ZN(_06274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30366_ (.A1(_06274_),
    .A2(_06240_),
    .B(_06232_),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30367_ (.A1(_06272_),
    .A2(_06275_),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30368_ (.A1(_06271_),
    .A2(_06276_),
    .A3(_06253_),
    .ZN(_06277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30369_ (.A1(_06267_),
    .A2(_06277_),
    .A3(_06143_),
    .ZN(_06278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30370_ (.A1(_06249_),
    .A2(_06159_),
    .A3(_06211_),
    .ZN(_06279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30371_ (.A1(_06161_),
    .A2(_16162_),
    .A3(_06112_),
    .ZN(_06280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30372_ (.A1(_06279_),
    .A2(_06280_),
    .A3(_06073_),
    .ZN(_06281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30373_ (.A1(_06032_),
    .A2(net23),
    .A3(_06258_),
    .ZN(_06282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30374_ (.A1(_06162_),
    .A2(_06240_),
    .A3(net1191),
    .ZN(_06283_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30375_ (.A1(_06282_),
    .A2(_06283_),
    .A3(_06247_),
    .ZN(_06284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30376_ (.A1(_06281_),
    .A2(_06284_),
    .A3(_06253_),
    .ZN(_06285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30377_ (.A1(net58),
    .A2(_16162_),
    .B(_06127_),
    .ZN(_06286_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30378_ (.A1(_06286_),
    .A2(_06200_),
    .ZN(_06287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30379_ (.A1(_06239_),
    .A2(_06124_),
    .B(_06072_),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30380_ (.A1(_06287_),
    .A2(_06288_),
    .B(_06237_),
    .ZN(_06289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30381_ (.A1(_06171_),
    .A2(_06081_),
    .Z(_06290_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _30382_ (.I(_06091_),
    .Z(_06291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30383_ (.A1(_06290_),
    .A2(net1195),
    .B(_06291_),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30384_ (.A1(_06292_),
    .A2(_06201_),
    .ZN(_06293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30385_ (.A1(_06289_),
    .A2(_06293_),
    .ZN(_06294_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30386_ (.A1(_06285_),
    .A2(_06294_),
    .A3(_06188_),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30387_ (.A1(_06278_),
    .A2(_06295_),
    .B(_06195_),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30388_ (.A1(_06077_),
    .A2(_06180_),
    .ZN(_06297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30389_ (.A1(_06109_),
    .A2(_06232_),
    .Z(_06298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30390_ (.A1(_06081_),
    .A2(_16155_),
    .ZN(_06299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30391_ (.I(_06299_),
    .ZN(_06300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30392_ (.A1(_06300_),
    .A2(_06262_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _30393_ (.A1(_06280_),
    .A2(_06297_),
    .A3(_06298_),
    .A4(_06301_),
    .ZN(_06302_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30394_ (.I(_16163_),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _30395_ (.A1(_06108_),
    .A2(_06303_),
    .A3(_06206_),
    .Z(_06304_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30396_ (.A1(_06304_),
    .A2(_06291_),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30397_ (.A1(_06217_),
    .A2(_06120_),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30398_ (.A1(_06305_),
    .A2(_06306_),
    .B(_06143_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30399_ (.A1(_06302_),
    .A2(_06307_),
    .ZN(_06308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30400_ (.A1(_06158_),
    .A2(_06166_),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30401_ (.A1(net24),
    .A2(net1181),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30402_ (.A1(_06058_),
    .A2(_06310_),
    .ZN(_06311_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _30403_ (.A1(_06309_),
    .A2(_06247_),
    .A3(_06311_),
    .A4(_06227_),
    .Z(_06312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30404_ (.A1(_06308_),
    .A2(_06312_),
    .B(_06195_),
    .ZN(_06313_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _30405_ (.I(_06176_),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30406_ (.A1(_06314_),
    .A2(_06206_),
    .ZN(_06315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30407_ (.A1(_06123_),
    .A2(_06127_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30408_ (.A1(_06315_),
    .A2(_06316_),
    .Z(_06317_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30409_ (.I(_06162_),
    .ZN(_06318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30410_ (.A1(_06318_),
    .A2(_06245_),
    .B(net1209),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30411_ (.I(_06209_),
    .ZN(_06320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30412_ (.A1(_06320_),
    .A2(_06081_),
    .Z(_06321_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30413_ (.I(_06321_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30414_ (.A1(_06317_),
    .A2(_06319_),
    .A3(_06322_),
    .ZN(_06323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30415_ (.A1(_06158_),
    .A2(_06180_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30416_ (.A1(_06324_),
    .A2(_06183_),
    .A3(_06311_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30417_ (.A1(_06323_),
    .A2(_06325_),
    .A3(_06253_),
    .ZN(_06326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30418_ (.A1(_06051_),
    .A2(_06120_),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30419_ (.A1(_06231_),
    .A2(_06072_),
    .Z(_06328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30420_ (.A1(_06327_),
    .A2(_06328_),
    .B(_06237_),
    .ZN(_06329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30421_ (.A1(_06116_),
    .A2(_06050_),
    .Z(_06330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30422_ (.A1(_06025_),
    .A2(_06122_),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30423_ (.A1(_06330_),
    .A2(_06331_),
    .ZN(_06332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30424_ (.A1(_06272_),
    .A2(_06247_),
    .A3(_06332_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30425_ (.A1(_06329_),
    .A2(_06333_),
    .ZN(_06334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30426_ (.A1(_06326_),
    .A2(_06334_),
    .B(_06243_),
    .ZN(_06335_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30427_ (.A1(_06313_),
    .A2(_06335_),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30428_ (.A1(_06336_),
    .A2(_06296_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30429_ (.A1(_06161_),
    .A2(_06249_),
    .A3(_06206_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30430_ (.A1(net1199),
    .A2(_06053_),
    .Z(_06338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30431_ (.A1(_06338_),
    .A2(_06080_),
    .ZN(_06339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30432_ (.A1(_06337_),
    .A2(_06339_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30433_ (.I(_06091_),
    .Z(_06341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30434_ (.A1(_06340_),
    .A2(_06341_),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30435_ (.A1(_06161_),
    .A2(_16155_),
    .ZN(_06343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30436_ (.A1(_06197_),
    .A2(_06056_),
    .Z(_06344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30437_ (.A1(_06343_),
    .A2(_06344_),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30438_ (.I(_06071_),
    .Z(_06346_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30439_ (.A1(_06345_),
    .A2(_06346_),
    .A3(_06250_),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30440_ (.A1(_06342_),
    .A2(_06347_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30441_ (.A1(_06348_),
    .A2(_06130_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30442_ (.A1(_06154_),
    .A2(_06151_),
    .A3(net1196),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30443_ (.A1(_06061_),
    .A2(_06127_),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30444_ (.A1(_06350_),
    .A2(_06351_),
    .A3(_06073_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30445_ (.A1(_06166_),
    .A2(_06240_),
    .A3(net23),
    .ZN(_06353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30446_ (.A1(_06157_),
    .A2(_06202_),
    .ZN(_06354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30447_ (.A1(_06354_),
    .A2(_06151_),
    .ZN(_06355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30448_ (.A1(_06353_),
    .A2(_06355_),
    .A3(_06247_),
    .ZN(_06356_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30449_ (.A1(_06352_),
    .A2(_06110_),
    .A3(_06356_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30450_ (.A1(_06349_),
    .A2(_06357_),
    .A3(_06188_),
    .ZN(_06358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30451_ (.A1(_06075_),
    .A2(_06224_),
    .A3(_06211_),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30452_ (.A1(_06086_),
    .A2(_06209_),
    .A3(_06112_),
    .ZN(_06360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30453_ (.A1(_06360_),
    .A2(_06359_),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30454_ (.A1(_06361_),
    .A2(_06346_),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30455_ (.A1(_06310_),
    .A2(_06112_),
    .A3(_06234_),
    .ZN(_06363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30456_ (.A1(_16162_),
    .A2(_16153_),
    .ZN(_06364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30457_ (.A1(_06157_),
    .A2(_06364_),
    .A3(_06124_),
    .ZN(_06365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30458_ (.A1(_06363_),
    .A2(_06365_),
    .A3(_06291_),
    .ZN(_06366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30459_ (.A1(_06362_),
    .A2(_06366_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30460_ (.A1(_06367_),
    .A2(_06110_),
    .ZN(_06368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30461_ (.A1(_06198_),
    .A2(_06151_),
    .ZN(_06369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30462_ (.A1(_06364_),
    .A2(_06234_),
    .ZN(_06370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30463_ (.A1(_06370_),
    .A2(_06169_),
    .ZN(_06371_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30464_ (.A1(_06369_),
    .A2(_06371_),
    .A3(_06118_),
    .ZN(_06372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30465_ (.A1(_16162_),
    .A2(_06052_),
    .ZN(_06373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30466_ (.A1(_06199_),
    .A2(_06258_),
    .A3(_06373_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30467_ (.A1(_06374_),
    .A2(_06236_),
    .A3(_06183_),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30468_ (.A1(_06372_),
    .A2(_06375_),
    .A3(_06185_),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30469_ (.A1(_06368_),
    .A2(_06376_),
    .A3(_06143_),
    .ZN(_06377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30470_ (.A1(_06358_),
    .A2(_06377_),
    .A3(_06195_),
    .ZN(_06378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30471_ (.A1(_06310_),
    .A2(_06032_),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30472_ (.A1(_06122_),
    .A2(_06052_),
    .Z(_06380_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30473_ (.A1(_16162_),
    .A2(_06380_),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30474_ (.A1(_06379_),
    .A2(_06381_),
    .B(_06151_),
    .ZN(_06382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30475_ (.A1(_06382_),
    .A2(_06092_),
    .A3(_06306_),
    .ZN(_06383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30476_ (.A1(_06314_),
    .A2(_06127_),
    .ZN(_06384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30477_ (.I(_06071_),
    .Z(_06385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30478_ (.A1(_06384_),
    .A2(_06385_),
    .Z(_06386_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30479_ (.I(_06231_),
    .ZN(_06387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30480_ (.A1(_06387_),
    .A2(_06373_),
    .ZN(_06388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30481_ (.A1(_06386_),
    .A2(_06388_),
    .B(_06227_),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30482_ (.A1(_06383_),
    .A2(_06389_),
    .ZN(_06390_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30483_ (.A1(_06076_),
    .A2(_16158_),
    .Z(_06391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30484_ (.A1(_06351_),
    .A2(_06391_),
    .ZN(_06392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30485_ (.A1(_06392_),
    .A2(_06341_),
    .Z(_06393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30486_ (.A1(_16167_),
    .A2(_06240_),
    .B(_06385_),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30487_ (.A1(_06337_),
    .A2(_06394_),
    .B(_06237_),
    .ZN(_06395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30488_ (.A1(_06393_),
    .A2(_06395_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30489_ (.A1(_06390_),
    .A2(_06396_),
    .A3(_06188_),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30490_ (.A1(_06149_),
    .A2(_06081_),
    .Z(_06398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30491_ (.A1(_06398_),
    .A2(_06209_),
    .Z(_06399_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _30492_ (.A1(_06249_),
    .A2(_06124_),
    .A3(_06146_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30493_ (.A1(_06399_),
    .A2(_06400_),
    .B(_06118_),
    .ZN(_06401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30494_ (.A1(_06249_),
    .A2(_06159_),
    .A3(_06081_),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30495_ (.A1(_06402_),
    .A2(net1209),
    .Z(_06403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30496_ (.A1(_06169_),
    .A2(net1197),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30497_ (.A1(_06403_),
    .A2(_06404_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30498_ (.A1(_06401_),
    .A2(_06405_),
    .A3(_06130_),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30499_ (.A1(_06290_),
    .A2(_06218_),
    .ZN(_06407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30500_ (.A1(_16160_),
    .A2(_06245_),
    .B(_06232_),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30501_ (.A1(_06407_),
    .A2(_06408_),
    .B(_06108_),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30502_ (.A1(_06310_),
    .A2(_06112_),
    .A3(_06075_),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30503_ (.A1(_06250_),
    .A2(_06410_),
    .A3(_06341_),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30504_ (.A1(_06409_),
    .A2(_06411_),
    .B(_06187_),
    .ZN(_06412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30505_ (.A1(_06406_),
    .A2(_06412_),
    .ZN(_06413_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30506_ (.I(_06194_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30507_ (.A1(_06397_),
    .A2(_06413_),
    .A3(_06414_),
    .ZN(_06415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30508_ (.A1(_06378_),
    .A2(_06415_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30509_ (.A1(_06217_),
    .A2(_06249_),
    .Z(_06416_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30510_ (.A1(_06416_),
    .A2(_06173_),
    .B(_06108_),
    .ZN(_06417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30511_ (.A1(_06257_),
    .A2(_06127_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30512_ (.I(_06418_),
    .ZN(_06419_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30513_ (.A1(_06419_),
    .A2(_06237_),
    .B(_06221_),
    .ZN(_06420_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30514_ (.A1(_06417_),
    .A2(_06420_),
    .B(_06143_),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30515_ (.A1(_06380_),
    .A2(_16155_),
    .B(net1200),
    .ZN(_06422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30516_ (.A1(_06422_),
    .A2(_06080_),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30517_ (.A1(_06051_),
    .A2(_06086_),
    .ZN(_06424_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30518_ (.A1(_06423_),
    .A2(_06424_),
    .A3(_06108_),
    .ZN(_06425_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30519_ (.A1(_06234_),
    .A2(_06076_),
    .Z(_06426_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30520_ (.A1(_06359_),
    .A2(_06109_),
    .A3(_06426_),
    .ZN(_06427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30521_ (.A1(_06425_),
    .A2(_06427_),
    .ZN(_06428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30522_ (.A1(_06428_),
    .A2(_06073_),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30523_ (.A1(_06429_),
    .A2(_06421_),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30524_ (.A1(_06279_),
    .A2(_06207_),
    .A3(_06385_),
    .ZN(_06431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30525_ (.A1(_06032_),
    .A2(_06234_),
    .ZN(_06432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30526_ (.A1(_06432_),
    .A2(_06206_),
    .ZN(_06433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30527_ (.A1(_06080_),
    .A2(_06086_),
    .A3(_06211_),
    .ZN(_06434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30528_ (.A1(_06433_),
    .A2(_06434_),
    .A3(_06232_),
    .ZN(_06435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30529_ (.A1(_06431_),
    .A2(_06435_),
    .ZN(_06436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30530_ (.A1(_06436_),
    .A2(_06253_),
    .ZN(_06437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30531_ (.A1(_06422_),
    .A2(_06224_),
    .ZN(_06438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30532_ (.A1(_06438_),
    .A2(_06306_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30533_ (.A1(_06439_),
    .A2(_06346_),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30534_ (.A1(_06365_),
    .A2(_06291_),
    .B(_06109_),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30535_ (.A1(_06440_),
    .A2(_06441_),
    .ZN(_06442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30536_ (.A1(_06437_),
    .A2(_06143_),
    .A3(_06442_),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30537_ (.A1(_06430_),
    .A2(_06443_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30538_ (.A1(_06444_),
    .A2(_06195_),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30539_ (.A1(_06309_),
    .A2(_06174_),
    .ZN(_06446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30540_ (.A1(_06446_),
    .A2(_06092_),
    .ZN(_06447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30541_ (.A1(_06158_),
    .A2(_06161_),
    .ZN(_06448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30542_ (.A1(_06168_),
    .A2(_06151_),
    .ZN(_06449_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30543_ (.A1(_06448_),
    .A2(_06449_),
    .A3(_06183_),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30544_ (.A1(_06447_),
    .A2(_06450_),
    .A3(_06130_),
    .ZN(_06451_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30545_ (.A1(_06314_),
    .A2(_06172_),
    .B(_06258_),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30546_ (.A1(_06318_),
    .A2(_06150_),
    .B(_06245_),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30547_ (.A1(_06452_),
    .A2(_06453_),
    .A3(_06247_),
    .ZN(_06454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30548_ (.A1(_06167_),
    .A2(_06076_),
    .Z(_06455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30549_ (.A1(_06455_),
    .A2(_06310_),
    .ZN(_06456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30550_ (.A1(net1195),
    .A2(_06373_),
    .A3(_06181_),
    .ZN(_06457_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30551_ (.A1(_06456_),
    .A2(_06183_),
    .A3(_06457_),
    .ZN(_06458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30552_ (.A1(_06454_),
    .A2(_06458_),
    .A3(_06253_),
    .ZN(_06459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30553_ (.A1(_06451_),
    .A2(_06459_),
    .A3(_06188_),
    .ZN(_06460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30554_ (.A1(_06398_),
    .A2(_06310_),
    .A3(_06162_),
    .ZN(_06461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30555_ (.I(_06268_),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30556_ (.A1(_06462_),
    .A2(_06210_),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30557_ (.A1(_06461_),
    .A2(_06463_),
    .A3(_06346_),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30558_ (.A1(_06153_),
    .A2(_06177_),
    .ZN(_06465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30559_ (.A1(_06465_),
    .A2(_06163_),
    .A3(_06341_),
    .ZN(_06466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30560_ (.A1(_06464_),
    .A2(_06466_),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30561_ (.A1(_06467_),
    .A2(_06110_),
    .ZN(_06468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30562_ (.A1(_06455_),
    .A2(_06224_),
    .ZN(_06469_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30563_ (.A1(_06469_),
    .A2(_06270_),
    .A3(_06247_),
    .ZN(_06470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30564_ (.A1(_06299_),
    .A2(net1209),
    .Z(_06471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30565_ (.A1(_06161_),
    .A2(_06157_),
    .ZN(_06472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30566_ (.A1(_06471_),
    .A2(_06472_),
    .B(_06237_),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30567_ (.A1(_06470_),
    .A2(_06473_),
    .B(_06187_),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30568_ (.A1(_06468_),
    .A2(_06474_),
    .ZN(_06475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30569_ (.A1(_06460_),
    .A2(_06475_),
    .A3(_06414_),
    .ZN(_06476_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30570_ (.A1(_06445_),
    .A2(_06476_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _30571_ (.A1(_06225_),
    .A2(_06385_),
    .A3(net1186),
    .ZN(_06477_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30572_ (.A1(_06477_),
    .A2(_06185_),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30573_ (.A1(_06286_),
    .A2(_06075_),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30574_ (.A1(_06479_),
    .A2(_06297_),
    .A3(_06073_),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30575_ (.A1(_06478_),
    .A2(_06480_),
    .B(_06243_),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30576_ (.A1(_06403_),
    .A2(_06309_),
    .ZN(_06482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30577_ (.A1(_06199_),
    .A2(_06206_),
    .Z(_06483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30578_ (.A1(_06483_),
    .A2(_06180_),
    .ZN(_06484_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30579_ (.A1(_06199_),
    .A2(_06262_),
    .A3(_06124_),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30580_ (.A1(_06484_),
    .A2(_06092_),
    .A3(_06485_),
    .ZN(_06486_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30581_ (.A1(_06482_),
    .A2(_06486_),
    .A3(_06130_),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30582_ (.A1(_06481_),
    .A2(_06487_),
    .B(_06195_),
    .ZN(_06488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30583_ (.A1(_06218_),
    .A2(_06206_),
    .ZN(_06489_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30584_ (.A1(_06126_),
    .A2(_06489_),
    .B(_06339_),
    .C(_06247_),
    .ZN(_06490_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30585_ (.A1(_06315_),
    .A2(_06072_),
    .Z(_06491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30586_ (.A1(net58),
    .A2(_06206_),
    .ZN(_06492_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30587_ (.A1(_06492_),
    .A2(_16155_),
    .Z(_06493_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30588_ (.A1(_06201_),
    .A2(_06491_),
    .A3(_06493_),
    .ZN(_06494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30589_ (.A1(_06490_),
    .A2(_06494_),
    .A3(_06130_),
    .ZN(_06495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30590_ (.A1(_06426_),
    .A2(_06232_),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30591_ (.A1(_06496_),
    .A2(_06236_),
    .A3(_06322_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30592_ (.A1(_06330_),
    .A2(_06171_),
    .ZN(_06498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30593_ (.A1(_06226_),
    .A2(_06498_),
    .A3(_06073_),
    .ZN(_06499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30594_ (.A1(_06497_),
    .A2(_06499_),
    .A3(_06110_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30595_ (.A1(_06495_),
    .A2(_06500_),
    .A3(_06188_),
    .ZN(_06501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30596_ (.A1(_06488_),
    .A2(_06501_),
    .ZN(_06502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30597_ (.A1(_06225_),
    .A2(_06157_),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30598_ (.A1(_06161_),
    .A2(_06310_),
    .A3(_06240_),
    .ZN(_06504_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30599_ (.A1(_06503_),
    .A2(_06504_),
    .A3(_06118_),
    .ZN(_06505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30600_ (.A1(_06246_),
    .A2(_06163_),
    .A3(_06183_),
    .ZN(_06506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30601_ (.A1(_06505_),
    .A2(_06506_),
    .A3(_06130_),
    .ZN(_06507_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30602_ (.I(_16151_),
    .ZN(_06508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30603_ (.A1(_06211_),
    .A2(_06508_),
    .ZN(_06509_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30604_ (.A1(_06124_),
    .A2(_06320_),
    .B(_06509_),
    .C(net1209),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30605_ (.A1(_06510_),
    .A2(_06237_),
    .ZN(_06511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30606_ (.I(_06511_),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30607_ (.A1(_06343_),
    .A2(_06112_),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30608_ (.A1(_06225_),
    .A2(_06199_),
    .ZN(_06514_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30609_ (.A1(_06513_),
    .A2(_06514_),
    .A3(_06118_),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30610_ (.A1(_06512_),
    .A2(_06515_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30611_ (.A1(_06507_),
    .A2(_06516_),
    .A3(_06188_),
    .ZN(_06517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30612_ (.A1(_06121_),
    .A2(_06385_),
    .Z(_06518_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30613_ (.A1(_06338_),
    .A2(_06209_),
    .Z(_06519_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30614_ (.I(_06519_),
    .ZN(_06520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30615_ (.A1(_06520_),
    .A2(_06518_),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30616_ (.A1(_06331_),
    .A2(_06127_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30617_ (.A1(_06522_),
    .A2(_06232_),
    .Z(_06523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30618_ (.A1(_06154_),
    .A2(_06151_),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30619_ (.A1(_06523_),
    .A2(_06524_),
    .B(_06227_),
    .ZN(_06525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30620_ (.A1(_06521_),
    .A2(_06525_),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30621_ (.A1(_06158_),
    .A2(_06080_),
    .ZN(_06527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30622_ (.A1(_16162_),
    .A2(_06181_),
    .B(_06232_),
    .ZN(_06528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30623_ (.A1(_06527_),
    .A2(_06528_),
    .B(_06237_),
    .ZN(_06529_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30624_ (.A1(_06057_),
    .A2(_06126_),
    .B(net1201),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30625_ (.A1(_06128_),
    .A2(_06384_),
    .ZN(_06531_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30626_ (.A1(_06530_),
    .A2(_06531_),
    .Z(_06532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30627_ (.A1(_06529_),
    .A2(_06532_),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30628_ (.A1(_06143_),
    .A2(_06533_),
    .A3(_06526_),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30629_ (.A1(_06517_),
    .A2(_06534_),
    .A3(_06195_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30630_ (.A1(_06535_),
    .A2(_06502_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30631_ (.I(_06249_),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30632_ (.A1(_06522_),
    .A2(_06536_),
    .ZN(_06537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30633_ (.A1(_06537_),
    .A2(_06321_),
    .B(_06291_),
    .ZN(_06538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30634_ (.A1(_06387_),
    .A2(_06146_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30635_ (.A1(_06124_),
    .A2(_06364_),
    .B(net1201),
    .ZN(_06540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30636_ (.A1(_06539_),
    .A2(_06540_),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30637_ (.A1(_06538_),
    .A2(_06185_),
    .A3(_06541_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30638_ (.A1(_06542_),
    .A2(_06243_),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30639_ (.A1(_06051_),
    .A2(_06262_),
    .ZN(_06544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30640_ (.A1(_06544_),
    .A2(_06291_),
    .ZN(_06545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30641_ (.A1(_06120_),
    .A2(_06216_),
    .B(_06245_),
    .ZN(_06546_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30642_ (.A1(_06545_),
    .A2(_06546_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30643_ (.A1(_06485_),
    .A2(_06492_),
    .B(_06341_),
    .ZN(_06548_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _30644_ (.A1(_06547_),
    .A2(_06548_),
    .A3(_06185_),
    .ZN(_06549_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30645_ (.A1(_06543_),
    .A2(_06549_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30646_ (.A1(_06224_),
    .A2(_06127_),
    .Z(_06551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30647_ (.A1(_06551_),
    .A2(_06218_),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30648_ (.A1(_06123_),
    .A2(net1207),
    .B(_06181_),
    .ZN(_06553_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30649_ (.A1(_06552_),
    .A2(_06247_),
    .A3(_06553_),
    .ZN(_06554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30650_ (.A1(_06080_),
    .A2(net1191),
    .A3(_06181_),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30651_ (.A1(_06125_),
    .A2(_06128_),
    .A3(_06555_),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30652_ (.A1(_06554_),
    .A2(_06556_),
    .A3(_06253_),
    .ZN(_06557_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30653_ (.A1(_06153_),
    .A2(_06291_),
    .ZN(_06558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30654_ (.A1(_06433_),
    .A2(_06558_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30655_ (.A1(_06338_),
    .A2(_06346_),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30656_ (.A1(_06560_),
    .A2(_06280_),
    .ZN(_06561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30657_ (.A1(_06559_),
    .A2(_06561_),
    .A3(_06185_),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30658_ (.A1(_06562_),
    .A2(_06557_),
    .B(_06243_),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30659_ (.A1(_06563_),
    .A2(_06550_),
    .B(_06414_),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30660_ (.A1(net1189),
    .A2(_06258_),
    .B(_06232_),
    .ZN(_06565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30661_ (.A1(_06160_),
    .A2(_06565_),
    .B(_06227_),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30662_ (.A1(_06061_),
    .A2(_06387_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30663_ (.A1(_06551_),
    .A2(_06199_),
    .ZN(_06568_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30664_ (.A1(_06567_),
    .A2(_06568_),
    .A3(_06118_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30665_ (.A1(_06566_),
    .A2(_06569_),
    .B(_06243_),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30666_ (.A1(_06198_),
    .A2(_06169_),
    .ZN(_06571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30667_ (.A1(_06518_),
    .A2(_06571_),
    .ZN(_06572_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30668_ (.A1(_06120_),
    .A2(_06169_),
    .A3(_06080_),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30669_ (.I(_06177_),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30670_ (.A1(_06574_),
    .A2(_06258_),
    .B(_06385_),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30671_ (.A1(_06573_),
    .A2(_06575_),
    .B(_06253_),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30672_ (.A1(_06572_),
    .A2(_06576_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30673_ (.A1(_06570_),
    .A2(_06577_),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30674_ (.A1(_06455_),
    .A2(_06080_),
    .ZN(_06579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30675_ (.A1(_06387_),
    .A2(_06216_),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30676_ (.A1(_06579_),
    .A2(_06580_),
    .A3(_06092_),
    .ZN(_06581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30677_ (.A1(_06148_),
    .A2(_06258_),
    .B(_06232_),
    .ZN(_06582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30678_ (.A1(_06120_),
    .A2(_06169_),
    .ZN(_06583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30679_ (.A1(_06582_),
    .A2(_06583_),
    .B(_06237_),
    .ZN(_06584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30680_ (.A1(_06581_),
    .A2(_06584_),
    .ZN(_06585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30681_ (.A1(_06288_),
    .A2(_06082_),
    .B(_06227_),
    .ZN(_06586_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30682_ (.A1(_06061_),
    .A2(_06120_),
    .A3(_06240_),
    .ZN(_06587_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30683_ (.A1(_06422_),
    .A2(_06291_),
    .ZN(_06588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30684_ (.A1(_06587_),
    .A2(_06588_),
    .ZN(_06589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30685_ (.A1(_06586_),
    .A2(_06589_),
    .ZN(_06590_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30686_ (.A1(_06585_),
    .A2(_06590_),
    .A3(_06188_),
    .ZN(_06591_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30687_ (.A1(_06578_),
    .A2(_06591_),
    .A3(_06195_),
    .ZN(_06592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30688_ (.A1(_06564_),
    .A2(_06592_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30689_ (.I(_06217_),
    .ZN(_06593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30690_ (.A1(_06514_),
    .A2(_06593_),
    .ZN(_06594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30691_ (.A1(_06594_),
    .A2(_06341_),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30692_ (.A1(_06345_),
    .A2(_06346_),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30693_ (.A1(_06595_),
    .A2(_06596_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30694_ (.A1(_06597_),
    .A2(_06130_),
    .ZN(_06598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30695_ (.A1(_06083_),
    .A2(_06167_),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30696_ (.A1(_06319_),
    .A2(_06599_),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30697_ (.I(_16157_),
    .ZN(_06601_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30698_ (.A1(_06601_),
    .A2(_06258_),
    .B(_06291_),
    .ZN(_06602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30699_ (.A1(_06568_),
    .A2(_06602_),
    .ZN(_06603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30700_ (.A1(_06600_),
    .A2(_06603_),
    .A3(_06110_),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30701_ (.A1(_06598_),
    .A2(_06188_),
    .A3(_06604_),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30702_ (.A1(net58),
    .A2(_06151_),
    .B(_06472_),
    .C(_06183_),
    .ZN(_06606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30703_ (.A1(_06472_),
    .A2(_06151_),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30704_ (.A1(_06330_),
    .A2(_06162_),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30705_ (.A1(_06607_),
    .A2(_06608_),
    .A3(_06118_),
    .ZN(_06609_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30706_ (.A1(_06606_),
    .A2(_06609_),
    .A3(_06110_),
    .ZN(_06610_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30707_ (.A1(_06167_),
    .A2(_06112_),
    .Z(_06611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30708_ (.A1(_06433_),
    .A2(_06073_),
    .A3(_06611_),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30709_ (.A1(_06286_),
    .A2(_06346_),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30710_ (.A1(_06613_),
    .A2(_06078_),
    .ZN(_06614_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30711_ (.A1(_06612_),
    .A2(_06614_),
    .A3(_06185_),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30712_ (.A1(_06610_),
    .A2(_06143_),
    .A3(_06615_),
    .ZN(_06616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30713_ (.A1(_06605_),
    .A2(_06616_),
    .A3(_06195_),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30714_ (.A1(_06203_),
    .A2(_06112_),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30715_ (.A1(_06384_),
    .A2(_06618_),
    .Z(_06619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30716_ (.A1(_06496_),
    .A2(_06619_),
    .B(_06227_),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30717_ (.A1(_06310_),
    .A2(_06206_),
    .Z(_06621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30718_ (.A1(_06621_),
    .A2(_06161_),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30719_ (.A1(_16156_),
    .A2(_16165_),
    .B(_06245_),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30720_ (.A1(_06622_),
    .A2(_06073_),
    .A3(_06623_),
    .ZN(_06624_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30721_ (.A1(_06620_),
    .A2(_06624_),
    .B(_06243_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30722_ (.A1(_06379_),
    .A2(_06112_),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30723_ (.A1(_06626_),
    .A2(_06220_),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30724_ (.A1(_06330_),
    .A2(_06224_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30725_ (.A1(_06628_),
    .A2(_06385_),
    .Z(_06629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30726_ (.A1(_06627_),
    .A2(_06629_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30727_ (.A1(_06235_),
    .A2(_06203_),
    .B(_06258_),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30728_ (.A1(_06210_),
    .A2(_06157_),
    .ZN(_06632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30729_ (.A1(_06631_),
    .A2(_06118_),
    .A3(_06632_),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30730_ (.A1(_06630_),
    .A2(_06633_),
    .A3(_06130_),
    .ZN(_06634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30731_ (.A1(_06625_),
    .A2(_06634_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30732_ (.A1(_06316_),
    .A2(net1209),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30733_ (.A1(_06519_),
    .A2(_06636_),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30734_ (.A1(_06489_),
    .A2(_06318_),
    .Z(_06638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30735_ (.A1(_06638_),
    .A2(_06637_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30736_ (.A1(_06574_),
    .A2(_06245_),
    .B(_06385_),
    .ZN(_06640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30737_ (.A1(_06157_),
    .A2(net58),
    .ZN(_06641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30738_ (.A1(_06641_),
    .A2(_06258_),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30739_ (.A1(_06640_),
    .A2(_06642_),
    .B(_06237_),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30740_ (.A1(_06643_),
    .A2(_06639_),
    .B(_06143_),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30741_ (.A1(_06392_),
    .A2(_06418_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30742_ (.A1(_06645_),
    .A2(_06092_),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30743_ (.A1(net23),
    .A2(_06202_),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30744_ (.A1(_06647_),
    .A2(_06240_),
    .B(_06291_),
    .ZN(_06648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30745_ (.A1(_06483_),
    .A2(_06061_),
    .ZN(_06649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30746_ (.A1(_06648_),
    .A2(_06649_),
    .B(_06227_),
    .ZN(_06650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30747_ (.A1(_06646_),
    .A2(_06650_),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30748_ (.A1(_06651_),
    .A2(_06644_),
    .ZN(_06652_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30749_ (.A1(_06652_),
    .A2(_06635_),
    .A3(_06414_),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30750_ (.A1(_06653_),
    .A2(_06617_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30751_ (.A1(_06199_),
    .A2(_06032_),
    .A3(_06211_),
    .ZN(_06654_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30752_ (.A1(_06167_),
    .A2(_06171_),
    .A3(_06206_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30753_ (.A1(_06654_),
    .A2(_06655_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30754_ (.A1(_06656_),
    .A2(_06341_),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30755_ (.A1(_06171_),
    .A2(_06234_),
    .A3(_06124_),
    .ZN(_06658_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30756_ (.A1(_06211_),
    .A2(_16165_),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30757_ (.A1(_06658_),
    .A2(_06346_),
    .A3(_06659_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30758_ (.A1(_06657_),
    .A2(_06185_),
    .A3(_06660_),
    .ZN(_06661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30759_ (.A1(_06641_),
    .A2(_06211_),
    .Z(_06662_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30760_ (.A1(_06076_),
    .A2(_16151_),
    .ZN(_06663_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30761_ (.A1(_06663_),
    .A2(_06091_),
    .ZN(_06664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30762_ (.A1(_06664_),
    .A2(_06204_),
    .ZN(_06665_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30763_ (.A1(_06530_),
    .A2(_06662_),
    .B(_06665_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30764_ (.A1(_06666_),
    .A2(_06253_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30765_ (.A1(_06661_),
    .A2(_06667_),
    .A3(_06243_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30766_ (.A1(_06668_),
    .A2(_06414_),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30767_ (.A1(_06249_),
    .A2(_06262_),
    .A3(_06245_),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30768_ (.A1(_06438_),
    .A2(_06670_),
    .B(_06346_),
    .ZN(_06671_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30769_ (.A1(_06231_),
    .A2(_06574_),
    .B(_06385_),
    .ZN(_06672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30770_ (.A1(_06176_),
    .A2(_06211_),
    .ZN(_06673_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30771_ (.A1(_06379_),
    .A2(_06673_),
    .ZN(_06674_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30772_ (.A1(_06672_),
    .A2(_06674_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30773_ (.A1(_06671_),
    .A2(_06675_),
    .B(_06110_),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30774_ (.A1(net1187),
    .A2(_06240_),
    .B(_06385_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30775_ (.A1(_06622_),
    .A2(_06677_),
    .B(_06253_),
    .ZN(_06678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30776_ (.A1(_06169_),
    .A2(_06126_),
    .B(_06673_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30777_ (.A1(_06679_),
    .A2(_06491_),
    .A3(_06204_),
    .ZN(_06680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30778_ (.A1(_06678_),
    .A2(_06680_),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30779_ (.A1(_06676_),
    .A2(_06681_),
    .B(_06243_),
    .ZN(_06682_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30780_ (.A1(_06669_),
    .A2(_06682_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30781_ (.A1(_06113_),
    .A2(_06154_),
    .ZN(_06684_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30782_ (.A1(_06684_),
    .A2(_06402_),
    .A3(_06183_),
    .ZN(_06685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30783_ (.A1(_06310_),
    .A2(_06181_),
    .A3(_06157_),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30784_ (.A1(_06240_),
    .A2(net1189),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30785_ (.A1(_06686_),
    .A2(_06341_),
    .A3(_06687_),
    .ZN(_06688_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30786_ (.A1(_06685_),
    .A2(_06110_),
    .A3(_06688_),
    .ZN(_06689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30787_ (.A1(_06455_),
    .A2(_06154_),
    .ZN(_06690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30788_ (.A1(_06690_),
    .A2(_06489_),
    .A3(_06341_),
    .ZN(_06691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30789_ (.A1(_06301_),
    .A2(_06346_),
    .A3(_06418_),
    .ZN(_06692_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30790_ (.A1(_06691_),
    .A2(_06185_),
    .A3(_06692_),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30791_ (.A1(_06689_),
    .A2(_06693_),
    .A3(_06188_),
    .ZN(_06694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30792_ (.A1(net1195),
    .A2(_06245_),
    .B(_06108_),
    .ZN(_06695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30793_ (.A1(_06514_),
    .A2(_06695_),
    .B(_06341_),
    .ZN(_06696_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30794_ (.A1(_06628_),
    .A2(_06410_),
    .A3(_06227_),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30795_ (.A1(_06696_),
    .A2(_06697_),
    .B(_06243_),
    .ZN(_06698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30796_ (.A1(_06051_),
    .A2(_06218_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30797_ (.A1(_06314_),
    .A2(_06181_),
    .B(_06108_),
    .ZN(_06700_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30798_ (.A1(_06626_),
    .A2(_06699_),
    .A3(_06700_),
    .ZN(_06701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30799_ (.A1(_06290_),
    .A2(net1195),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30800_ (.A1(_06424_),
    .A2(_06702_),
    .A3(_06227_),
    .ZN(_06703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30801_ (.A1(_06701_),
    .A2(_06703_),
    .A3(_06092_),
    .ZN(_06704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30802_ (.A1(_06698_),
    .A2(_06704_),
    .ZN(_06705_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30803_ (.A1(_06694_),
    .A2(_06705_),
    .B(_06414_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30804_ (.A1(_06683_),
    .A2(_06706_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30805_ (.A1(_03769_),
    .A2(_03780_),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30806_ (.A1(_12833_),
    .A2(_03776_),
    .ZN(_06708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30807_ (.A1(_06707_),
    .A2(_06708_),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30808_ (.I(_06709_),
    .ZN(_06710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30809_ (.A1(net914),
    .A2(net530),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30810_ (.A1(_12765_),
    .A2(net778),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30811_ (.A1(_06711_),
    .A2(_06712_),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30812_ (.A1(_06710_),
    .A2(net907),
    .ZN(_06714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30813_ (.I(_06713_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30814_ (.A1(_06715_),
    .A2(_06709_),
    .ZN(_06716_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30815_ (.A1(_06714_),
    .A2(_06716_),
    .A3(_10549_),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30816_ (.I(\u0.tmp_w[1] ),
    .ZN(_06718_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30817_ (.A1(_11989_),
    .A2(\text_in_r[1] ),
    .Z(_06719_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30818_ (.A1(_06717_),
    .A2(_06718_),
    .A3(_06719_),
    .ZN(_06720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30819_ (.A1(_06715_),
    .A2(_06710_),
    .ZN(_06721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30820_ (.A1(_06709_),
    .A2(net907),
    .ZN(_06722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30821_ (.A1(_06722_),
    .A2(_10479_),
    .A3(_06721_),
    .ZN(_06723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30822_ (.A1(_10483_),
    .A2(\text_in_r[1] ),
    .ZN(_06724_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30823_ (.A1(_06724_),
    .A2(\u0.tmp_w[1] ),
    .A3(_06723_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30824_ (.A1(_06720_),
    .A2(_06725_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _30825_ (.I(_06726_),
    .Z(_16175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30826_ (.A1(_12814_),
    .A2(_12816_),
    .A3(_13067_),
    .ZN(_06727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30827_ (.A1(_12780_),
    .A2(_12815_),
    .ZN(_06728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30828_ (.A1(\sa10_sub[0] ),
    .A2(net532),
    .ZN(_06729_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30829_ (.A1(_06728_),
    .A2(_03773_),
    .A3(_06729_),
    .ZN(_06730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30830_ (.A1(_06727_),
    .A2(_06730_),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30831_ (.A1(_06731_),
    .A2(net914),
    .ZN(_06732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30832_ (.A1(_06727_),
    .A2(_06730_),
    .A3(_12765_),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30833_ (.A1(_06732_),
    .A2(_06733_),
    .B(_10525_),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30834_ (.I(\text_in_r[0] ),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30835_ (.A1(_06735_),
    .A2(_10381_),
    .Z(_06736_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30836_ (.A1(_06734_),
    .A2(_06736_),
    .B(\u0.tmp_w[0] ),
    .ZN(_06737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30837_ (.A1(_06732_),
    .A2(_06733_),
    .ZN(_06738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30838_ (.A1(_06738_),
    .A2(_10405_),
    .ZN(_06739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30839_ (.I(\u0.tmp_w[0] ),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30840_ (.I(_06736_),
    .ZN(_06741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30841_ (.A1(_06739_),
    .A2(_06740_),
    .A3(_06741_),
    .ZN(_06742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30842_ (.A1(_06737_),
    .A2(_06742_),
    .ZN(_16178_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30843_ (.A1(net38),
    .A2(_12836_),
    .Z(_06743_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30844_ (.A1(net38),
    .A2(_12836_),
    .ZN(_06744_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30845_ (.A1(_06743_),
    .A2(_06744_),
    .B(\sa03_sr[2] ),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30846_ (.A1(_12766_),
    .A2(_12834_),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30847_ (.A1(net38),
    .A2(_12836_),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30848_ (.A1(_06746_),
    .A2(_12864_),
    .A3(_06747_),
    .ZN(_06748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30849_ (.A1(_06745_),
    .A2(_06748_),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30850_ (.A1(net737),
    .A2(\sa10_sub[2] ),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30851_ (.I(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30852_ (.A1(_06749_),
    .A2(_06751_),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30853_ (.A1(_06750_),
    .A2(_06748_),
    .A3(_06745_),
    .ZN(_06753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30854_ (.A1(_06753_),
    .A2(_06752_),
    .B(net596),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30855_ (.I(\text_in_r[2] ),
    .ZN(_06755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30856_ (.A1(_06755_),
    .A2(net476),
    .Z(_06756_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _30857_ (.A1(_06756_),
    .A2(_06754_),
    .B(\u0.tmp_w[2] ),
    .ZN(_06757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30858_ (.A1(_06752_),
    .A2(_06753_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30859_ (.A1(_06758_),
    .A2(_10378_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30860_ (.I(_06756_),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30861_ (.A1(_06759_),
    .A2(_07556_),
    .A3(_06760_),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30862_ (.A1(_06757_),
    .A2(_06761_),
    .ZN(_06762_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30863_ (.I(_06762_),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30864_ (.I(_06763_),
    .Z(_16194_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30865_ (.A1(_06734_),
    .A2(_06736_),
    .B(_06740_),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30866_ (.A1(_06739_),
    .A2(\u0.tmp_w[0] ),
    .A3(_06741_),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30867_ (.A1(_06764_),
    .A2(_06765_),
    .ZN(_16169_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30868_ (.I(net901),
    .Z(_16187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30869_ (.A1(_06763_),
    .A2(_16169_),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30870_ (.A1(_12867_),
    .A2(\sa21_sub[3] ),
    .ZN(_06767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30871_ (.A1(_12876_),
    .A2(_12870_),
    .ZN(_06768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30872_ (.A1(_06767_),
    .A2(_06768_),
    .ZN(_06769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30873_ (.A1(_03848_),
    .A2(_06769_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30874_ (.A1(_06767_),
    .A2(_06768_),
    .Z(_06771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30875_ (.A1(_03852_),
    .A2(_06771_),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30876_ (.A1(_06770_),
    .A2(_10479_),
    .A3(_06772_),
    .ZN(_06773_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30877_ (.I(\u0.tmp_w[3] ),
    .ZN(_06774_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30878_ (.A1(_10489_),
    .A2(\text_in_r[3] ),
    .Z(_06775_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30879_ (.A1(_06773_),
    .A2(_06774_),
    .A3(_06775_),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30880_ (.A1(_03848_),
    .A2(_06771_),
    .ZN(_06777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30881_ (.A1(_03852_),
    .A2(_06769_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30882_ (.A1(_06777_),
    .A2(_10479_),
    .A3(_06778_),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30883_ (.A1(_10483_),
    .A2(\text_in_r[3] ),
    .ZN(_06780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30884_ (.A1(_06779_),
    .A2(\u0.tmp_w[3] ),
    .A3(_06780_),
    .ZN(_06781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30885_ (.A1(_06776_),
    .A2(_06781_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30886_ (.I(_06782_),
    .Z(_06783_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30887_ (.A1(_06766_),
    .A2(_06783_),
    .Z(_06784_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _30888_ (.I(net903),
    .Z(_06785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30889_ (.A1(net892),
    .A2(_16178_),
    .A3(_06785_),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30890_ (.A1(_06784_),
    .A2(_06786_),
    .ZN(_06787_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _30891_ (.I(net910),
    .Z(_06788_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _30892_ (.I(_06761_),
    .Z(_06789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30893_ (.A1(_06788_),
    .A2(_06789_),
    .A3(_16176_),
    .ZN(_06790_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30894_ (.A1(_06790_),
    .A2(_06782_),
    .Z(_06791_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30895_ (.A1(_12931_),
    .A2(_03869_),
    .B(_10522_),
    .ZN(_06792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30896_ (.A1(_12931_),
    .A2(_03869_),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30897_ (.I(_06793_),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30898_ (.A1(_11203_),
    .A2(\text_in_r[4] ),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30899_ (.A1(_06792_),
    .A2(_06794_),
    .B(_06795_),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30900_ (.A1(_06796_),
    .A2(\u0.tmp_w[4] ),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30901_ (.I(\u0.tmp_w[4] ),
    .ZN(_06798_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _30902_ (.A1(_06792_),
    .A2(_06794_),
    .B(_06798_),
    .C(_06795_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30903_ (.A1(_06799_),
    .A2(_06797_),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30904_ (.A1(_06791_),
    .A2(net85),
    .Z(_06801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30905_ (.A1(_06787_),
    .A2(_06801_),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30906_ (.I(\u0.tmp_w[5] ),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30907_ (.A1(\sa32_sub[4] ),
    .A2(\sa21_sub[5] ),
    .Z(_06804_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30908_ (.A1(_06804_),
    .A2(_00956_),
    .Z(_06805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30909_ (.A1(_06804_),
    .A2(_00956_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30910_ (.A1(_06805_),
    .A2(_06806_),
    .ZN(_06807_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30911_ (.A1(\sa03_sr[4] ),
    .A2(\sa10_sub[5] ),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30912_ (.I(_06808_),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30913_ (.A1(_06807_),
    .A2(_06809_),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30914_ (.A1(_06805_),
    .A2(_06808_),
    .A3(_06806_),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30915_ (.A1(_06810_),
    .A2(_06811_),
    .A3(_10549_),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30916_ (.A1(_10483_),
    .A2(\text_in_r[5] ),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30917_ (.A1(_06812_),
    .A2(_06813_),
    .ZN(_06814_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _30918_ (.A1(_06803_),
    .A2(_06814_),
    .Z(_06815_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30919_ (.I(_06815_),
    .Z(_06816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30920_ (.I(_16172_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30921_ (.A1(_06817_),
    .A2(net904),
    .ZN(_06818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30922_ (.A1(_06782_),
    .A2(_06818_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30923_ (.I(_06800_),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30924_ (.I(_06820_),
    .Z(_06821_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30925_ (.A1(_06819_),
    .A2(_06821_),
    .Z(_06822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30926_ (.A1(_06762_),
    .A2(_16181_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30927_ (.A1(_06823_),
    .A2(_06790_),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30928_ (.A1(_06779_),
    .A2(_06774_),
    .A3(_06780_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30929_ (.A1(_06773_),
    .A2(\u0.tmp_w[3] ),
    .A3(_06775_),
    .ZN(_06826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30930_ (.A1(_06825_),
    .A2(_06826_),
    .ZN(_06827_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30931_ (.I(_06827_),
    .Z(_06828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30932_ (.A1(_06824_),
    .A2(_06828_),
    .ZN(_06829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30933_ (.A1(_06822_),
    .A2(_06829_),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30934_ (.A1(_06802_),
    .A2(_06816_),
    .A3(_06830_),
    .ZN(_06831_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _30935_ (.I(_16176_),
    .ZN(_06832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30936_ (.A1(_06832_),
    .A2(_06785_),
    .ZN(_06833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30937_ (.A1(_06833_),
    .A2(_06783_),
    .ZN(_06834_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30938_ (.A1(_06834_),
    .A2(_06821_),
    .Z(_06835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30939_ (.A1(_06785_),
    .A2(_16173_),
    .ZN(_06836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30940_ (.I(_16171_),
    .ZN(_06837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30941_ (.A1(net1040),
    .A2(_06789_),
    .A3(_06837_),
    .ZN(_06838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30942_ (.A1(_06836_),
    .A2(_06838_),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30943_ (.I(_06827_),
    .Z(_06840_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30944_ (.I(_06840_),
    .Z(_06841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30945_ (.A1(_06839_),
    .A2(_06841_),
    .ZN(_06842_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30946_ (.I(_06815_),
    .Z(_06843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30947_ (.A1(_06835_),
    .A2(_06842_),
    .B(_06843_),
    .ZN(_06844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30948_ (.A1(net892),
    .A2(_06785_),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30949_ (.I(_06827_),
    .Z(_06846_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30950_ (.A1(_06788_),
    .A2(_06789_),
    .A3(_16172_),
    .ZN(_06847_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30951_ (.A1(_06845_),
    .A2(_06846_),
    .A3(_06847_),
    .ZN(_06848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30952_ (.A1(_06763_),
    .A2(_16179_),
    .ZN(_06849_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30953_ (.I(_06783_),
    .Z(_06850_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30954_ (.A1(_06785_),
    .A2(_16169_),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30955_ (.A1(_06849_),
    .A2(_06850_),
    .A3(_06851_),
    .ZN(_06852_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _30956_ (.I(_06800_),
    .Z(_06853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30957_ (.A1(_06848_),
    .A2(_06852_),
    .A3(_06853_),
    .ZN(_06854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30958_ (.A1(_06844_),
    .A2(_06854_),
    .ZN(_06855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30959_ (.A1(_06831_),
    .A2(_06855_),
    .ZN(_06856_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _30960_ (.A1(\sa32_sub[5] ),
    .A2(\sa21_sub[6] ),
    .A3(\sa03_sr[6] ),
    .Z(_06857_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30961_ (.A1(\sa03_sr[5] ),
    .A2(\sa10_sub[6] ),
    .Z(_06858_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30962_ (.A1(_06857_),
    .A2(_06858_),
    .Z(_06859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30963_ (.A1(_06857_),
    .A2(_06858_),
    .ZN(_06860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30964_ (.A1(_06859_),
    .A2(_10523_),
    .A3(_06860_),
    .ZN(_06861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30965_ (.A1(_12115_),
    .A2(\text_in_r[6] ),
    .ZN(_06862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30966_ (.A1(_06861_),
    .A2(_06862_),
    .Z(_06863_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30967_ (.A1(_06863_),
    .A2(\u0.tmp_w[6] ),
    .Z(_06864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30968_ (.A1(_06863_),
    .A2(\u0.tmp_w[6] ),
    .ZN(_06865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30969_ (.A1(_06864_),
    .A2(_06865_),
    .ZN(_06866_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30970_ (.I(_06866_),
    .Z(_06867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30971_ (.A1(_06856_),
    .A2(_06867_),
    .ZN(_06868_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _30972_ (.A1(\sa32_sub[6] ),
    .A2(net976),
    .A3(_13068_),
    .ZN(_06869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30973_ (.A1(_10639_),
    .A2(\text_in_r[7] ),
    .Z(_06870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30974_ (.A1(_06869_),
    .A2(_12965_),
    .B(_06870_),
    .ZN(_06871_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30975_ (.A1(\u0.tmp_w[7] ),
    .A2(_06871_),
    .Z(_06872_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30976_ (.I(_06872_),
    .Z(_06873_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30977_ (.I(_06873_),
    .ZN(_06874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30978_ (.A1(_06868_),
    .A2(_06874_),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30979_ (.A1(_06849_),
    .A2(_06827_),
    .ZN(_06876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30980_ (.I(_06876_),
    .ZN(_06877_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30981_ (.A1(net81),
    .A2(_16169_),
    .A3(_06785_),
    .ZN(_06878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30982_ (.A1(_06877_),
    .A2(_06878_),
    .ZN(_06879_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30983_ (.I(_06821_),
    .Z(_06880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30984_ (.I(_06836_),
    .ZN(_06881_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30985_ (.I(_06782_),
    .Z(_06882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30986_ (.A1(_06881_),
    .A2(_06882_),
    .ZN(_06883_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30987_ (.A1(_06879_),
    .A2(_06880_),
    .A3(_06883_),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30988_ (.A1(_06881_),
    .A2(_06828_),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30989_ (.A1(_06885_),
    .A2(_06853_),
    .Z(_06886_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30990_ (.I(_16181_),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30991_ (.A1(_06887_),
    .A2(_06789_),
    .A3(_06788_),
    .ZN(_06888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30992_ (.A1(_06888_),
    .A2(_06782_),
    .Z(_06889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30993_ (.A1(_06878_),
    .A2(_06889_),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30994_ (.A1(_06886_),
    .A2(_06890_),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _30995_ (.I(_06815_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30996_ (.I(_06892_),
    .Z(_06893_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _30997_ (.I(_06893_),
    .Z(_06894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30998_ (.A1(_06884_),
    .A2(_06891_),
    .A3(_06894_),
    .ZN(_06895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30999_ (.A1(_06837_),
    .A2(net902),
    .ZN(_06896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31000_ (.A1(_06896_),
    .A2(_06840_),
    .B(net85),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31001_ (.A1(_16194_),
    .A2(_16178_),
    .ZN(_06898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31002_ (.A1(_06898_),
    .A2(_06846_),
    .ZN(_06899_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31003_ (.A1(_06897_),
    .A2(_06899_),
    .ZN(_06900_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31004_ (.I(_06840_),
    .Z(_06901_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31005_ (.A1(_06832_),
    .A2(_06789_),
    .A3(net1040),
    .ZN(_06902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31006_ (.A1(_06878_),
    .A2(_06901_),
    .A3(_06902_),
    .ZN(_06903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31007_ (.A1(_16194_),
    .A2(_16173_),
    .Z(_06904_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31008_ (.I(_06846_),
    .Z(_06905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31009_ (.A1(_06904_),
    .A2(_06905_),
    .ZN(_06906_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31010_ (.A1(_06900_),
    .A2(_06903_),
    .A3(_06906_),
    .ZN(_06907_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31011_ (.A1(_06847_),
    .A2(_06840_),
    .Z(_06908_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31012_ (.A1(_06841_),
    .A2(_16192_),
    .ZN(_06909_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31013_ (.A1(_06908_),
    .A2(_06909_),
    .Z(_06910_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31014_ (.I(_06821_),
    .Z(_06911_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31015_ (.I(_06892_),
    .Z(_06912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31016_ (.A1(_06910_),
    .A2(_06911_),
    .B(_06912_),
    .ZN(_06913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31017_ (.A1(_06907_),
    .A2(_06913_),
    .ZN(_06914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31018_ (.A1(_06895_),
    .A2(_06914_),
    .B(_06867_),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31019_ (.A1(_06875_),
    .A2(_06915_),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31020_ (.A1(_06717_),
    .A2(\u0.tmp_w[1] ),
    .A3(_06719_),
    .ZN(_06917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31021_ (.A1(_06723_),
    .A2(_06718_),
    .A3(_06724_),
    .ZN(_06918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31022_ (.A1(_06917_),
    .A2(_06918_),
    .ZN(_16170_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31023_ (.A1(net18),
    .A2(_16194_),
    .Z(_06919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31024_ (.A1(_06919_),
    .A2(_06881_),
    .B(_06828_),
    .ZN(_06920_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31025_ (.I(net85),
    .Z(_06921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31026_ (.A1(_06787_),
    .A2(_06920_),
    .A3(_06921_),
    .ZN(_06922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31027_ (.A1(_16187_),
    .A2(_16185_),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31028_ (.A1(_06898_),
    .A2(_06923_),
    .ZN(_06924_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _31029_ (.I(_06882_),
    .Z(_06925_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _31030_ (.I(_06800_),
    .Z(_06926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31031_ (.A1(_06924_),
    .A2(_06925_),
    .B(_06926_),
    .ZN(_06927_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _31032_ (.A1(net904),
    .A2(_16178_),
    .ZN(_06928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31033_ (.A1(_06928_),
    .A2(net81),
    .ZN(_06929_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31034_ (.I(_06846_),
    .Z(_06930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31035_ (.A1(_16170_),
    .A2(_06785_),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31036_ (.I(_06931_),
    .Z(_06932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31037_ (.A1(_06929_),
    .A2(_06930_),
    .A3(_06932_),
    .ZN(_06933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31038_ (.A1(_06927_),
    .A2(_06933_),
    .ZN(_06934_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31039_ (.I(_06843_),
    .Z(_06935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31040_ (.A1(_06922_),
    .A2(_06934_),
    .A3(_06935_),
    .ZN(_06936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _31041_ (.I(_06834_),
    .ZN(_06937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31042_ (.A1(_06937_),
    .A2(_06929_),
    .ZN(_06938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31043_ (.A1(_06766_),
    .A2(_06840_),
    .Z(_06939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31044_ (.I(_06939_),
    .ZN(_06940_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31045_ (.I(_06800_),
    .Z(_06941_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31046_ (.A1(_06938_),
    .A2(_06940_),
    .A3(_06941_),
    .ZN(_06942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31047_ (.A1(_06785_),
    .A2(net906),
    .ZN(_06943_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31048_ (.A1(net1040),
    .A2(_06789_),
    .A3(_16185_),
    .ZN(_06944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31049_ (.A1(_06943_),
    .A2(_06944_),
    .ZN(_06945_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31050_ (.I(_06882_),
    .Z(_06946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31051_ (.A1(_06945_),
    .A2(_06946_),
    .B(_06926_),
    .ZN(_06947_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31052_ (.A1(_06929_),
    .A2(_06828_),
    .A3(_06851_),
    .ZN(_06948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31053_ (.A1(_06947_),
    .A2(_06948_),
    .ZN(_06949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31054_ (.A1(_06942_),
    .A2(_06949_),
    .A3(_06912_),
    .ZN(_06950_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _31055_ (.I(_06866_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31056_ (.I(_06951_),
    .Z(_06952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31057_ (.A1(_06936_),
    .A2(_06950_),
    .B(_06952_),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _31058_ (.I(_06819_),
    .ZN(_06954_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31059_ (.A1(net1040),
    .A2(_06789_),
    .A3(_16171_),
    .ZN(_06955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31060_ (.A1(_06954_),
    .A2(_06955_),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _31061_ (.I(_06896_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _31062_ (.A1(_06785_),
    .A2(_16179_),
    .ZN(_06958_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31063_ (.A1(_06957_),
    .A2(_06958_),
    .B(_06905_),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31064_ (.I(_06821_),
    .Z(_06960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31065_ (.A1(_06956_),
    .A2(_06959_),
    .B(_06960_),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31066_ (.A1(_06788_),
    .A2(_06817_),
    .A3(_06789_),
    .ZN(_06962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31067_ (.A1(_06783_),
    .A2(_06962_),
    .Z(_06963_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31068_ (.A1(_06963_),
    .A2(_06853_),
    .ZN(_06964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31069_ (.A1(net81),
    .A2(_16194_),
    .ZN(_06965_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31070_ (.A1(_06965_),
    .A2(_06901_),
    .A3(_06943_),
    .ZN(_06966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31071_ (.A1(_06964_),
    .A2(_06966_),
    .ZN(_06967_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31072_ (.I(_06815_),
    .Z(_06968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31073_ (.A1(_06967_),
    .A2(_06968_),
    .ZN(_06969_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31074_ (.A1(_06961_),
    .A2(_06969_),
    .B(_06951_),
    .ZN(_06970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31075_ (.A1(_06785_),
    .A2(_16178_),
    .ZN(_06971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31076_ (.A1(_06971_),
    .A2(_06840_),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31077_ (.A1(net18),
    .A2(_16169_),
    .ZN(_06973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31078_ (.A1(_06972_),
    .A2(_06973_),
    .ZN(_06974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31079_ (.A1(net912),
    .A2(_16169_),
    .ZN(_06975_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31080_ (.A1(_06975_),
    .A2(_06898_),
    .A3(_06850_),
    .ZN(_06976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31081_ (.A1(_06974_),
    .A2(_06976_),
    .A3(_06960_),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31082_ (.A1(_06818_),
    .A2(_06840_),
    .ZN(_06978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31083_ (.I(_06978_),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31084_ (.A1(net81),
    .A2(_16194_),
    .A3(_16178_),
    .ZN(_06980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31085_ (.A1(_06979_),
    .A2(_06980_),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31086_ (.I(_06800_),
    .Z(_06982_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31087_ (.I(_16179_),
    .ZN(_06983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31088_ (.A1(_16187_),
    .A2(_06983_),
    .ZN(_06984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31089_ (.A1(_06984_),
    .A2(_06838_),
    .ZN(_06985_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _31090_ (.I(_06783_),
    .Z(_06986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31091_ (.A1(_06985_),
    .A2(_06986_),
    .ZN(_06987_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31092_ (.A1(_06981_),
    .A2(_06982_),
    .A3(_06987_),
    .ZN(_06988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31093_ (.A1(_06977_),
    .A2(_06988_),
    .B(_06968_),
    .ZN(_06989_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31094_ (.A1(_06970_),
    .A2(_06989_),
    .B(_06873_),
    .ZN(_06990_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31095_ (.A1(_06953_),
    .A2(_06990_),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31096_ (.A1(_06916_),
    .A2(_06991_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31097_ (.A1(_06975_),
    .A2(_16194_),
    .ZN(_06992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31098_ (.A1(net892),
    .A2(_16178_),
    .ZN(_06993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31099_ (.A1(_06993_),
    .A2(_16187_),
    .ZN(_06994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31100_ (.A1(_06992_),
    .A2(_06994_),
    .Z(_06995_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31101_ (.A1(_06851_),
    .A2(_06828_),
    .A3(_06955_),
    .ZN(_06996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31102_ (.A1(_06996_),
    .A2(_06892_),
    .Z(_06997_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31103_ (.A1(_06930_),
    .A2(_06995_),
    .B(_06997_),
    .ZN(_06998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31104_ (.A1(_06972_),
    .A2(_06965_),
    .ZN(_06999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31105_ (.A1(net900),
    .A2(_06763_),
    .ZN(_07000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31106_ (.A1(_06937_),
    .A2(_07000_),
    .ZN(_07001_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31107_ (.A1(_06999_),
    .A2(_07001_),
    .A3(_06968_),
    .ZN(_07002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31108_ (.A1(_06998_),
    .A2(_06880_),
    .A3(_07002_),
    .ZN(_07003_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31109_ (.A1(_06892_),
    .A2(_16195_),
    .A3(_06901_),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31110_ (.A1(_06877_),
    .A2(_06786_),
    .ZN(_07005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31111_ (.A1(_07004_),
    .A2(_07005_),
    .ZN(_07006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31112_ (.A1(_07006_),
    .A2(_06921_),
    .B(_06866_),
    .ZN(_07007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31113_ (.A1(_07003_),
    .A2(_07007_),
    .B(_06874_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31114_ (.A1(_06786_),
    .A2(_06846_),
    .ZN(_07009_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31115_ (.A1(_07009_),
    .A2(_06928_),
    .B(_06941_),
    .C(_06819_),
    .ZN(_07010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31116_ (.A1(_06980_),
    .A2(_06882_),
    .ZN(_07011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _31117_ (.I(_06943_),
    .ZN(_07012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31118_ (.A1(_07011_),
    .A2(_07012_),
    .Z(_07013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _31119_ (.I(_16185_),
    .ZN(_07014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31120_ (.A1(net904),
    .A2(_07014_),
    .ZN(_07015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31121_ (.A1(_07015_),
    .A2(_06840_),
    .Z(_07016_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31122_ (.I(_16173_),
    .ZN(_07017_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31123_ (.A1(net1040),
    .A2(_06789_),
    .A3(_07017_),
    .ZN(_07018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31124_ (.A1(_07016_),
    .A2(_07018_),
    .B(_06926_),
    .ZN(_07019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31125_ (.A1(_07013_),
    .A2(_07019_),
    .ZN(_07020_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31126_ (.A1(_07010_),
    .A2(_07020_),
    .A3(_06935_),
    .ZN(_07021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31127_ (.A1(_06957_),
    .A2(_06850_),
    .ZN(_07022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31128_ (.A1(_06885_),
    .A2(_07022_),
    .Z(_07023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31129_ (.I(_06898_),
    .ZN(_07024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31130_ (.A1(_07024_),
    .A2(_06841_),
    .B(net85),
    .ZN(_07025_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31131_ (.I(_06847_),
    .ZN(_07026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31132_ (.A1(_07026_),
    .A2(_06882_),
    .ZN(_07027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31133_ (.A1(_07023_),
    .A2(_07025_),
    .A3(_07027_),
    .ZN(_07028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31134_ (.A1(_06972_),
    .A2(_06955_),
    .ZN(_07029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31135_ (.A1(_07029_),
    .A2(_07001_),
    .A3(_06941_),
    .ZN(_07030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31136_ (.A1(_07028_),
    .A2(_06894_),
    .A3(_07030_),
    .ZN(_07031_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31137_ (.A1(_07021_),
    .A2(_07031_),
    .A3(_06867_),
    .ZN(_07032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31138_ (.A1(_07008_),
    .A2(_07032_),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31139_ (.A1(_06783_),
    .A2(_16187_),
    .ZN(_07034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31140_ (.A1(_06782_),
    .A2(net18),
    .ZN(_07035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31141_ (.A1(_07034_),
    .A2(_07035_),
    .ZN(_07036_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31142_ (.A1(_07036_),
    .A2(net85),
    .ZN(_07037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31143_ (.A1(_06791_),
    .A2(_06932_),
    .Z(_07038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31144_ (.A1(_07037_),
    .A2(_07038_),
    .B(_06893_),
    .ZN(_07039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31145_ (.A1(_06963_),
    .A2(_07015_),
    .ZN(_07040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31146_ (.A1(_06903_),
    .A2(_06941_),
    .A3(_07040_),
    .ZN(_07041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31147_ (.A1(_07039_),
    .A2(_07041_),
    .B(_06866_),
    .ZN(_07042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31148_ (.A1(_06898_),
    .A2(_06846_),
    .Z(_07043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31149_ (.A1(_07043_),
    .A2(_06833_),
    .ZN(_07044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31150_ (.A1(_06784_),
    .A2(_06818_),
    .ZN(_07045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31151_ (.A1(_07044_),
    .A2(_07045_),
    .A3(_06911_),
    .ZN(_07046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31152_ (.A1(_06845_),
    .A2(_06973_),
    .A3(_06841_),
    .ZN(_07047_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31153_ (.A1(_06783_),
    .A2(_16194_),
    .Z(_07048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31154_ (.A1(_07048_),
    .A2(_06975_),
    .ZN(_07049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31155_ (.A1(_07047_),
    .A2(_06941_),
    .A3(_07049_),
    .ZN(_07050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31156_ (.A1(_07046_),
    .A2(_07050_),
    .A3(_06894_),
    .ZN(_07051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31157_ (.A1(_07042_),
    .A2(_07051_),
    .B(_06873_),
    .ZN(_07052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31158_ (.A1(_06788_),
    .A2(_06789_),
    .A3(_07014_),
    .ZN(_07053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31159_ (.A1(_06783_),
    .A2(_07053_),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31160_ (.A1(_07054_),
    .A2(_06932_),
    .ZN(_07055_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31161_ (.A1(_06925_),
    .A2(_06994_),
    .B(_07055_),
    .C(_06960_),
    .ZN(_07056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31162_ (.A1(_06828_),
    .A2(_16176_),
    .Z(_07057_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _31163_ (.I(_06820_),
    .Z(_07058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31164_ (.A1(_07057_),
    .A2(_16187_),
    .B(_07058_),
    .ZN(_07059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31165_ (.A1(_07013_),
    .A2(_07059_),
    .ZN(_07060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31166_ (.A1(_07056_),
    .A2(_07060_),
    .A3(_06894_),
    .ZN(_07061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31167_ (.A1(_07043_),
    .A2(_06896_),
    .ZN(_07062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31168_ (.A1(_06954_),
    .A2(_06790_),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31169_ (.A1(_07062_),
    .A2(_07063_),
    .ZN(_07064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31170_ (.A1(_07064_),
    .A2(_06880_),
    .ZN(_07065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31171_ (.I(_06993_),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31172_ (.I(_06851_),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31173_ (.A1(_07066_),
    .A2(_07067_),
    .B(_06986_),
    .ZN(_07068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31174_ (.A1(_06908_),
    .A2(_06851_),
    .ZN(_07069_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31175_ (.A1(_07068_),
    .A2(_06941_),
    .A3(_07069_),
    .ZN(_07070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31176_ (.A1(_07065_),
    .A2(_07070_),
    .A3(_06935_),
    .ZN(_07071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31177_ (.A1(_07061_),
    .A2(_07071_),
    .A3(_06867_),
    .ZN(_07072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31178_ (.A1(_07072_),
    .A2(_07052_),
    .ZN(_07073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31179_ (.A1(_07033_),
    .A2(_07073_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31180_ (.A1(_06929_),
    .A2(_06930_),
    .B(_07058_),
    .ZN(_07074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31181_ (.A1(_06980_),
    .A2(_06925_),
    .A3(_07015_),
    .ZN(_07075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31182_ (.A1(_07074_),
    .A2(_07075_),
    .B(_06968_),
    .ZN(_07076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31183_ (.A1(_16187_),
    .A2(_16178_),
    .Z(_07077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31184_ (.A1(_06904_),
    .A2(_07077_),
    .B(_06925_),
    .ZN(_07078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31185_ (.A1(_06965_),
    .A2(_06930_),
    .A3(_06818_),
    .ZN(_07079_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31186_ (.A1(_07078_),
    .A2(_07079_),
    .A3(_06880_),
    .ZN(_07080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31187_ (.A1(_07076_),
    .A2(_07080_),
    .B(_06866_),
    .ZN(_07081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31188_ (.A1(_06845_),
    .A2(net913),
    .A3(_06850_),
    .ZN(_07082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31189_ (.I(_07082_),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31190_ (.A1(_06833_),
    .A2(_06840_),
    .ZN(_07084_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31191_ (.I(_07053_),
    .ZN(_07085_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31192_ (.A1(_07084_),
    .A2(_07085_),
    .ZN(_07086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31193_ (.A1(_07083_),
    .A2(_07086_),
    .B(_07058_),
    .ZN(_07087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31194_ (.A1(_06851_),
    .A2(_06902_),
    .ZN(_07088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31195_ (.A1(_07088_),
    .A2(_06986_),
    .A3(_06932_),
    .ZN(_07089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31196_ (.A1(_07089_),
    .A2(_06982_),
    .A3(_06848_),
    .ZN(_07090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31197_ (.A1(_07087_),
    .A2(_07090_),
    .ZN(_07091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31198_ (.A1(_07091_),
    .A2(_06935_),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31199_ (.A1(_07081_),
    .A2(_07092_),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31200_ (.A1(_07000_),
    .A2(_06986_),
    .A3(_06823_),
    .ZN(_07094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31201_ (.A1(_06971_),
    .A2(_06841_),
    .A3(_06944_),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31202_ (.A1(_07094_),
    .A2(_07058_),
    .A3(_07095_),
    .ZN(_07096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31203_ (.A1(_06851_),
    .A2(_06828_),
    .A3(_06888_),
    .ZN(_07097_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31204_ (.A1(_06818_),
    .A2(_06847_),
    .A3(_06850_),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31205_ (.A1(_07097_),
    .A2(_07098_),
    .ZN(_07099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31206_ (.A1(_07099_),
    .A2(_06982_),
    .ZN(_07100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31207_ (.A1(_07096_),
    .A2(_07100_),
    .ZN(_07101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31208_ (.A1(_07101_),
    .A2(_06894_),
    .ZN(_07102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31209_ (.A1(_06932_),
    .A2(_06946_),
    .A3(net1041),
    .ZN(_07103_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31210_ (.A1(_07103_),
    .A2(_06829_),
    .A3(_06941_),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31211_ (.A1(_06823_),
    .A2(_06944_),
    .ZN(_07105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31212_ (.A1(_07105_),
    .A2(_06930_),
    .ZN(_07106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31213_ (.A1(_06851_),
    .A2(_06986_),
    .A3(net1041),
    .ZN(_07107_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31214_ (.A1(_07106_),
    .A2(_07107_),
    .A3(_06960_),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31215_ (.A1(_07104_),
    .A2(_07108_),
    .A3(_06968_),
    .ZN(_07109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31216_ (.A1(_07102_),
    .A2(_07109_),
    .A3(_06867_),
    .ZN(_07110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31217_ (.A1(_07093_),
    .A2(_06873_),
    .A3(_07110_),
    .ZN(_07111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31218_ (.A1(_06984_),
    .A2(_06882_),
    .Z(_07112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31219_ (.A1(_07112_),
    .A2(_06847_),
    .Z(_07113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31220_ (.A1(_06845_),
    .A2(_06841_),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31221_ (.I(_06838_),
    .ZN(_07115_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31222_ (.A1(_07114_),
    .A2(_07115_),
    .ZN(_07116_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31223_ (.A1(_07113_),
    .A2(_07116_),
    .B(_06880_),
    .ZN(_07117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31224_ (.A1(_06845_),
    .A2(_06973_),
    .A3(_06882_),
    .ZN(_07118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31225_ (.A1(_07118_),
    .A2(_06853_),
    .Z(_07119_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31226_ (.A1(_06986_),
    .A2(_16195_),
    .Z(_07120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31227_ (.A1(_07119_),
    .A2(_07120_),
    .ZN(_07121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31228_ (.A1(_07117_),
    .A2(_07121_),
    .A3(_06935_),
    .ZN(_07122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31229_ (.A1(_07000_),
    .A2(_06882_),
    .Z(_07123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31230_ (.A1(_07123_),
    .A2(_06851_),
    .ZN(_07124_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31231_ (.A1(_07124_),
    .A2(_06911_),
    .A3(_06848_),
    .ZN(_07125_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _31232_ (.I(_06820_),
    .Z(_07126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31233_ (.A1(_16192_),
    .A2(_06905_),
    .B(_07126_),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31234_ (.A1(_06878_),
    .A2(_06963_),
    .ZN(_07128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31235_ (.A1(_07127_),
    .A2(_07128_),
    .B(_06816_),
    .ZN(_07129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31236_ (.A1(_07125_),
    .A2(_07129_),
    .B(_06952_),
    .ZN(_07130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31237_ (.A1(_07122_),
    .A2(_07130_),
    .ZN(_07131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31238_ (.A1(_07000_),
    .A2(_06766_),
    .ZN(_07132_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31239_ (.I(_07132_),
    .ZN(_07133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31240_ (.A1(_07017_),
    .A2(_06832_),
    .ZN(_07134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31241_ (.A1(_16187_),
    .A2(_07134_),
    .ZN(_07135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31242_ (.A1(_07133_),
    .A2(_07135_),
    .ZN(_07136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31243_ (.A1(_07136_),
    .A2(_06925_),
    .ZN(_07137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31244_ (.A1(_06877_),
    .A2(_06786_),
    .B(_06926_),
    .ZN(_07138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31245_ (.A1(_07137_),
    .A2(_07138_),
    .ZN(_07139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31246_ (.A1(_06957_),
    .A2(_06828_),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31247_ (.A1(_07140_),
    .A2(_06853_),
    .Z(_07141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31248_ (.A1(_06954_),
    .A2(net1042),
    .ZN(_07142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31249_ (.A1(_07141_),
    .A2(_07142_),
    .B(_06816_),
    .ZN(_07143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31250_ (.A1(_07139_),
    .A2(_07143_),
    .ZN(_07144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31251_ (.A1(_06929_),
    .A2(_06841_),
    .ZN(_07145_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31252_ (.A1(_06846_),
    .A2(_16190_),
    .Z(_07146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31253_ (.A1(_07145_),
    .A2(_07146_),
    .ZN(_07147_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31254_ (.A1(_07147_),
    .A2(_07058_),
    .Z(_07148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31255_ (.A1(_16199_),
    .A2(_06905_),
    .B(_06853_),
    .ZN(_07149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31256_ (.A1(_07082_),
    .A2(_07149_),
    .B(_06893_),
    .ZN(_07150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31257_ (.A1(_07148_),
    .A2(_07150_),
    .ZN(_07151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31258_ (.A1(_07144_),
    .A2(_07151_),
    .A3(_06952_),
    .ZN(_07152_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31259_ (.A1(_07131_),
    .A2(_07152_),
    .A3(_06874_),
    .ZN(_07153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31260_ (.A1(_07111_),
    .A2(_07153_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31261_ (.A1(_06900_),
    .A2(_07047_),
    .ZN(_07154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31262_ (.I(_06823_),
    .ZN(_07155_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31263_ (.A1(_07155_),
    .A2(_06928_),
    .B(_06882_),
    .ZN(_07156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31264_ (.A1(_06945_),
    .A2(_06841_),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31265_ (.A1(_07156_),
    .A2(_07126_),
    .A3(_07157_),
    .ZN(_07158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31266_ (.A1(_07154_),
    .A2(_07158_),
    .ZN(_07159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31267_ (.A1(_07159_),
    .A2(_06912_),
    .ZN(_07160_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31268_ (.A1(_16194_),
    .A2(_07134_),
    .B(_06888_),
    .C(_06882_),
    .ZN(_07161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31269_ (.A1(_07005_),
    .A2(_07161_),
    .ZN(_07162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31270_ (.A1(_07162_),
    .A2(_06982_),
    .ZN(_07163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31271_ (.A1(_07095_),
    .A2(_07058_),
    .B(_06893_),
    .ZN(_07164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31272_ (.A1(_07163_),
    .A2(_07164_),
    .ZN(_07165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31273_ (.A1(_07160_),
    .A2(_07165_),
    .A3(_06867_),
    .ZN(_07166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31274_ (.A1(_06939_),
    .A2(_06818_),
    .ZN(_07167_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31275_ (.A1(_16194_),
    .A2(_07134_),
    .B(_07053_),
    .C(_06850_),
    .ZN(_07168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31276_ (.A1(_07167_),
    .A2(_07168_),
    .A3(_06843_),
    .ZN(_07169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31277_ (.A1(_07155_),
    .A2(_06850_),
    .ZN(_07170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31278_ (.A1(_07097_),
    .A2(_07170_),
    .A3(_06893_),
    .ZN(_07171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31279_ (.A1(_07169_),
    .A2(_07171_),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31280_ (.A1(_07172_),
    .A2(_06921_),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31281_ (.I(_06818_),
    .ZN(_07174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31282_ (.A1(_07174_),
    .A2(_06828_),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31283_ (.I(_07175_),
    .ZN(_07176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31284_ (.A1(_06883_),
    .A2(_07126_),
    .ZN(_07177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31285_ (.A1(_06893_),
    .A2(_07176_),
    .B(_07177_),
    .ZN(_07178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31286_ (.I(_06845_),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31287_ (.A1(_06876_),
    .A2(_07179_),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _31288_ (.I(_06962_),
    .ZN(_07181_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31289_ (.A1(_07181_),
    .A2(_06783_),
    .Z(_07182_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31290_ (.A1(_07180_),
    .A2(_07182_),
    .B(_06843_),
    .ZN(_07183_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31291_ (.A1(_07178_),
    .A2(_07183_),
    .B(_06866_),
    .ZN(_07184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31292_ (.A1(_07173_),
    .A2(_07184_),
    .ZN(_07185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31293_ (.A1(_07166_),
    .A2(_07185_),
    .ZN(_07186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31294_ (.A1(_07186_),
    .A2(_06873_),
    .ZN(_07187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31295_ (.I(_07182_),
    .ZN(_07188_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31296_ (.A1(_06999_),
    .A2(_06816_),
    .A3(_07188_),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31297_ (.A1(_06963_),
    .A2(_06896_),
    .ZN(_07190_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31298_ (.A1(_06898_),
    .A2(_06901_),
    .A3(_06984_),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31299_ (.A1(_07190_),
    .A2(_07191_),
    .A3(_06893_),
    .ZN(_07192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31300_ (.A1(_07192_),
    .A2(_07189_),
    .ZN(_07193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31301_ (.A1(_07193_),
    .A2(_06880_),
    .ZN(_07194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31302_ (.A1(_06972_),
    .A2(net913),
    .ZN(_07195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31303_ (.A1(_06954_),
    .A2(_07000_),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31304_ (.A1(_07195_),
    .A2(_07196_),
    .A3(_06968_),
    .ZN(_07197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31305_ (.A1(_06943_),
    .A2(_06846_),
    .Z(_07198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31306_ (.A1(_07198_),
    .A2(_07000_),
    .ZN(_07199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31307_ (.A1(_07015_),
    .A2(net1042),
    .A3(_06986_),
    .ZN(_07200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31308_ (.A1(_07199_),
    .A2(_06912_),
    .A3(_07200_),
    .ZN(_07201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31309_ (.A1(_07197_),
    .A2(_07201_),
    .A3(_06921_),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31310_ (.A1(_07194_),
    .A2(_07202_),
    .A3(_06952_),
    .ZN(_07203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31311_ (.A1(_07198_),
    .A2(_06888_),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31312_ (.A1(_07204_),
    .A2(_07055_),
    .A3(_06911_),
    .ZN(_07205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31313_ (.A1(_07034_),
    .A2(_06853_),
    .Z(_07206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31314_ (.A1(_06975_),
    .A2(_06971_),
    .ZN(_07207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31315_ (.A1(_07206_),
    .A2(_07207_),
    .B(_06893_),
    .ZN(_07208_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31316_ (.A1(_07205_),
    .A2(_07208_),
    .B(_06951_),
    .ZN(_07209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31317_ (.A1(_06992_),
    .A2(_07112_),
    .ZN(_07210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31318_ (.A1(_06994_),
    .A2(_06908_),
    .ZN(_07211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31319_ (.A1(_07210_),
    .A2(_07211_),
    .A3(_06982_),
    .ZN(_07212_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31320_ (.A1(_06978_),
    .A2(_06958_),
    .Z(_07213_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31321_ (.A1(_07213_),
    .A2(_06976_),
    .A3(_07058_),
    .ZN(_07214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31322_ (.A1(_07212_),
    .A2(_07214_),
    .ZN(_07215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31323_ (.A1(_07215_),
    .A2(_06894_),
    .ZN(_07216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31324_ (.A1(_07209_),
    .A2(_07216_),
    .ZN(_07217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31325_ (.A1(_07203_),
    .A2(_07217_),
    .A3(_06874_),
    .ZN(_07218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31326_ (.A1(_07187_),
    .A2(_07218_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31327_ (.A1(_07048_),
    .A2(net81),
    .Z(_07219_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31328_ (.A1(_07219_),
    .A2(_06897_),
    .ZN(_07220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31329_ (.A1(_07220_),
    .A2(_06903_),
    .ZN(_07221_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31330_ (.A1(_07086_),
    .A2(_06926_),
    .ZN(_07222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31331_ (.A1(_07123_),
    .A2(_06878_),
    .ZN(_07223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31332_ (.A1(_07222_),
    .A2(_07223_),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31333_ (.A1(_07221_),
    .A2(_06935_),
    .A3(_07224_),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31334_ (.A1(_07027_),
    .A2(_07126_),
    .Z(_07226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31335_ (.A1(_07226_),
    .A2(_06829_),
    .A3(_07170_),
    .ZN(_07227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31336_ (.A1(_07016_),
    .A2(_06962_),
    .ZN(_07228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31337_ (.A1(_07228_),
    .A2(_06890_),
    .A3(_06921_),
    .ZN(_07229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31338_ (.A1(_07227_),
    .A2(_07229_),
    .A3(_06894_),
    .ZN(_07230_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31339_ (.A1(_07225_),
    .A2(_07230_),
    .A3(_06952_),
    .ZN(_07231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31340_ (.A1(_06999_),
    .A2(_07118_),
    .A3(_06921_),
    .ZN(_07233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31341_ (.A1(_06932_),
    .A2(_06993_),
    .A3(_06905_),
    .ZN(_07234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31342_ (.A1(_06932_),
    .A2(_06946_),
    .A3(_06955_),
    .ZN(_07235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31343_ (.A1(_07234_),
    .A2(_07235_),
    .A3(_06911_),
    .ZN(_07236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31344_ (.A1(_07233_),
    .A2(_07236_),
    .A3(_06935_),
    .ZN(_07237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31345_ (.A1(_07036_),
    .A2(_06851_),
    .ZN(_07238_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31346_ (.A1(_07238_),
    .A2(_06921_),
    .A3(_06996_),
    .ZN(_07239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31347_ (.A1(_07126_),
    .A2(_06836_),
    .Z(_07240_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31348_ (.I(_06889_),
    .ZN(_07241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31349_ (.A1(_07240_),
    .A2(_07241_),
    .B(_06816_),
    .ZN(_07242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31350_ (.A1(_07239_),
    .A2(_07242_),
    .ZN(_07244_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31351_ (.A1(_07237_),
    .A2(_06867_),
    .A3(_07244_),
    .ZN(_07245_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31352_ (.A1(_07231_),
    .A2(_07245_),
    .A3(_06874_),
    .ZN(_07246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31353_ (.A1(net913),
    .A2(_16187_),
    .A3(_06905_),
    .ZN(_07247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31354_ (.A1(_06889_),
    .A2(_06931_),
    .ZN(_07248_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31355_ (.A1(_07247_),
    .A2(_07248_),
    .B(_06982_),
    .ZN(_07249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31356_ (.A1(_06901_),
    .A2(_16183_),
    .ZN(_07250_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31357_ (.A1(_07027_),
    .A2(_06926_),
    .A3(_07250_),
    .Z(_07251_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31358_ (.A1(_07249_),
    .A2(_07251_),
    .B(_06912_),
    .ZN(_07252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31359_ (.A1(_07000_),
    .A2(net913),
    .A3(_06901_),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31360_ (.A1(_06889_),
    .A2(_06971_),
    .ZN(_07255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31361_ (.A1(_07253_),
    .A2(_07255_),
    .A3(_06911_),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31362_ (.A1(_06976_),
    .A2(_06941_),
    .A3(_06842_),
    .ZN(_07257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31363_ (.A1(_07256_),
    .A2(_07257_),
    .A3(_06935_),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31364_ (.A1(_07252_),
    .A2(_07258_),
    .A3(_06952_),
    .ZN(_07259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31365_ (.A1(_07000_),
    .A2(net905),
    .ZN(_07260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31366_ (.A1(_07260_),
    .A2(_06930_),
    .ZN(_07261_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31367_ (.A1(_07261_),
    .A2(_07001_),
    .A3(_06911_),
    .ZN(_07262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31368_ (.A1(_06972_),
    .A2(_07053_),
    .ZN(_07263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31369_ (.I(_07048_),
    .ZN(_07264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31370_ (.A1(_07263_),
    .A2(_06941_),
    .A3(_07264_),
    .ZN(_07266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31371_ (.A1(_07262_),
    .A2(_07266_),
    .A3(_06935_),
    .ZN(_07267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31372_ (.A1(_06908_),
    .A2(_06833_),
    .ZN(_07268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31373_ (.A1(_06787_),
    .A2(_06941_),
    .A3(_07268_),
    .ZN(_07269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31374_ (.A1(_07018_),
    .A2(_06846_),
    .ZN(_07270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31375_ (.A1(_07270_),
    .A2(_06821_),
    .Z(_07271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31376_ (.A1(_07011_),
    .A2(_07271_),
    .B(_06816_),
    .ZN(_07272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31377_ (.A1(_07269_),
    .A2(_07272_),
    .ZN(_07273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31378_ (.A1(_07267_),
    .A2(_06867_),
    .A3(_07273_),
    .ZN(_07274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31379_ (.A1(_07259_),
    .A2(_07274_),
    .A3(_06873_),
    .ZN(_07275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31380_ (.A1(_07246_),
    .A2(_07275_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31381_ (.A1(net1039),
    .A2(_16187_),
    .B(_06828_),
    .ZN(_07277_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31382_ (.A1(_07067_),
    .A2(_06958_),
    .ZN(_07278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31383_ (.A1(_07277_),
    .A2(_07278_),
    .ZN(_07279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31384_ (.A1(_06993_),
    .A2(_06766_),
    .A3(_06901_),
    .ZN(_07280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31385_ (.A1(_07279_),
    .A2(_06960_),
    .A3(_07280_),
    .ZN(_07281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31386_ (.A1(_07253_),
    .A2(_06982_),
    .A3(_07035_),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31387_ (.A1(_07281_),
    .A2(_07282_),
    .A3(_06912_),
    .ZN(_07283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31388_ (.A1(_07179_),
    .A2(_07270_),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31389_ (.I(_07027_),
    .ZN(_07285_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31390_ (.A1(_07284_),
    .A2(_07285_),
    .B(_07058_),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31391_ (.A1(_06944_),
    .A2(_06901_),
    .ZN(_07288_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31392_ (.A1(_06819_),
    .A2(_07115_),
    .B(_06926_),
    .C(_07288_),
    .ZN(_07289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31393_ (.A1(_07287_),
    .A2(_07289_),
    .A3(_06968_),
    .ZN(_07290_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31394_ (.A1(_07283_),
    .A2(_06952_),
    .A3(_07290_),
    .ZN(_07291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31395_ (.A1(_06783_),
    .A2(_16176_),
    .ZN(_07292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31396_ (.A1(_07292_),
    .A2(_06820_),
    .ZN(_07293_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31397_ (.A1(_06836_),
    .A2(_06846_),
    .ZN(_07294_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31398_ (.A1(_07293_),
    .A2(_07294_),
    .ZN(_07295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31399_ (.A1(_06888_),
    .A2(_06840_),
    .Z(_07296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31400_ (.A1(_06878_),
    .A2(_07296_),
    .ZN(_07298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31401_ (.A1(_07295_),
    .A2(_07298_),
    .B(_06843_),
    .ZN(_07299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31402_ (.A1(_07054_),
    .A2(_06833_),
    .ZN(_07300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31403_ (.A1(_06920_),
    .A2(_07300_),
    .A3(_06926_),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31404_ (.A1(_07299_),
    .A2(_07301_),
    .ZN(_07302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31405_ (.A1(_07084_),
    .A2(_06821_),
    .Z(_07303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31406_ (.A1(_07303_),
    .A2(_07049_),
    .B(_06892_),
    .ZN(_07304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31407_ (.A1(_07156_),
    .A2(_06853_),
    .A3(_06978_),
    .ZN(_07305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31408_ (.A1(_07304_),
    .A2(_07305_),
    .ZN(_07306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31409_ (.A1(_07302_),
    .A2(_07306_),
    .ZN(_07307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31410_ (.A1(_07307_),
    .A2(_06867_),
    .ZN(_07309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31411_ (.A1(_07309_),
    .A2(_07291_),
    .ZN(_07310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31412_ (.A1(_07310_),
    .A2(_06874_),
    .ZN(_07311_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31413_ (.A1(_06925_),
    .A2(_07088_),
    .B(_06787_),
    .C(_06921_),
    .ZN(_07312_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31414_ (.A1(_07009_),
    .A2(_07085_),
    .Z(_07313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31415_ (.A1(_06958_),
    .A2(_06925_),
    .B(_06926_),
    .ZN(_07314_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31416_ (.A1(_07313_),
    .A2(_07314_),
    .B(_06912_),
    .ZN(_07315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31417_ (.A1(_07312_),
    .A2(_07315_),
    .ZN(_07316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31418_ (.A1(_16178_),
    .A2(_06946_),
    .B(_07126_),
    .ZN(_07317_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31419_ (.A1(_07317_),
    .A2(_06974_),
    .B(_06816_),
    .ZN(_07318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31420_ (.A1(_06954_),
    .A2(_06929_),
    .ZN(_07320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31421_ (.A1(_07296_),
    .A2(_06931_),
    .ZN(_07321_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31422_ (.A1(_07320_),
    .A2(_07321_),
    .A3(_06911_),
    .ZN(_07322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31423_ (.A1(_07318_),
    .A2(_07322_),
    .B(_06951_),
    .ZN(_07323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31424_ (.A1(_07323_),
    .A2(_07316_),
    .ZN(_07324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31425_ (.A1(_06791_),
    .A2(_07126_),
    .Z(_07325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31426_ (.I(_07054_),
    .ZN(_07326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31427_ (.A1(_07325_),
    .A2(_07326_),
    .B(_06968_),
    .ZN(_07327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31428_ (.A1(_06850_),
    .A2(_16173_),
    .ZN(_07328_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31429_ (.A1(_06834_),
    .A2(_06853_),
    .A3(_07328_),
    .Z(_07329_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31430_ (.A1(_06929_),
    .A2(_06786_),
    .A3(_06930_),
    .ZN(_07331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31431_ (.A1(_07329_),
    .A2(_07331_),
    .ZN(_07332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31432_ (.A1(_07327_),
    .A2(_07332_),
    .ZN(_07333_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31433_ (.A1(_06983_),
    .A2(_06946_),
    .B(_07126_),
    .ZN(_07334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31434_ (.A1(_07334_),
    .A2(_07009_),
    .B(_06893_),
    .ZN(_07335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31435_ (.A1(_07198_),
    .A2(_07053_),
    .ZN(_07336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31436_ (.A1(_06849_),
    .A2(_06954_),
    .ZN(_07337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31437_ (.A1(_07337_),
    .A2(_07336_),
    .A3(_06960_),
    .ZN(_07338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31438_ (.A1(_07338_),
    .A2(_07335_),
    .ZN(_07339_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31439_ (.A1(_07333_),
    .A2(_06952_),
    .A3(_07339_),
    .ZN(_07340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31440_ (.A1(_07340_),
    .A2(_07324_),
    .A3(_06873_),
    .ZN(_07342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31441_ (.A1(_07342_),
    .A2(_07311_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31442_ (.A1(_07054_),
    .A2(_06943_),
    .ZN(_07343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31443_ (.A1(_07343_),
    .A2(_07025_),
    .ZN(_07344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31444_ (.I(_16189_),
    .ZN(_07345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31445_ (.A1(_07345_),
    .A2(_06850_),
    .B(_06821_),
    .ZN(_07346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31446_ (.A1(_07346_),
    .A2(_07321_),
    .ZN(_07347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31447_ (.A1(_07344_),
    .A2(_07347_),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31448_ (.A1(_07348_),
    .A2(_06912_),
    .B(_06866_),
    .ZN(_07349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31449_ (.A1(_07248_),
    .A2(_06876_),
    .Z(_07350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31450_ (.A1(_07089_),
    .A2(_06982_),
    .ZN(_07351_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31451_ (.A1(_06921_),
    .A2(_07350_),
    .B(_07351_),
    .C(_06968_),
    .ZN(_07352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31452_ (.A1(_07349_),
    .A2(_07352_),
    .ZN(_07353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31453_ (.A1(_07037_),
    .A2(_06948_),
    .ZN(_07354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31454_ (.A1(_07012_),
    .A2(_06841_),
    .B(_06821_),
    .ZN(_07355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31455_ (.A1(_07355_),
    .A2(_07156_),
    .ZN(_07356_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31456_ (.A1(_07354_),
    .A2(_07356_),
    .A3(_06816_),
    .ZN(_07357_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31457_ (.A1(net18),
    .A2(_06841_),
    .B(_06821_),
    .ZN(_07358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31458_ (.A1(_07358_),
    .A2(_07207_),
    .B(_06843_),
    .ZN(_07359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31459_ (.A1(_07207_),
    .A2(_06986_),
    .ZN(_07360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31460_ (.A1(_07016_),
    .A2(_06898_),
    .ZN(_07362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31461_ (.A1(_07360_),
    .A2(_07362_),
    .A3(_07126_),
    .ZN(_07363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31462_ (.A1(_07359_),
    .A2(_07363_),
    .ZN(_07364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31463_ (.A1(_07357_),
    .A2(_07364_),
    .ZN(_07365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31464_ (.A1(_07365_),
    .A2(_06867_),
    .ZN(_07366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31465_ (.A1(_07353_),
    .A2(_07366_),
    .ZN(_07367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31466_ (.A1(_07367_),
    .A2(_06873_),
    .ZN(_07368_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31467_ (.A1(_16188_),
    .A2(_16197_),
    .Z(_07369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31468_ (.A1(_06905_),
    .A2(_07369_),
    .B(_06843_),
    .ZN(_07370_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31469_ (.A1(_07000_),
    .A2(_06975_),
    .A3(_06986_),
    .ZN(_07371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31470_ (.A1(_07370_),
    .A2(_07371_),
    .B(_06960_),
    .ZN(_07373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31471_ (.A1(_07132_),
    .A2(_06925_),
    .B(_07294_),
    .ZN(_07374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31472_ (.A1(_07296_),
    .A2(_07015_),
    .B(_06892_),
    .ZN(_07375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31473_ (.A1(_07374_),
    .A2(_07375_),
    .ZN(_07376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31474_ (.A1(_07373_),
    .A2(_07376_),
    .B(_06951_),
    .ZN(_07377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31475_ (.A1(_06908_),
    .A2(_06971_),
    .A3(_06843_),
    .ZN(_07378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31476_ (.A1(_06824_),
    .A2(_06986_),
    .A3(_06843_),
    .ZN(_07379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31477_ (.A1(_06904_),
    .A2(_06946_),
    .ZN(_07380_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31478_ (.A1(_07378_),
    .A2(_07379_),
    .A3(_07380_),
    .ZN(_07381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31479_ (.A1(_07140_),
    .A2(_07170_),
    .B(_06816_),
    .ZN(_07382_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31480_ (.A1(_07381_),
    .A2(_07382_),
    .B(_06880_),
    .ZN(_07384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31481_ (.A1(_07377_),
    .A2(_07384_),
    .B(_06873_),
    .ZN(_07385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31482_ (.A1(_07147_),
    .A2(_07058_),
    .A3(_07175_),
    .Z(_07386_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31483_ (.A1(_06929_),
    .A2(_06946_),
    .A3(_06932_),
    .ZN(_07387_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31484_ (.A1(_07270_),
    .A2(_07012_),
    .Z(_07388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31485_ (.A1(_07387_),
    .A2(_07388_),
    .B(_06960_),
    .ZN(_07389_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31486_ (.A1(_07386_),
    .A2(_07389_),
    .B(_06894_),
    .ZN(_07390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31487_ (.A1(_06878_),
    .A2(_06850_),
    .ZN(_07391_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31488_ (.A1(_07391_),
    .A2(_07024_),
    .Z(_07392_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31489_ (.A1(_07392_),
    .A2(_06886_),
    .A3(_07268_),
    .ZN(_07393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31490_ (.A1(_06958_),
    .A2(_06905_),
    .B(_06853_),
    .ZN(_07395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31491_ (.A1(_06971_),
    .A2(net81),
    .ZN(_07396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31492_ (.A1(_07396_),
    .A2(_06946_),
    .ZN(_07397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31493_ (.A1(_07395_),
    .A2(_07397_),
    .B(_06893_),
    .ZN(_07398_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31494_ (.A1(_07393_),
    .A2(_07398_),
    .B(_06866_),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31495_ (.A1(_07390_),
    .A2(_07399_),
    .ZN(_07400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31496_ (.A1(_07385_),
    .A2(_07400_),
    .ZN(_07401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31497_ (.A1(_07368_),
    .A2(_07401_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31498_ (.A1(_07114_),
    .A2(_07066_),
    .B(_07161_),
    .ZN(_07402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31499_ (.A1(_07402_),
    .A2(_06911_),
    .ZN(_07403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31500_ (.A1(_07133_),
    .A2(_06905_),
    .A3(_06896_),
    .ZN(_07405_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31501_ (.A1(_06958_),
    .A2(_06819_),
    .Z(_07406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31502_ (.A1(_07406_),
    .A2(_06982_),
    .A3(_07405_),
    .ZN(_07407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31503_ (.A1(_07403_),
    .A2(_07407_),
    .ZN(_07408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31504_ (.A1(_07408_),
    .A2(_06894_),
    .ZN(_07409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31505_ (.A1(_06919_),
    .A2(_06925_),
    .ZN(_07410_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _31506_ (.A1(_06921_),
    .A2(_07410_),
    .A3(_06906_),
    .A4(net905),
    .ZN(_07411_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31507_ (.A1(_07057_),
    .A2(_06926_),
    .ZN(_07412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31508_ (.A1(_07371_),
    .A2(_07412_),
    .B(_06912_),
    .ZN(_07413_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31509_ (.A1(_07411_),
    .A2(_07413_),
    .B(_06952_),
    .ZN(_07414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31510_ (.A1(_07409_),
    .A2(_07414_),
    .ZN(_07416_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31511_ (.I(_16183_),
    .ZN(_07417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31512_ (.A1(_07417_),
    .A2(_06946_),
    .B(_07126_),
    .ZN(_07418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31513_ (.A1(_07418_),
    .A2(_06906_),
    .B(_06816_),
    .ZN(_07419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31514_ (.A1(_07396_),
    .A2(_06930_),
    .ZN(_07420_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31515_ (.A1(_07001_),
    .A2(_06911_),
    .A3(_07420_),
    .ZN(_07421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31516_ (.A1(_07419_),
    .A2(_07421_),
    .B(_06866_),
    .ZN(_07422_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31517_ (.A1(_07181_),
    .A2(_06901_),
    .A3(_07012_),
    .Z(_07423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31518_ (.A1(_06939_),
    .A2(_06932_),
    .ZN(_07424_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31519_ (.A1(_06880_),
    .A2(_07424_),
    .A3(_07423_),
    .ZN(_07425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31520_ (.A1(_16197_),
    .A2(_06946_),
    .B(_07058_),
    .ZN(_07427_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31521_ (.A1(_07155_),
    .A2(_07181_),
    .B(_06905_),
    .ZN(_07428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31522_ (.A1(_07427_),
    .A2(_07428_),
    .B(_06912_),
    .ZN(_07429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31523_ (.A1(_07429_),
    .A2(_07425_),
    .ZN(_07430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31524_ (.A1(_07430_),
    .A2(_07422_),
    .B(_06873_),
    .ZN(_07431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31525_ (.A1(_07416_),
    .A2(_07431_),
    .ZN(_07432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31526_ (.A1(_07375_),
    .A2(_07124_),
    .ZN(_07433_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31527_ (.A1(_07016_),
    .A2(_06843_),
    .ZN(_07434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31528_ (.A1(_07434_),
    .A2(_07248_),
    .B(_06960_),
    .ZN(_07435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31529_ (.A1(_07433_),
    .A2(_07435_),
    .B(_06951_),
    .ZN(_07436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31530_ (.A1(_07022_),
    .A2(_06892_),
    .Z(_07438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31531_ (.A1(_06939_),
    .A2(_06878_),
    .ZN(_07439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31532_ (.A1(_07132_),
    .A2(_06925_),
    .ZN(_07440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31533_ (.A1(_07438_),
    .A2(_07439_),
    .A3(_07440_),
    .ZN(_07441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31534_ (.A1(_07167_),
    .A2(_06968_),
    .A3(_07040_),
    .ZN(_07442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31535_ (.A1(_07441_),
    .A2(_07442_),
    .A3(_06880_),
    .ZN(_07443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31536_ (.A1(_07443_),
    .A2(_07436_),
    .B(_06874_),
    .ZN(_07444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31537_ (.A1(_06980_),
    .A2(_06930_),
    .A3(_06932_),
    .ZN(_07445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31538_ (.A1(_07119_),
    .A2(_07445_),
    .ZN(_07446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31539_ (.A1(_06901_),
    .A2(_16169_),
    .ZN(_07447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31540_ (.A1(_07238_),
    .A2(_07447_),
    .ZN(_07449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31541_ (.A1(_07449_),
    .A2(_06880_),
    .ZN(_07450_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31542_ (.A1(_07446_),
    .A2(_07450_),
    .A3(_06894_),
    .ZN(_07451_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31543_ (.A1(_06994_),
    .A2(_06930_),
    .B(_07175_),
    .C(_06982_),
    .ZN(_07452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31544_ (.A1(_07198_),
    .A2(_06980_),
    .ZN(_07453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31545_ (.A1(_07453_),
    .A2(_07391_),
    .A3(_06960_),
    .ZN(_07454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31546_ (.A1(_07452_),
    .A2(_07454_),
    .A3(_06935_),
    .ZN(_07455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31547_ (.A1(_07451_),
    .A2(_06952_),
    .A3(_07455_),
    .ZN(_07456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31548_ (.A1(_07456_),
    .A2(_07444_),
    .ZN(_07457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31549_ (.A1(_07457_),
    .A2(_07432_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31550_ (.I(\dcnt[3] ),
    .ZN(_07459_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31551_ (.I(\dcnt[2] ),
    .ZN(_07460_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31552_ (.A1(_07459_),
    .A2(_07460_),
    .Z(_07461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31553_ (.I(\dcnt[1] ),
    .ZN(_07462_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _31554_ (.A1(_07461_),
    .A2(_07911_),
    .A3(_07462_),
    .A4(\dcnt[0] ),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31555_ (.A1(\u0.w[0][24] ),
    .A2(net75),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31556_ (.A1(net631),
    .A2(net620),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31557_ (.A1(\u0.w[0][26] ),
    .A2(\sa00_sr[2] ),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31558_ (.A1(\u0.w[0][27] ),
    .A2(\sa00_sr[3] ),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31559_ (.A1(\u0.w[0][28] ),
    .A2(\sa00_sr[4] ),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31560_ (.A1(\u0.w[0][29] ),
    .A2(\sa00_sr[5] ),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31561_ (.A1(\u0.w[0][30] ),
    .A2(\sa00_sr[6] ),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31562_ (.A1(\u0.w[0][31] ),
    .A2(net76),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31563_ (.A1(net700),
    .A2(\sa01_sr[0] ),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31564_ (.A1(net655),
    .A2(\sa01_sr[1] ),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31565_ (.A1(net768),
    .A2(\sa01_sr[2] ),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31566_ (.A1(\u0.w[1][27] ),
    .A2(\sa01_sr[3] ),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31567_ (.A1(\u0.w[1][28] ),
    .A2(\sa01_sr[4] ),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31568_ (.A1(\u0.w[1][29] ),
    .A2(\sa01_sr[5] ),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31569_ (.A1(\u0.w[1][30] ),
    .A2(\sa01_sr[6] ),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31570_ (.A1(\u0.w[1][31] ),
    .A2(net35),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31571_ (.A1(net490),
    .A2(net1176),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31572_ (.A1(net622),
    .A2(net1198),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31573_ (.A1(net709),
    .A2(\sa02_sr[2] ),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31574_ (.A1(\u0.w[2][27] ),
    .A2(\sa02_sr[3] ),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31575_ (.A1(\u0.w[2][28] ),
    .A2(\sa02_sr[4] ),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _31576_ (.A1(\u0.w[2][29] ),
    .A2(\sa02_sr[5] ),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31577_ (.A1(\u0.w[2][30] ),
    .A2(\sa02_sr[6] ),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31578_ (.A1(\u0.w[2][31] ),
    .A2(net57),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31579_ (.A1(\u0.tmp_w[24] ),
    .A2(net716),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31580_ (.A1(net628),
    .A2(net739),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31581_ (.A1(\u0.tmp_w[26] ),
    .A2(\sa03_sr[2] ),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31582_ (.A1(\u0.tmp_w[27] ),
    .A2(\sa03_sr[3] ),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31583_ (.A1(\u0.tmp_w[28] ),
    .A2(\sa03_sr[4] ),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31584_ (.A1(\u0.tmp_w[29] ),
    .A2(\sa03_sr[5] ),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31585_ (.A1(\u0.tmp_w[30] ),
    .A2(\sa03_sr[6] ),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31586_ (.A1(\u0.tmp_w[31] ),
    .A2(net39),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31587_ (.A1(\u0.w[0][16] ),
    .A2(net575),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31588_ (.A1(\u0.w[0][17] ),
    .A2(net493),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31589_ (.A1(\u0.w[0][18] ),
    .A2(net859),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31590_ (.A1(\u0.w[0][19] ),
    .A2(\sa10_sr[3] ),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31591_ (.A1(\u0.w[0][20] ),
    .A2(\sa10_sr[4] ),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31592_ (.A1(\u0.w[0][21] ),
    .A2(\sa10_sr[5] ),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31593_ (.A1(\u0.w[0][22] ),
    .A2(\sa10_sr[6] ),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31594_ (.A1(\u0.w[0][23] ),
    .A2(net46),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31595_ (.A1(\u0.w[1][16] ),
    .A2(net795),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31596_ (.A1(net1032),
    .A2(net806),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31597_ (.A1(\u0.w[1][18] ),
    .A2(\sa11_sr[2] ),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31598_ (.A1(\u0.w[1][19] ),
    .A2(\sa11_sr[3] ),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31599_ (.A1(\u0.w[1][20] ),
    .A2(\sa11_sr[4] ),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31600_ (.A1(\u0.w[1][21] ),
    .A2(\sa11_sr[5] ),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31601_ (.A1(\u0.w[1][22] ),
    .A2(\sa11_sr[6] ),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31602_ (.A1(\u0.w[1][23] ),
    .A2(net525),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31603_ (.A1(\u0.w[2][16] ),
    .A2(net1180),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31604_ (.A1(\u0.w[2][17] ),
    .A2(\sa12_sr[1] ),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31605_ (.A1(\u0.w[2][18] ),
    .A2(\sa12_sr[2] ),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31606_ (.A1(\u0.w[2][19] ),
    .A2(\sa12_sr[3] ),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31607_ (.A1(\u0.w[2][20] ),
    .A2(\sa12_sr[4] ),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31608_ (.A1(\u0.w[2][21] ),
    .A2(\sa12_sr[5] ),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31609_ (.A1(\u0.w[2][22] ),
    .A2(\sa12_sr[6] ),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31610_ (.A1(\u0.w[2][23] ),
    .A2(net72),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31611_ (.A1(\u0.tmp_w[16] ),
    .A2(\sa10_sub[0] ),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31612_ (.A1(\u0.tmp_w[17] ),
    .A2(net733),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31613_ (.A1(\u0.tmp_w[18] ),
    .A2(\sa10_sub[2] ),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31614_ (.A1(\u0.tmp_w[19] ),
    .A2(\sa10_sub[3] ),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31615_ (.A1(\u0.tmp_w[20] ),
    .A2(\sa10_sub[4] ),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31616_ (.A1(\u0.tmp_w[21] ),
    .A2(\sa10_sub[5] ),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31617_ (.A1(\u0.tmp_w[22] ),
    .A2(\sa10_sub[6] ),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31618_ (.A1(\u0.tmp_w[23] ),
    .A2(net772),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31619_ (.A1(\u0.w[0][8] ),
    .A2(net573),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31620_ (.A1(\u0.w[0][9] ),
    .A2(net613),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31621_ (.A1(\u0.w[0][10] ),
    .A2(\sa20_sr[2] ),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31622_ (.A1(\u0.w[0][11] ),
    .A2(\sa20_sr[3] ),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31623_ (.A1(\u0.w[0][12] ),
    .A2(\sa20_sr[4] ),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31624_ (.A1(\u0.w[0][13] ),
    .A2(\sa20_sr[5] ),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31625_ (.A1(\u0.w[0][14] ),
    .A2(\sa20_sr[6] ),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31626_ (.A1(\u0.w[0][15] ),
    .A2(net47),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _31627_ (.A1(\u0.w[1][8] ),
    .A2(net815),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31628_ (.A1(\u0.w[1][9] ),
    .A2(\sa21_sr[1] ),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31629_ (.A1(\u0.w[1][10] ),
    .A2(_11218_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31630_ (.A1(\u0.w[1][11] ),
    .A2(\sa21_sr[3] ),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31631_ (.A1(\u0.w[1][12] ),
    .A2(\sa21_sr[4] ),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31632_ (.A1(\u0.w[1][13] ),
    .A2(\sa21_sr[5] ),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31633_ (.A1(\u0.w[1][14] ),
    .A2(\sa21_sr[6] ),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31634_ (.A1(\u0.w[1][15] ),
    .A2(net26),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31635_ (.A1(\u0.w[2][8] ),
    .A2(\sa20_sub[0] ),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31636_ (.A1(\u0.w[2][9] ),
    .A2(net1169),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31637_ (.A1(\u0.w[2][10] ),
    .A2(_12027_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31638_ (.A1(\u0.w[2][11] ),
    .A2(\sa20_sub[3] ),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31639_ (.A1(\u0.w[2][12] ),
    .A2(\sa20_sub[4] ),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31640_ (.A1(\u0.w[2][13] ),
    .A2(\sa20_sub[5] ),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31641_ (.A1(\u0.w[2][14] ),
    .A2(\sa20_sub[6] ),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31642_ (.A1(\u0.w[2][15] ),
    .A2(net49),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31643_ (.A1(\u0.tmp_w[8] ),
    .A2(\sa21_sub[0] ),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31644_ (.A1(\u0.tmp_w[9] ),
    .A2(net528),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31645_ (.A1(\u0.tmp_w[10] ),
    .A2(_12836_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31646_ (.A1(\u0.tmp_w[11] ),
    .A2(\sa21_sub[3] ),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31647_ (.A1(\u0.tmp_w[12] ),
    .A2(\sa21_sub[4] ),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31648_ (.A1(\u0.tmp_w[13] ),
    .A2(\sa21_sub[5] ),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31649_ (.A1(\u0.tmp_w[14] ),
    .A2(\sa21_sub[6] ),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31650_ (.A1(\u0.tmp_w[15] ),
    .A2(net50),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31651_ (.A1(\u0.w[0][0] ),
    .A2(net584),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31652_ (.A1(\u0.w[0][1] ),
    .A2(net605),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31653_ (.A1(\u0.w[0][2] ),
    .A2(\sa30_sr[2] ),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31654_ (.A1(\u0.w[0][3] ),
    .A2(\sa30_sr[3] ),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31655_ (.A1(\u0.w[0][4] ),
    .A2(\sa30_sr[4] ),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31656_ (.A1(\u0.w[0][5] ),
    .A2(\sa30_sr[5] ),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31657_ (.A1(\u0.w[0][6] ),
    .A2(\sa30_sr[6] ),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31658_ (.A1(\u0.w[0][7] ),
    .A2(net68),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31659_ (.A1(\u0.w[1][0] ),
    .A2(net519),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31660_ (.A1(\u0.w[1][1] ),
    .A2(net1029),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31661_ (.A1(\u0.w[1][2] ),
    .A2(\sa30_sub[2] ),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31662_ (.A1(\u0.w[1][3] ),
    .A2(\sa30_sub[3] ),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31663_ (.A1(\u0.w[1][4] ),
    .A2(\sa30_sub[4] ),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31664_ (.A1(\u0.w[1][5] ),
    .A2(\sa30_sub[5] ),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31665_ (.A1(\u0.w[1][6] ),
    .A2(\sa30_sub[6] ),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31666_ (.A1(\u0.w[1][7] ),
    .A2(net819),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31667_ (.A1(\u0.w[2][0] ),
    .A2(\sa31_sub[0] ),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31668_ (.A1(\u0.w[2][1] ),
    .A2(\sa31_sub[1] ),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31669_ (.A1(\u0.w[2][2] ),
    .A2(\sa31_sub[2] ),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31670_ (.A1(\u0.w[2][3] ),
    .A2(\sa31_sub[3] ),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31671_ (.A1(\u0.w[2][4] ),
    .A2(\sa31_sub[4] ),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31672_ (.A1(\u0.w[2][5] ),
    .A2(\sa31_sub[5] ),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _31673_ (.A1(\u0.w[2][6] ),
    .A2(\sa31_sub[6] ),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31674_ (.A1(\u0.w[2][7] ),
    .A2(net642),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31675_ (.A1(\u0.tmp_w[0] ),
    .A2(\sa32_sub[0] ),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31676_ (.A1(\u0.tmp_w[1] ),
    .A2(net38),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31677_ (.A1(\u0.tmp_w[2] ),
    .A2(\sa32_sub[2] ),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31678_ (.A1(\u0.tmp_w[3] ),
    .A2(\sa32_sub[3] ),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31679_ (.A1(\u0.tmp_w[4] ),
    .A2(\sa32_sub[4] ),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31680_ (.A1(\u0.tmp_w[5] ),
    .A2(\sa32_sub[5] ),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31681_ (.A1(\u0.tmp_w[6] ),
    .A2(\sa32_sub[6] ),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31682_ (.A1(\u0.tmp_w[7] ),
    .A2(net54),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31683_ (.I(\u0.r0.rcnt[0] ),
    .ZN(\u0.r0.rcnt_next[0] ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31684_ (.I(\u0.r0.rcnt[1] ),
    .ZN(_16201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31685_ (.I0(\text_in_r[0] ),
    .I1(net218),
    .S(_07774_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31686_ (.I(_07773_),
    .Z(_07474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31687_ (.I0(\text_in_r[100] ),
    .I1(net219),
    .S(_07474_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31688_ (.I0(\text_in_r[101] ),
    .I1(net220),
    .S(_07474_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31689_ (.I0(\text_in_r[102] ),
    .I1(net221),
    .S(_07474_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31690_ (.I0(\text_in_r[103] ),
    .I1(net222),
    .S(_07474_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31691_ (.I0(\text_in_r[104] ),
    .I1(net223),
    .S(_07474_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31692_ (.I0(\text_in_r[105] ),
    .I1(net224),
    .S(_07474_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31693_ (.I0(\text_in_r[106] ),
    .I1(net225),
    .S(_07474_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31694_ (.I0(\text_in_r[107] ),
    .I1(net226),
    .S(_07474_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31695_ (.I0(\text_in_r[108] ),
    .I1(net227),
    .S(_07474_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31696_ (.I0(\text_in_r[109] ),
    .I1(net228),
    .S(_07474_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31697_ (.I(_07773_),
    .Z(_07476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31698_ (.I0(\text_in_r[10] ),
    .I1(net229),
    .S(_07476_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31699_ (.I0(\text_in_r[110] ),
    .I1(net230),
    .S(_07476_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31700_ (.I0(\text_in_r[111] ),
    .I1(net231),
    .S(_07476_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31701_ (.I0(\text_in_r[112] ),
    .I1(net232),
    .S(_07476_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31702_ (.I0(\text_in_r[113] ),
    .I1(net233),
    .S(_07476_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31703_ (.I0(\text_in_r[114] ),
    .I1(net234),
    .S(_07476_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31704_ (.I0(\text_in_r[115] ),
    .I1(net235),
    .S(_07476_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31705_ (.I0(\text_in_r[116] ),
    .I1(net236),
    .S(_07476_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31706_ (.I0(\text_in_r[117] ),
    .I1(net237),
    .S(_07476_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31707_ (.I0(\text_in_r[118] ),
    .I1(net238),
    .S(_07476_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31708_ (.I(_07773_),
    .Z(_07478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31709_ (.I0(\text_in_r[119] ),
    .I1(net239),
    .S(_07478_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31710_ (.I0(\text_in_r[11] ),
    .I1(net240),
    .S(_07478_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31711_ (.I0(\text_in_r[120] ),
    .I1(net241),
    .S(_07478_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31712_ (.I0(\text_in_r[121] ),
    .I1(net242),
    .S(_07478_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31713_ (.I0(\text_in_r[122] ),
    .I1(net243),
    .S(_07478_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31714_ (.I0(\text_in_r[123] ),
    .I1(net244),
    .S(_07478_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31715_ (.I0(\text_in_r[124] ),
    .I1(net245),
    .S(_07478_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31716_ (.I0(\text_in_r[125] ),
    .I1(net246),
    .S(_07478_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31717_ (.I0(\text_in_r[126] ),
    .I1(net247),
    .S(_07478_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31718_ (.I0(\text_in_r[127] ),
    .I1(net248),
    .S(_07478_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31719_ (.I(_07773_),
    .Z(_07480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31720_ (.I0(\text_in_r[12] ),
    .I1(net249),
    .S(_07480_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31721_ (.I0(\text_in_r[13] ),
    .I1(net250),
    .S(_07480_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31722_ (.I0(\text_in_r[14] ),
    .I1(net251),
    .S(_07480_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31723_ (.I0(\text_in_r[15] ),
    .I1(net252),
    .S(_07480_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31724_ (.I0(\text_in_r[16] ),
    .I1(net253),
    .S(_07480_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31725_ (.I0(\text_in_r[17] ),
    .I1(net254),
    .S(_07480_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31726_ (.I0(\text_in_r[18] ),
    .I1(net255),
    .S(_07480_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31727_ (.I0(\text_in_r[19] ),
    .I1(net256),
    .S(_07480_),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31728_ (.I0(\text_in_r[1] ),
    .I1(net257),
    .S(_07480_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31729_ (.I0(\text_in_r[20] ),
    .I1(net258),
    .S(_07480_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31730_ (.I(_07773_),
    .Z(_07483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31731_ (.I0(\text_in_r[21] ),
    .I1(net259),
    .S(_07483_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31732_ (.I0(\text_in_r[22] ),
    .I1(net260),
    .S(_07483_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31733_ (.I0(\text_in_r[23] ),
    .I1(net261),
    .S(_07483_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31734_ (.I0(\text_in_r[24] ),
    .I1(net262),
    .S(_07483_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31735_ (.I0(\text_in_r[25] ),
    .I1(net263),
    .S(_07483_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31736_ (.I0(\text_in_r[26] ),
    .I1(net264),
    .S(_07483_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31737_ (.I0(\text_in_r[27] ),
    .I1(net265),
    .S(_07483_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31738_ (.I0(\text_in_r[28] ),
    .I1(net266),
    .S(_07483_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31739_ (.I0(\text_in_r[29] ),
    .I1(net267),
    .S(_07483_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31740_ (.I0(\text_in_r[2] ),
    .I1(net268),
    .S(_07483_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31741_ (.I(_07773_),
    .Z(_07485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31742_ (.I0(\text_in_r[30] ),
    .I1(net269),
    .S(_07485_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31743_ (.I0(\text_in_r[31] ),
    .I1(net270),
    .S(_07485_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31744_ (.I0(\text_in_r[32] ),
    .I1(net271),
    .S(_07485_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31745_ (.I0(\text_in_r[33] ),
    .I1(net272),
    .S(_07485_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31746_ (.I0(\text_in_r[34] ),
    .I1(net273),
    .S(_07485_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31747_ (.I0(\text_in_r[35] ),
    .I1(net274),
    .S(_07485_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31748_ (.I0(\text_in_r[36] ),
    .I1(net275),
    .S(_07485_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31749_ (.I0(\text_in_r[37] ),
    .I1(net276),
    .S(_07485_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31750_ (.I0(\text_in_r[38] ),
    .I1(net277),
    .S(_07485_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31751_ (.I0(\text_in_r[39] ),
    .I1(net278),
    .S(_07485_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _31752_ (.I(_07773_),
    .Z(_07487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31753_ (.I0(\text_in_r[3] ),
    .I1(net279),
    .S(_07487_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31754_ (.I0(\text_in_r[40] ),
    .I1(net280),
    .S(_07487_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31755_ (.I0(\text_in_r[41] ),
    .I1(net281),
    .S(_07487_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31756_ (.I0(\text_in_r[42] ),
    .I1(net282),
    .S(_07487_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31757_ (.I0(\text_in_r[43] ),
    .I1(net283),
    .S(_07487_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31758_ (.I0(\text_in_r[44] ),
    .I1(net284),
    .S(_07487_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31759_ (.I0(\text_in_r[45] ),
    .I1(net285),
    .S(_07487_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31760_ (.I0(\text_in_r[46] ),
    .I1(net286),
    .S(_07487_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31761_ (.I0(\text_in_r[47] ),
    .I1(net287),
    .S(_07487_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31762_ (.I0(\text_in_r[48] ),
    .I1(net288),
    .S(_07487_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31763_ (.I(_07773_),
    .Z(_07488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31764_ (.I0(\text_in_r[49] ),
    .I1(net289),
    .S(_07488_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31765_ (.I0(\text_in_r[4] ),
    .I1(net290),
    .S(_07488_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31766_ (.I0(\text_in_r[50] ),
    .I1(net291),
    .S(_07488_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31767_ (.I0(\text_in_r[51] ),
    .I1(net292),
    .S(_07488_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31768_ (.I0(\text_in_r[52] ),
    .I1(net293),
    .S(_07488_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31769_ (.I0(\text_in_r[53] ),
    .I1(net294),
    .S(_07488_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31770_ (.I0(\text_in_r[54] ),
    .I1(net295),
    .S(_07488_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31771_ (.I0(\text_in_r[55] ),
    .I1(net296),
    .S(_07488_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31772_ (.I0(\text_in_r[56] ),
    .I1(net297),
    .S(_07488_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31773_ (.I0(\text_in_r[57] ),
    .I1(net298),
    .S(_07488_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31774_ (.I(_07773_),
    .Z(_07490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31775_ (.I0(\text_in_r[58] ),
    .I1(net299),
    .S(_07490_),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31776_ (.I0(\text_in_r[59] ),
    .I1(net300),
    .S(_07490_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31777_ (.I0(\text_in_r[5] ),
    .I1(net301),
    .S(_07490_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31778_ (.I0(\text_in_r[60] ),
    .I1(net302),
    .S(_07490_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31779_ (.I0(\text_in_r[61] ),
    .I1(net303),
    .S(_07490_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31780_ (.I0(\text_in_r[62] ),
    .I1(net304),
    .S(_07490_),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31781_ (.I0(\text_in_r[63] ),
    .I1(net305),
    .S(_07490_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31782_ (.I0(\text_in_r[64] ),
    .I1(net306),
    .S(_07490_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31783_ (.I0(\text_in_r[65] ),
    .I1(net307),
    .S(_07490_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31784_ (.I0(\text_in_r[66] ),
    .I1(net308),
    .S(_07490_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _31785_ (.I(_07789_),
    .Z(_07492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31786_ (.I0(\text_in_r[67] ),
    .I1(net309),
    .S(_07492_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31787_ (.I0(\text_in_r[68] ),
    .I1(net310),
    .S(_07492_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31788_ (.I0(\text_in_r[69] ),
    .I1(net311),
    .S(_07492_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31789_ (.I0(\text_in_r[6] ),
    .I1(net312),
    .S(_07492_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31790_ (.I0(\text_in_r[70] ),
    .I1(net313),
    .S(_07492_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31791_ (.I0(\text_in_r[71] ),
    .I1(net314),
    .S(_07492_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31792_ (.I0(\text_in_r[72] ),
    .I1(net315),
    .S(_07492_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31793_ (.I0(\text_in_r[73] ),
    .I1(net316),
    .S(_07492_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31794_ (.I0(\text_in_r[74] ),
    .I1(net317),
    .S(_07492_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31795_ (.I0(\text_in_r[75] ),
    .I1(net318),
    .S(_07492_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _31796_ (.I(_07789_),
    .Z(_07494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31797_ (.I0(\text_in_r[76] ),
    .I1(net319),
    .S(_07494_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31798_ (.I0(\text_in_r[77] ),
    .I1(net320),
    .S(_07494_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31799_ (.I0(\text_in_r[78] ),
    .I1(net321),
    .S(_07494_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31800_ (.I0(\text_in_r[79] ),
    .I1(net322),
    .S(_07494_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31801_ (.I0(\text_in_r[7] ),
    .I1(net323),
    .S(_07494_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31802_ (.I0(\text_in_r[80] ),
    .I1(net324),
    .S(_07494_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31803_ (.I0(\text_in_r[81] ),
    .I1(net325),
    .S(_07494_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31804_ (.I0(\text_in_r[82] ),
    .I1(net326),
    .S(_07494_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31805_ (.I0(\text_in_r[83] ),
    .I1(net327),
    .S(_07494_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31806_ (.I0(\text_in_r[84] ),
    .I1(net328),
    .S(_07494_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _31807_ (.I(_07789_),
    .Z(_07496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31808_ (.I0(\text_in_r[85] ),
    .I1(net329),
    .S(_07496_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31809_ (.I0(\text_in_r[86] ),
    .I1(net330),
    .S(_07496_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31810_ (.I0(\text_in_r[87] ),
    .I1(net331),
    .S(_07496_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31811_ (.I0(\text_in_r[88] ),
    .I1(net332),
    .S(_07496_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31812_ (.I0(\text_in_r[89] ),
    .I1(net333),
    .S(_07496_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31813_ (.I0(\text_in_r[8] ),
    .I1(net334),
    .S(_07496_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31814_ (.I0(\text_in_r[90] ),
    .I1(net335),
    .S(_07496_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31815_ (.I0(\text_in_r[91] ),
    .I1(net336),
    .S(_07496_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31816_ (.I0(\text_in_r[92] ),
    .I1(net337),
    .S(_07496_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31817_ (.I0(\text_in_r[93] ),
    .I1(net338),
    .S(_07496_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31818_ (.I0(\text_in_r[94] ),
    .I1(net339),
    .S(_07942_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31819_ (.I0(\text_in_r[95] ),
    .I1(net340),
    .S(_07942_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31820_ (.I0(\text_in_r[96] ),
    .I1(net341),
    .S(_07942_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31821_ (.I0(\text_in_r[97] ),
    .I1(net342),
    .S(_07942_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31822_ (.I0(\text_in_r[98] ),
    .I1(net343),
    .S(_07942_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31823_ (.I0(\text_in_r[99] ),
    .I1(net344),
    .S(_07942_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31824_ (.I0(\text_in_r[9] ),
    .I1(net345),
    .S(_07942_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31825_ (.A1(\dcnt[1] ),
    .A2(\dcnt[0] ),
    .ZN(_07499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31826_ (.A1(_07461_),
    .A2(_07499_),
    .ZN(_07500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31827_ (.A1(_07500_),
    .A2(net217),
    .ZN(_07501_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31828_ (.A1(_07499_),
    .A2(_07460_),
    .Z(_07502_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31829_ (.A1(_07499_),
    .A2(_07460_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31830_ (.A1(_07502_),
    .A2(_07503_),
    .ZN(_07505_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31831_ (.A1(_07501_),
    .A2(_07505_),
    .A3(_07747_),
    .Z(_07506_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31832_ (.I(_07506_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31833_ (.A1(\u0.r0.rcnt[2] ),
    .A2(_16209_),
    .Z(_07507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31834_ (.A1(\u0.r0.rcnt[2] ),
    .A2(_16209_),
    .ZN(_07508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31835_ (.A1(_07507_),
    .A2(_07508_),
    .ZN(_07509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31836_ (.A1(_07509_),
    .A2(_16207_),
    .Z(_07510_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31837_ (.A1(_07510_),
    .A2(_07940_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31838_ (.A1(\u0.r0.rcnt[2] ),
    .A2(\u0.r0.rcnt[1] ),
    .A3(\u0.r0.rcnt[0] ),
    .ZN(_07511_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31839_ (.A1(\u0.r0.rcnt[3] ),
    .A2(_07511_),
    .Z(_07512_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31840_ (.I(_07512_),
    .ZN(_07514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31841_ (.I(_16202_),
    .ZN(_07515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31842_ (.I(_07509_),
    .ZN(_07516_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31843_ (.A1(_07514_),
    .A2(_07515_),
    .A3(_07516_),
    .Z(_07517_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31844_ (.A1(_07512_),
    .A2(\u0.r0.rcnt_next[1] ),
    .A3(_07516_),
    .Z(_07518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31845_ (.A1(_07517_),
    .A2(_07518_),
    .B(_07940_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31846_ (.A1(_07512_),
    .A2(_07515_),
    .A3(_07516_),
    .Z(_07519_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31847_ (.A1(_07512_),
    .A2(_16205_),
    .A3(_07509_),
    .ZN(_07520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31848_ (.A1(_07519_),
    .A2(_07520_),
    .B(_07940_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31849_ (.A1(_07512_),
    .A2(_16203_),
    .A3(_07509_),
    .ZN(_07521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31850_ (.A1(_07514_),
    .A2(_07510_),
    .ZN(_07522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31851_ (.A1(_07521_),
    .A2(_07522_),
    .B(_07940_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31852_ (.A1(_07512_),
    .A2(_07516_),
    .Z(_07523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31853_ (.A1(_07523_),
    .A2(_16207_),
    .ZN(_07524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31854_ (.A1(_07518_),
    .A2(_07524_),
    .B(_07940_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31855_ (.A1(_07523_),
    .A2(_16202_),
    .ZN(_07525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31856_ (.A1(_07519_),
    .A2(_07525_),
    .B(_07940_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31857_ (.A1(_07523_),
    .A2(_07911_),
    .A3(_16205_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31858_ (.A1(_07523_),
    .A2(_07911_),
    .A3(_16203_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31859_ (.A1(_07911_),
    .A2(\u0.r0.rcnt_next[0] ),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31860_ (.A1(_07911_),
    .A2(\u0.r0.rcnt_next[1] ),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31861_ (.A1(_07516_),
    .A2(_07911_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31862_ (.A1(_07514_),
    .A2(_07911_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31863_ (.A1(_07747_),
    .A2(net217),
    .ZN(_07527_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31864_ (.A1(_07501_),
    .A2(\dcnt[0] ),
    .B(_07527_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31865_ (.A1(_07461_),
    .A2(\dcnt[1] ),
    .A3(\dcnt[0] ),
    .Z(_07528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31866_ (.A1(\dcnt[1] ),
    .A2(\dcnt[0] ),
    .B(_07747_),
    .ZN(_07529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31867_ (.I(net217),
    .ZN(_07530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31868_ (.A1(_07528_),
    .A2(_07529_),
    .B(_07530_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _31869_ (.A1(_07502_),
    .A2(_07530_),
    .A3(_07459_),
    .B(_07527_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31870_ (.A(_15537_),
    .B(_15538_),
    .CO(_15539_),
    .S(_15540_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31871_ (.A(_15537_),
    .B(_15538_),
    .CO(_15541_),
    .S(_15542_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31872_ (.A(_15537_),
    .B(_15543_),
    .CO(_15544_),
    .S(_15545_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31873_ (.A(_15537_),
    .B(_15543_),
    .CO(_15546_),
    .S(_15547_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31874_ (.A(_15548_),
    .B(_15538_),
    .CO(_15549_),
    .S(_15550_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31875_ (.A(_15548_),
    .B(_15538_),
    .CO(_15551_),
    .S(_15552_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31876_ (.A(_15548_),
    .B(_15543_),
    .CO(_15553_),
    .S(_15554_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31877_ (.A(_15548_),
    .B(_15543_),
    .CO(_15555_),
    .S(_15556_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31878_ (.A(net895),
    .B(_15557_),
    .CO(_15558_),
    .S(_15559_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31879_ (.A(net6),
    .B(_15557_),
    .CO(_15560_),
    .S(_15561_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31880_ (.A(net6),
    .B(_15562_),
    .CO(_15563_),
    .S(_15564_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31881_ (.A(net6),
    .B(_15562_),
    .CO(_15565_),
    .S(_15566_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31882_ (.A(net82),
    .B(_15557_),
    .CO(_15567_),
    .S(_15568_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31883_ (.A(net82),
    .B(_15557_),
    .CO(_15569_),
    .S(_15570_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31884_ (.A(_15572_),
    .B(_15571_),
    .CO(_15573_),
    .S(_15574_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31885_ (.A(_15571_),
    .B(_15572_),
    .CO(_15575_),
    .S(_15576_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31886_ (.A(_15571_),
    .B(_15577_),
    .CO(_15578_),
    .S(_15579_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31887_ (.A(_15571_),
    .B(_15577_),
    .CO(_15580_),
    .S(_15581_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31888_ (.A(_15582_),
    .B(_15572_),
    .CO(_15583_),
    .S(_15584_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31889_ (.A(_15582_),
    .B(_15572_),
    .CO(_15585_),
    .S(_15586_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31890_ (.A(_15582_),
    .B(_15577_),
    .CO(_15587_),
    .S(_15588_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31891_ (.A(_15582_),
    .B(_15577_),
    .CO(_15589_),
    .S(_15590_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31892_ (.A(_15571_),
    .B(_15591_),
    .CO(_15592_),
    .S(_15593_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31893_ (.A(_15571_),
    .B(_15591_),
    .CO(_15594_),
    .S(_15595_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31894_ (.A(net30),
    .B(_15596_),
    .CO(_15597_),
    .S(_15598_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31895_ (.A(_15571_),
    .B(_15596_),
    .CO(_15599_),
    .S(_15600_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31896_ (.A(net78),
    .B(_15591_),
    .CO(_15601_),
    .S(_15602_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31897_ (.A(net78),
    .B(_15591_),
    .CO(_15603_),
    .S(_15604_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31898_ (.A(_15606_),
    .B(_15605_),
    .CO(_15607_),
    .S(_15608_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31899_ (.A(_15605_),
    .B(_15606_),
    .CO(_15609_),
    .S(_15610_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31900_ (.A(_15605_),
    .B(_15611_),
    .CO(_15612_),
    .S(_15613_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31901_ (.A(_15605_),
    .B(_15611_),
    .CO(_15614_),
    .S(_15615_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31902_ (.A(_15616_),
    .B(_15606_),
    .CO(_15617_),
    .S(_15618_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31903_ (.A(_15616_),
    .B(_15606_),
    .CO(_15619_),
    .S(_15620_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31904_ (.A(_15616_),
    .B(_15611_),
    .CO(_15621_),
    .S(_15622_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31905_ (.A(_15616_),
    .B(_15611_),
    .CO(_15623_),
    .S(_15624_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31906_ (.A(_15605_),
    .B(_15625_),
    .CO(_15626_),
    .S(_15627_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31907_ (.A(_15605_),
    .B(_15625_),
    .CO(_15628_),
    .S(_15629_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31908_ (.A(net86),
    .B(_15630_),
    .CO(_15631_),
    .S(_15632_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31909_ (.A(_15605_),
    .B(_15630_),
    .CO(_15633_),
    .S(_15634_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31910_ (.A(net89),
    .B(_15625_),
    .CO(_15635_),
    .S(_15636_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31911_ (.A(_15616_),
    .B(_15625_),
    .CO(_15637_),
    .S(_15638_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31912_ (.A(_15639_),
    .B(_15640_),
    .CO(_15641_),
    .S(_15642_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31913_ (.A(net762),
    .B(_15640_),
    .CO(_15643_),
    .S(_15644_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31914_ (.A(net762),
    .B(net962),
    .CO(_15646_),
    .S(_15647_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31915_ (.A(net762),
    .B(net962),
    .CO(_15648_),
    .S(_15649_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31916_ (.A(net480),
    .B(_15640_),
    .CO(_15651_),
    .S(_15652_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31917_ (.A(net482),
    .B(net625),
    .CO(_15653_),
    .S(_15654_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31918_ (.A(net482),
    .B(net962),
    .CO(_15655_),
    .S(_15656_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31919_ (.A(net482),
    .B(net962),
    .CO(_15657_),
    .S(_15658_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31920_ (.A(net763),
    .B(_15659_),
    .CO(_15660_),
    .S(_15661_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31921_ (.A(_15659_),
    .B(_15639_),
    .CO(_15662_),
    .S(_15663_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31922_ (.A(_15664_),
    .B(net37),
    .CO(_15665_),
    .S(_15666_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31923_ (.A(_15664_),
    .B(net762),
    .CO(_15667_),
    .S(_15668_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31924_ (.A(_15664_),
    .B(net11),
    .CO(_15669_),
    .S(_15670_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31925_ (.A(_15664_),
    .B(net11),
    .CO(_15671_),
    .S(_15672_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31926_ (.A(_15674_),
    .B(_15673_),
    .CO(_15675_),
    .S(_15676_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31927_ (.A(_15673_),
    .B(_15674_),
    .CO(_15677_),
    .S(_15678_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31928_ (.A(net1260),
    .B(_15673_),
    .CO(_15680_),
    .S(_15681_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31929_ (.A(net828),
    .B(net610),
    .CO(_15683_),
    .S(_15684_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31930_ (.A(_15682_),
    .B(_15674_),
    .CO(_15685_),
    .S(_15686_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31931_ (.A(net600),
    .B(net828),
    .CO(_15687_),
    .S(_15688_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31932_ (.A(net828),
    .B(net1259),
    .CO(_15689_),
    .S(_15690_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31933_ (.A(_15691_),
    .B(net612),
    .CO(_15692_),
    .S(_15693_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31934_ (.A(_15691_),
    .B(net32),
    .CO(_15694_),
    .S(_15695_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31935_ (.A(_15691_),
    .B(net602),
    .CO(_15696_),
    .S(_15697_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31936_ (.A(_15698_),
    .B(net1263),
    .CO(_15699_),
    .S(_15700_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31937_ (.A(_15698_),
    .B(net1264),
    .CO(_15701_),
    .S(_15702_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31938_ (.A(_15698_),
    .B(net32),
    .CO(_15703_),
    .S(_15704_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31939_ (.A(_15705_),
    .B(_15706_),
    .CO(_15707_),
    .S(_15708_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31940_ (.A(net842),
    .B(_15706_),
    .CO(_15709_),
    .S(_15710_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31941_ (.A(net845),
    .B(_15711_),
    .CO(_15712_),
    .S(_15713_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31942_ (.A(_15714_),
    .B(net1024),
    .CO(_15715_),
    .S(_15716_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31943_ (.A(_15714_),
    .B(_15706_),
    .CO(_15717_),
    .S(_15718_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31944_ (.A(_15714_),
    .B(_15711_),
    .CO(_15719_),
    .S(_15720_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31945_ (.A(_15714_),
    .B(_15711_),
    .CO(_15721_),
    .S(_15722_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31946_ (.A(_15723_),
    .B(net1024),
    .CO(_15724_),
    .S(_15725_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31947_ (.A(_15723_),
    .B(_15711_),
    .CO(_15726_),
    .S(_15727_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31948_ (.A(_15723_),
    .B(_15711_),
    .CO(_15728_),
    .S(_15729_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31949_ (.A(_15730_),
    .B(net1),
    .CO(_15731_),
    .S(_15732_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31950_ (.A(_15730_),
    .B(net1024),
    .CO(_15733_),
    .S(_15734_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31951_ (.A(_15730_),
    .B(net42),
    .CO(_15735_),
    .S(_15736_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31952_ (.A(_15737_),
    .B(_15738_),
    .CO(_15739_),
    .S(_15740_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31953_ (.A(_15738_),
    .B(_15737_),
    .CO(_15741_),
    .S(_15742_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31954_ (.A(_15737_),
    .B(_15743_),
    .CO(_15744_),
    .S(_15745_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31955_ (.A(net1150),
    .B(_15738_),
    .CO(_15747_),
    .S(_15748_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31956_ (.A(_15746_),
    .B(_15738_),
    .CO(_15749_),
    .S(_15750_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31957_ (.A(net1150),
    .B(_15743_),
    .CO(_15751_),
    .S(_15752_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31958_ (.A(net1150),
    .B(_15743_),
    .CO(_15753_),
    .S(_15754_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31959_ (.A(_15755_),
    .B(net1162),
    .CO(_15756_),
    .S(_15757_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31960_ (.A(_15755_),
    .B(_15743_),
    .CO(_15758_),
    .S(_15759_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31961_ (.A(_15755_),
    .B(_15743_),
    .CO(_15760_),
    .S(_15761_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31962_ (.A(_15762_),
    .B(net17),
    .CO(_15763_),
    .S(_15764_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31963_ (.A(_15762_),
    .B(net1162),
    .CO(_15765_),
    .S(_15766_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31964_ (.A(_15762_),
    .B(_15743_),
    .CO(_15767_),
    .S(_15768_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31965_ (.A(_15769_),
    .B(_15770_),
    .CO(_15771_),
    .S(_15772_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31966_ (.A(net549),
    .B(net968),
    .CO(_15773_),
    .S(_15774_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31967_ (.A(_15775_),
    .B(net549),
    .CO(_15776_),
    .S(_15777_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31968_ (.A(net542),
    .B(net486),
    .CO(_15779_),
    .S(_15780_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31969_ (.A(net486),
    .B(net540),
    .CO(_15781_),
    .S(_15782_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31970_ (.A(net538),
    .B(net41),
    .CO(_15783_),
    .S(_15784_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31971_ (.A(net542),
    .B(_15775_),
    .CO(_15785_),
    .S(_15786_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31972_ (.A(_15787_),
    .B(net486),
    .CO(_15788_),
    .S(_15789_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31973_ (.A(_15787_),
    .B(net41),
    .CO(_15790_),
    .S(_15791_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31974_ (.A(_15787_),
    .B(net41),
    .CO(_15792_),
    .S(_15793_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31975_ (.A(_15794_),
    .B(_15770_),
    .CO(_15795_),
    .S(_15796_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31976_ (.A(_15794_),
    .B(net4),
    .CO(_15797_),
    .S(_15798_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31977_ (.A(_15794_),
    .B(net41),
    .CO(_15799_),
    .S(_15800_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31978_ (.A(_15801_),
    .B(_15802_),
    .CO(_15803_),
    .S(_15804_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31979_ (.A(_15801_),
    .B(_15802_),
    .CO(_15805_),
    .S(_15806_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31980_ (.A(net676),
    .B(_15801_),
    .CO(_15808_),
    .S(_15809_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31981_ (.A(net664),
    .B(_15802_),
    .CO(_15811_),
    .S(_15812_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31982_ (.A(_15810_),
    .B(_15802_),
    .CO(_15813_),
    .S(_15814_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31983_ (.A(_15810_),
    .B(net677),
    .CO(_15815_),
    .S(_15816_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31984_ (.A(_15810_),
    .B(net676),
    .CO(_15817_),
    .S(_15818_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31985_ (.A(_15819_),
    .B(net547),
    .CO(_15820_),
    .S(_15821_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31986_ (.A(_15819_),
    .B(net28),
    .CO(_15822_),
    .S(_15823_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31987_ (.A(_15819_),
    .B(net658),
    .CO(_15824_),
    .S(_15825_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31988_ (.A(_15826_),
    .B(net19),
    .CO(_15827_),
    .S(_15828_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31989_ (.A(_15826_),
    .B(net547),
    .CO(_15829_),
    .S(_15830_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31990_ (.A(_15826_),
    .B(net28),
    .CO(_15831_),
    .S(_15832_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31991_ (.A(_15833_),
    .B(_15834_),
    .CO(_15835_),
    .S(_15836_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31992_ (.A(net1273),
    .B(net504),
    .CO(_15837_),
    .S(_15838_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31993_ (.A(_15833_),
    .B(_15839_),
    .CO(_15840_),
    .S(_15841_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31994_ (.A(_15842_),
    .B(net505),
    .CO(_15843_),
    .S(_15844_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31995_ (.A(_15842_),
    .B(net504),
    .CO(_15845_),
    .S(_15846_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31996_ (.A(_15842_),
    .B(_15839_),
    .CO(_15847_),
    .S(_15848_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31997_ (.A(_15842_),
    .B(net552),
    .CO(_15849_),
    .S(_15850_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31998_ (.A(_15851_),
    .B(net2),
    .CO(_15852_),
    .S(_15853_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _31999_ (.A(_15851_),
    .B(net553),
    .CO(_15854_),
    .S(_15855_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32000_ (.A(_15851_),
    .B(net554),
    .CO(_15856_),
    .S(_15857_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32001_ (.A(_15858_),
    .B(net506),
    .CO(_15859_),
    .S(_15860_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32002_ (.A(_15858_),
    .B(net505),
    .CO(_15861_),
    .S(_15862_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32003_ (.A(_15858_),
    .B(net14),
    .CO(_15863_),
    .S(_15864_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32004_ (.A(_15866_),
    .B(net1258),
    .CO(_15867_),
    .S(_15868_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32005_ (.A(net1050),
    .B(net545),
    .CO(_15869_),
    .S(_15870_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32006_ (.A(_15865_),
    .B(_15871_),
    .CO(_15872_),
    .S(_15873_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32007_ (.A(_15874_),
    .B(net543),
    .CO(_15875_),
    .S(_15876_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32008_ (.A(_15874_),
    .B(_15866_),
    .CO(_15877_),
    .S(_15878_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32009_ (.A(net1217),
    .B(_15871_),
    .CO(_15879_),
    .S(_15880_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32010_ (.A(_15874_),
    .B(_15871_),
    .CO(_15881_),
    .S(_15882_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32011_ (.A(_15883_),
    .B(net544),
    .CO(_15884_),
    .S(_15885_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32012_ (.A(_15883_),
    .B(net8),
    .CO(_15886_),
    .S(_15887_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32013_ (.A(_15883_),
    .B(net836),
    .CO(_15888_),
    .S(_15889_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32014_ (.A(_15890_),
    .B(net10),
    .CO(_15891_),
    .S(_15892_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32015_ (.A(_15890_),
    .B(net545),
    .CO(_15893_),
    .S(_15894_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32016_ (.A(_15890_),
    .B(net8),
    .CO(_15895_),
    .S(_15896_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32017_ (.A(_15897_),
    .B(_15898_),
    .CO(_15899_),
    .S(_15900_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32018_ (.A(net483),
    .B(net1088),
    .CO(_15901_),
    .S(_15902_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32019_ (.A(net500),
    .B(net483),
    .CO(_15904_),
    .S(_15905_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32020_ (.A(_15906_),
    .B(net1088),
    .CO(_15907_),
    .S(_15908_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32021_ (.A(_15906_),
    .B(net1088),
    .CO(_15909_),
    .S(_15910_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32022_ (.A(_15906_),
    .B(net16),
    .CO(_15911_),
    .S(_15912_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32023_ (.A(_15906_),
    .B(net500),
    .CO(_15913_),
    .S(_15914_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32024_ (.A(_15915_),
    .B(net21),
    .CO(_15916_),
    .S(_15917_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32025_ (.A(net501),
    .B(_15915_),
    .CO(_15918_),
    .S(_15919_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32026_ (.A(_15915_),
    .B(net16),
    .CO(_15920_),
    .S(_15921_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32027_ (.A(_15922_),
    .B(net21),
    .CO(_15923_),
    .S(_15924_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32028_ (.A(_15922_),
    .B(net1089),
    .CO(_15925_),
    .S(_15926_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32029_ (.A(_15922_),
    .B(net16),
    .CO(_15927_),
    .S(_15928_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32030_ (.A(_15929_),
    .B(_15930_),
    .CO(_15931_),
    .S(_15932_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32031_ (.A(_15929_),
    .B(net1118),
    .CO(_15933_),
    .S(_15934_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32032_ (.A(net1116),
    .B(net557),
    .CO(_15936_),
    .S(_15937_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32033_ (.A(net494),
    .B(_15935_),
    .CO(_15938_),
    .S(_15939_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32034_ (.A(_15940_),
    .B(_15930_),
    .CO(_15941_),
    .S(_15942_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32035_ (.A(_15940_),
    .B(net1118),
    .CO(_15943_),
    .S(_15944_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32036_ (.A(_15940_),
    .B(_15935_),
    .CO(_15945_),
    .S(_15946_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32037_ (.A(_15940_),
    .B(_15935_),
    .CO(_15947_),
    .S(_15948_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32038_ (.A(_15949_),
    .B(net1118),
    .CO(_15950_),
    .S(_15951_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32039_ (.A(_15949_),
    .B(net479),
    .CO(_15952_),
    .S(_15953_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32040_ (.A(_15949_),
    .B(net588),
    .CO(_15954_),
    .S(_15955_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32041_ (.A(_15956_),
    .B(net27),
    .CO(_15957_),
    .S(_15958_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32042_ (.A(_15956_),
    .B(net27),
    .CO(_15959_),
    .S(_15960_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32043_ (.A(_15956_),
    .B(net479),
    .CO(_15961_),
    .S(_15962_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32044_ (.A(_15956_),
    .B(net588),
    .CO(_15963_),
    .S(_15964_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32045_ (.A(_15966_),
    .B(_15965_),
    .CO(_15967_),
    .S(_15968_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32046_ (.A(_15965_),
    .B(_15966_),
    .CO(_15969_),
    .S(_15970_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32047_ (.A(_15965_),
    .B(_15971_),
    .CO(_15972_),
    .S(_15973_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32048_ (.A(_15965_),
    .B(_15971_),
    .CO(_15974_),
    .S(_15975_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32049_ (.A(_15976_),
    .B(_15966_),
    .CO(_15977_),
    .S(_15978_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32050_ (.A(_15976_),
    .B(_15966_),
    .CO(_15979_),
    .S(_15980_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32051_ (.A(_15976_),
    .B(_15971_),
    .CO(_15981_),
    .S(_15982_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32052_ (.A(_15976_),
    .B(_15971_),
    .CO(_15983_),
    .S(_15984_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32053_ (.A(_15985_),
    .B(net797),
    .CO(_15986_),
    .S(_15987_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32054_ (.A(_15985_),
    .B(net92),
    .CO(_15988_),
    .S(_15989_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32055_ (.A(_15985_),
    .B(_15971_),
    .CO(_15990_),
    .S(_15991_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32056_ (.A(_15992_),
    .B(net31),
    .CO(_15993_),
    .S(_15994_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32057_ (.A(_15992_),
    .B(net31),
    .CO(_15995_),
    .S(_15996_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32058_ (.A(_15992_),
    .B(net92),
    .CO(_15997_),
    .S(_15998_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32059_ (.A(_15992_),
    .B(net92),
    .CO(_15999_),
    .S(_16000_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32060_ (.A(_16002_),
    .B(_16001_),
    .CO(_16003_),
    .S(_16004_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32061_ (.A(_16001_),
    .B(net884),
    .CO(_16005_),
    .S(_16006_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32062_ (.A(_16001_),
    .B(_16007_),
    .CO(_16008_),
    .S(_16009_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32063_ (.A(_16007_),
    .B(_16001_),
    .CO(_16010_),
    .S(_16011_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32064_ (.A(_16012_),
    .B(net636),
    .CO(_16013_),
    .S(_16014_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32065_ (.A(net632),
    .B(_16002_),
    .CO(_16015_),
    .S(_16016_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32066_ (.A(net632),
    .B(_16007_),
    .CO(_16017_),
    .S(_16018_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32067_ (.A(_16012_),
    .B(_16007_),
    .CO(_16019_),
    .S(_16020_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32068_ (.A(_16021_),
    .B(net636),
    .CO(_16022_),
    .S(_16023_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32069_ (.A(_16021_),
    .B(_16007_),
    .CO(_16024_),
    .S(_16025_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32070_ (.A(_16021_),
    .B(_16007_),
    .CO(_16026_),
    .S(_16027_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32071_ (.A(_16028_),
    .B(net15),
    .CO(_16029_),
    .S(_16030_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32072_ (.A(_16028_),
    .B(net15),
    .CO(_16031_),
    .S(_16032_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32073_ (.A(_16028_),
    .B(net48),
    .CO(_16033_),
    .S(_16034_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32074_ (.A(_16028_),
    .B(net48),
    .CO(_16035_),
    .S(_16036_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32075_ (.A(_16037_),
    .B(_16038_),
    .CO(_16039_),
    .S(_16040_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32076_ (.A(net713),
    .B(net740),
    .CO(_16041_),
    .S(_16042_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32077_ (.A(net719),
    .B(_16043_),
    .CO(_16044_),
    .S(_16045_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32078_ (.A(net713),
    .B(_16043_),
    .CO(_16046_),
    .S(_16047_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32079_ (.A(_16048_),
    .B(_16038_),
    .CO(_16049_),
    .S(_16050_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32080_ (.A(_16048_),
    .B(_16038_),
    .CO(_16051_),
    .S(_16052_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32081_ (.A(_16048_),
    .B(_16043_),
    .CO(_16053_),
    .S(_16054_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32082_ (.A(_16048_),
    .B(_16043_),
    .CO(_16055_),
    .S(_16056_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32083_ (.A(_16057_),
    .B(net741),
    .CO(_16058_),
    .S(_16059_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32084_ (.A(_16057_),
    .B(net60),
    .CO(_16060_),
    .S(_16061_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32085_ (.A(_16057_),
    .B(_16043_),
    .CO(_16062_),
    .S(_16063_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32086_ (.A(_16064_),
    .B(net9),
    .CO(_16065_),
    .S(_16066_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32087_ (.A(_16064_),
    .B(net740),
    .CO(_16067_),
    .S(_16068_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32088_ (.A(_16064_),
    .B(net60),
    .CO(_16069_),
    .S(_16070_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32089_ (.A(_16064_),
    .B(net60),
    .CO(_16071_),
    .S(_16072_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32090_ (.A(_16074_),
    .B(_16073_),
    .CO(_16075_),
    .S(_16076_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32091_ (.A(net1065),
    .B(net1068),
    .CO(_16077_),
    .S(_16078_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32092_ (.A(net1065),
    .B(net1143),
    .CO(_16080_),
    .S(_16081_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32093_ (.A(_16082_),
    .B(net1068),
    .CO(_16083_),
    .S(_16084_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32094_ (.A(_16082_),
    .B(_16074_),
    .CO(_16085_),
    .S(_16086_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32095_ (.A(_16082_),
    .B(net22),
    .CO(_16087_),
    .S(_16088_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32096_ (.A(_16082_),
    .B(_16079_),
    .CO(_16089_),
    .S(_16090_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32097_ (.A(_16091_),
    .B(net73),
    .CO(_16092_),
    .S(_16093_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32098_ (.A(_16091_),
    .B(net22),
    .CO(_16094_),
    .S(_16095_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32099_ (.A(_16091_),
    .B(net22),
    .CO(_16096_),
    .S(_16097_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32100_ (.A(_16098_),
    .B(net73),
    .CO(_16099_),
    .S(_16100_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32101_ (.A(_16098_),
    .B(net73),
    .CO(_16101_),
    .S(_16102_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32102_ (.A(_16098_),
    .B(net22),
    .CO(_16103_),
    .S(_16104_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32103_ (.A(_16105_),
    .B(_16106_),
    .CO(_16107_),
    .S(_16108_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32104_ (.A(_16105_),
    .B(_16106_),
    .CO(_16109_),
    .S(_16110_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32105_ (.A(net1121),
    .B(_16111_),
    .CO(_16112_),
    .S(_16113_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32106_ (.A(_16114_),
    .B(_16106_),
    .CO(_16115_),
    .S(_16116_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32107_ (.A(_16114_),
    .B(_16106_),
    .CO(_16117_),
    .S(_16118_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32108_ (.A(_16114_),
    .B(_16111_),
    .CO(_16119_),
    .S(_16120_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32109_ (.A(_16114_),
    .B(_16111_),
    .CO(_16121_),
    .S(_16122_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32110_ (.A(_16123_),
    .B(_16106_),
    .CO(_16124_),
    .S(_16125_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32111_ (.A(_16123_),
    .B(_16111_),
    .CO(_16126_),
    .S(_16127_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32112_ (.A(_16123_),
    .B(_16111_),
    .CO(_16128_),
    .S(_16129_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32113_ (.A(_16130_),
    .B(net7),
    .CO(_16131_),
    .S(_16132_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32114_ (.A(_16130_),
    .B(_16106_),
    .CO(_16133_),
    .S(_16134_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32115_ (.A(_16130_),
    .B(net3),
    .CO(_16135_),
    .S(_16136_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32116_ (.A(_16137_),
    .B(_16138_),
    .CO(_16139_),
    .S(_16140_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32117_ (.A(_16137_),
    .B(_16138_),
    .CO(_16141_),
    .S(_16142_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32118_ (.A(net1188),
    .B(_16143_),
    .CO(_16144_),
    .S(_16145_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32119_ (.A(net1189),
    .B(net1210),
    .CO(_16147_),
    .S(_16148_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32120_ (.A(_16146_),
    .B(_16138_),
    .CO(_16149_),
    .S(_16150_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32121_ (.A(net1189),
    .B(_16143_),
    .CO(_16151_),
    .S(_16152_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32122_ (.A(net1189),
    .B(_16143_),
    .CO(_16153_),
    .S(_16154_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32123_ (.A(_16155_),
    .B(net24),
    .CO(_16156_),
    .S(_16157_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32124_ (.A(_16155_),
    .B(_16143_),
    .CO(_16158_),
    .S(_16159_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32125_ (.A(_16155_),
    .B(net1202),
    .CO(_16160_),
    .S(_16161_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32126_ (.A(_16162_),
    .B(_16138_),
    .CO(_16163_),
    .S(_16164_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32127_ (.A(_16162_),
    .B(net24),
    .CO(_16165_),
    .S(_16166_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32128_ (.A(_16162_),
    .B(net58),
    .CO(_16167_),
    .S(_16168_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32129_ (.A(_16170_),
    .B(_16169_),
    .CO(_16171_),
    .S(_16172_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32130_ (.A(_16169_),
    .B(_16170_),
    .CO(_16173_),
    .S(_16174_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32131_ (.A(_16169_),
    .B(_16175_),
    .CO(_16176_),
    .S(_16177_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32132_ (.A(_16178_),
    .B(_16170_),
    .CO(_16179_),
    .S(_16180_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32133_ (.A(_16178_),
    .B(_16170_),
    .CO(_16181_),
    .S(_16182_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32134_ (.A(_16178_),
    .B(_16175_),
    .CO(_16183_),
    .S(_16184_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32135_ (.A(_16178_),
    .B(_16175_),
    .CO(_16185_),
    .S(_16186_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32136_ (.A(_16187_),
    .B(_16170_),
    .CO(_16188_),
    .S(_16189_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32137_ (.A(_16187_),
    .B(net892),
    .CO(_16190_),
    .S(_16191_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32138_ (.A(_16187_),
    .B(_16175_),
    .CO(_16192_),
    .S(_16193_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32139_ (.A(_16194_),
    .B(net18),
    .CO(_16195_),
    .S(_16196_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32140_ (.A(_16194_),
    .B(net18),
    .CO(_16197_),
    .S(_16198_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32141_ (.A(_16194_),
    .B(net81),
    .CO(_16199_),
    .S(_16200_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32142_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_16201_),
    .CO(_16202_),
    .S(\u0.r0.rcnt_next[1] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32143_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_16203_),
    .S(_16204_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32144_ (.A(\u0.r0.rcnt[0] ),
    .B(_16201_),
    .CO(_16205_),
    .S(_16206_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32145_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_16207_),
    .S(_16208_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _32146_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_16209_),
    .S(_16210_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[0]$_SDFFE_PN0P_  (.D(_00405_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dcnt[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[1]$_SDFFE_PN0P_  (.D(_00406_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dcnt[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[2]$_SDFFE_PP0P_  (.D(_00407_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dcnt[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[3]$_SDFFE_PN0P_  (.D(_00408_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dcnt[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \done$_DFF_P_  (.D(_00160_),
    .CLK(clknet_leaf_8_clk),
    .Q(net346));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \ld_r$_DFF_P_  (.D(net953),
    .CLK(clknet_leaf_23_clk),
    .Q(ld_r));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[0]$_DFF_P_  (.D(_00032_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa00_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[1]$_DFF_P_  (.D(_00033_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa00_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[2]$_DFF_P_  (.D(_00034_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa00_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[3]$_DFF_P_  (.D(_00035_),
    .CLK(clknet_leaf_8_clk),
    .Q(\sa00_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[4]$_DFF_P_  (.D(_00036_),
    .CLK(clknet_leaf_8_clk),
    .Q(\sa00_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[5]$_DFF_P_  (.D(_00037_),
    .CLK(clknet_leaf_8_clk),
    .Q(\sa00_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[6]$_DFF_P_  (.D(_00038_),
    .CLK(clknet_leaf_8_clk),
    .Q(\sa00_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[7]$_DFF_P_  (.D(_00039_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa00_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[0]$_DFF_P_  (.D(_00040_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa01_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[1]$_DFF_P_  (.D(_00041_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa01_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[2]$_DFF_P_  (.D(_00042_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa01_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[3]$_DFF_P_  (.D(_00043_),
    .CLK(clknet_leaf_9_clk),
    .Q(\sa01_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[4]$_DFF_P_  (.D(_00044_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa01_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[5]$_DFF_P_  (.D(_00045_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa01_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[6]$_DFF_P_  (.D(_00046_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa01_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[7]$_DFF_P_  (.D(_00047_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa01_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[0]$_DFF_P_  (.D(_00048_),
    .CLK(clknet_leaf_15_clk),
    .Q(\sa02_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[1]$_DFF_P_  (.D(_00049_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa02_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[2]$_DFF_P_  (.D(_00050_),
    .CLK(clknet_leaf_14_clk),
    .Q(\sa02_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[3]$_DFF_P_  (.D(_00051_),
    .CLK(clknet_leaf_14_clk),
    .Q(\sa02_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[4]$_DFF_P_  (.D(_00052_),
    .CLK(clknet_leaf_15_clk),
    .Q(\sa02_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[5]$_DFF_P_  (.D(_00053_),
    .CLK(clknet_leaf_15_clk),
    .Q(\sa02_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[6]$_DFF_P_  (.D(_00054_),
    .CLK(clknet_leaf_15_clk),
    .Q(\sa02_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[7]$_DFF_P_  (.D(_00055_),
    .CLK(clknet_leaf_14_clk),
    .Q(\sa02_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[0]$_DFF_P_  (.D(_00056_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa03_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[1]$_DFF_P_  (.D(_00057_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa03_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[2]$_DFF_P_  (.D(_00058_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa03_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[3]$_DFF_P_  (.D(_00059_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa03_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[4]$_DFF_P_  (.D(_00060_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa03_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[5]$_DFF_P_  (.D(_00061_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa03_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[6]$_DFF_P_  (.D(_00062_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa03_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[7]$_DFF_P_  (.D(_00063_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa03_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[0]$_DFF_P_  (.D(_00072_),
    .CLK(clknet_leaf_8_clk),
    .Q(\sa10_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[1]$_DFF_P_  (.D(_00073_),
    .CLK(clknet_leaf_7_clk),
    .Q(\sa10_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[2]$_DFF_P_  (.D(_00074_),
    .CLK(clknet_leaf_7_clk),
    .Q(\sa10_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[3]$_DFF_P_  (.D(_00075_),
    .CLK(clknet_leaf_8_clk),
    .Q(\sa10_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[4]$_DFF_P_  (.D(_00076_),
    .CLK(clknet_leaf_7_clk),
    .Q(\sa10_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[5]$_DFF_P_  (.D(_00077_),
    .CLK(clknet_leaf_7_clk),
    .Q(\sa10_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[6]$_DFF_P_  (.D(_00078_),
    .CLK(clknet_leaf_7_clk),
    .Q(\sa10_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[7]$_DFF_P_  (.D(_00079_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa10_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[0]$_DFF_P_  (.D(_00080_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa11_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[1]$_DFF_P_  (.D(_00081_),
    .CLK(clknet_leaf_12_clk),
    .Q(\sa11_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[2]$_DFF_P_  (.D(_00082_),
    .CLK(clknet_leaf_12_clk),
    .Q(\sa11_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[3]$_DFF_P_  (.D(_00083_),
    .CLK(clknet_leaf_12_clk),
    .Q(\sa11_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[4]$_DFF_P_  (.D(_00084_),
    .CLK(clknet_leaf_12_clk),
    .Q(\sa11_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[5]$_DFF_P_  (.D(_00085_),
    .CLK(clknet_leaf_12_clk),
    .Q(\sa11_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[6]$_DFF_P_  (.D(_00086_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa11_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[7]$_DFF_P_  (.D(_00087_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa11_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[0]$_DFF_P_  (.D(_00088_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[1]$_DFF_P_  (.D(_00089_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[2]$_DFF_P_  (.D(_00090_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[3]$_DFF_P_  (.D(_00091_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[4]$_DFF_P_  (.D(_00092_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[5]$_DFF_P_  (.D(_00093_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[6]$_DFF_P_  (.D(_00094_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[7]$_DFF_P_  (.D(_00095_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa12_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[0]$_DFF_P_  (.D(_00064_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa10_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[1]$_DFF_P_  (.D(_00065_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa10_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[2]$_DFF_P_  (.D(_00066_),
    .CLK(clknet_leaf_23_clk),
    .Q(\sa10_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[3]$_DFF_P_  (.D(_00067_),
    .CLK(clknet_leaf_23_clk),
    .Q(\sa10_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[4]$_DFF_P_  (.D(_00068_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa10_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[5]$_DFF_P_  (.D(_00069_),
    .CLK(clknet_leaf_3_clk),
    .Q(\sa10_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[6]$_DFF_P_  (.D(_00070_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa10_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[7]$_DFF_P_  (.D(_00071_),
    .CLK(clknet_leaf_23_clk),
    .Q(\sa10_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[0]$_DFF_P_  (.D(_00112_),
    .CLK(clknet_leaf_11_clk),
    .Q(\sa20_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[1]$_DFF_P_  (.D(_00113_),
    .CLK(clknet_leaf_11_clk),
    .Q(\sa20_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[2]$_DFF_P_  (.D(_00114_),
    .CLK(clknet_leaf_5_clk),
    .Q(\sa20_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[3]$_DFF_P_  (.D(_00115_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa20_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[4]$_DFF_P_  (.D(_00116_),
    .CLK(clknet_leaf_4_clk),
    .Q(\sa20_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[5]$_DFF_P_  (.D(_00117_),
    .CLK(clknet_leaf_4_clk),
    .Q(\sa20_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[6]$_DFF_P_  (.D(_00118_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa20_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[7]$_DFF_P_  (.D(_00119_),
    .CLK(clknet_leaf_4_clk),
    .Q(\sa20_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[0]$_DFF_P_  (.D(_00120_),
    .CLK(clknet_leaf_24_clk),
    .Q(\sa21_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[1]$_DFF_P_  (.D(_00121_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[2]$_DFF_P_  (.D(_00122_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[3]$_DFF_P_  (.D(_00123_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[4]$_DFF_P_  (.D(_00124_),
    .CLK(clknet_leaf_23_clk),
    .Q(\sa21_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[5]$_DFF_P_  (.D(_00125_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[6]$_DFF_P_  (.D(_00126_),
    .CLK(clknet_leaf_24_clk),
    .Q(\sa21_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[7]$_DFF_P_  (.D(_00127_),
    .CLK(clknet_leaf_3_clk),
    .Q(\sa21_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[0]$_DFF_P_  (.D(_00096_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa20_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[1]$_DFF_P_  (.D(_00097_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa20_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[2]$_DFF_P_  (.D(_00098_),
    .CLK(clknet_leaf_11_clk),
    .Q(\sa20_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[3]$_DFF_P_  (.D(_00099_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa20_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[4]$_DFF_P_  (.D(_00100_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa20_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[5]$_DFF_P_  (.D(_00101_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa20_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[6]$_DFF_P_  (.D(_00102_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa20_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[7]$_DFF_P_  (.D(_00103_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa20_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[0]$_DFF_P_  (.D(_00104_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[1]$_DFF_P_  (.D(_00105_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[2]$_DFF_P_  (.D(_00106_),
    .CLK(clknet_leaf_26_clk),
    .Q(\sa21_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[3]$_DFF_P_  (.D(_00107_),
    .CLK(clknet_leaf_26_clk),
    .Q(\sa21_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[4]$_DFF_P_  (.D(_00108_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa21_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[5]$_DFF_P_  (.D(_00109_),
    .CLK(clknet_leaf_25_clk),
    .Q(\sa21_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[6]$_DFF_P_  (.D(_00110_),
    .CLK(clknet_leaf_26_clk),
    .Q(\sa21_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[7]$_DFF_P_  (.D(_00111_),
    .CLK(clknet_leaf_22_clk),
    .Q(\sa21_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[0]$_DFF_P_  (.D(_00152_),
    .CLK(clknet_leaf_11_clk),
    .Q(\sa30_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[1]$_DFF_P_  (.D(_00153_),
    .CLK(clknet_leaf_11_clk),
    .Q(\sa30_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[2]$_DFF_P_  (.D(_00154_),
    .CLK(clknet_leaf_11_clk),
    .Q(\sa30_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[3]$_DFF_P_  (.D(_00155_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa30_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[4]$_DFF_P_  (.D(_00156_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa30_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[5]$_DFF_P_  (.D(_00157_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa30_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[6]$_DFF_P_  (.D(_00158_),
    .CLK(clknet_leaf_17_clk),
    .Q(\sa30_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[7]$_DFF_P_  (.D(_00159_),
    .CLK(clknet_leaf_4_clk),
    .Q(\sa30_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[0]$_DFF_P_  (.D(_00128_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[1]$_DFF_P_  (.D(_00129_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[2]$_DFF_P_  (.D(_00130_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[3]$_DFF_P_  (.D(_00131_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[4]$_DFF_P_  (.D(_00132_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[5]$_DFF_P_  (.D(_00133_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[6]$_DFF_P_  (.D(_00134_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[7]$_DFF_P_  (.D(_00135_),
    .CLK(clknet_leaf_10_clk),
    .Q(\sa30_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[0]$_DFF_P_  (.D(_00136_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[1]$_DFF_P_  (.D(_00137_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[2]$_DFF_P_  (.D(_00138_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[3]$_DFF_P_  (.D(_00139_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[4]$_DFF_P_  (.D(_00140_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[5]$_DFF_P_  (.D(_00141_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[6]$_DFF_P_  (.D(_00142_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[7]$_DFF_P_  (.D(_00143_),
    .CLK(clknet_leaf_16_clk),
    .Q(\sa31_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[0]$_DFF_P_  (.D(_00144_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[1]$_DFF_P_  (.D(_00145_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[2]$_DFF_P_  (.D(_00146_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[3]$_DFF_P_  (.D(_00147_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[4]$_DFF_P_  (.D(_00148_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[5]$_DFF_P_  (.D(_00149_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[6]$_DFF_P_  (.D(_00150_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[7]$_DFF_P_  (.D(_00151_),
    .CLK(clknet_leaf_18_clk),
    .Q(\sa32_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[0]$_DFFE_PP_  (.D(_00409_),
    .CLK(clknet_leaf_24_clk),
    .Q(\text_in_r[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[100]$_DFFE_PP_  (.D(_00410_),
    .CLK(clknet_leaf_4_clk),
    .Q(\text_in_r[100] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[101]$_DFFE_PP_  (.D(_00411_),
    .CLK(clknet_leaf_4_clk),
    .Q(\text_in_r[101] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[102]$_DFFE_PP_  (.D(_00412_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[102] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[103]$_DFFE_PP_  (.D(_00413_),
    .CLK(clknet_leaf_4_clk),
    .Q(\text_in_r[103] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[104]$_DFFE_PP_  (.D(_00414_),
    .CLK(clknet_leaf_10_clk),
    .Q(\text_in_r[104] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[105]$_DFFE_PP_  (.D(_00415_),
    .CLK(clknet_leaf_10_clk),
    .Q(\text_in_r[105] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[106]$_DFFE_PP_  (.D(_00416_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[106] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[107]$_DFFE_PP_  (.D(_00417_),
    .CLK(clknet_leaf_10_clk),
    .Q(\text_in_r[107] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[108]$_DFFE_PP_  (.D(_00418_),
    .CLK(clknet_leaf_10_clk),
    .Q(\text_in_r[108] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[109]$_DFFE_PP_  (.D(_00419_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[109] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[10]$_DFFE_PP_  (.D(_00420_),
    .CLK(clknet_leaf_23_clk),
    .Q(\text_in_r[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[110]$_DFFE_PP_  (.D(_00421_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[110] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[111]$_DFFE_PP_  (.D(_00422_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[111] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[112]$_DFFE_PP_  (.D(_00423_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[112] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[113]$_DFFE_PP_  (.D(_00424_),
    .CLK(clknet_leaf_25_clk),
    .Q(\text_in_r[113] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[114]$_DFFE_PP_  (.D(_00425_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[114] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[115]$_DFFE_PP_  (.D(_00426_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[115] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[116]$_DFFE_PP_  (.D(_00427_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[116] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[117]$_DFFE_PP_  (.D(_00428_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[117] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[118]$_DFFE_PP_  (.D(_00429_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[118] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[119]$_DFFE_PP_  (.D(_00430_),
    .CLK(clknet_leaf_0_clk),
    .Q(\text_in_r[119] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[11]$_DFFE_PP_  (.D(_00431_),
    .CLK(clknet_leaf_17_clk),
    .Q(\text_in_r[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[120]$_DFFE_PP_  (.D(_00432_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[120] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[121]$_DFFE_PP_  (.D(_00433_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[121] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[122]$_DFFE_PP_  (.D(_00434_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[122] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[123]$_DFFE_PP_  (.D(_00435_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[123] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[124]$_DFFE_PP_  (.D(_00436_),
    .CLK(clknet_leaf_7_clk),
    .Q(\text_in_r[124] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[125]$_DFFE_PP_  (.D(_00437_),
    .CLK(clknet_leaf_7_clk),
    .Q(\text_in_r[125] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[126]$_DFFE_PP_  (.D(_00438_),
    .CLK(clknet_leaf_7_clk),
    .Q(\text_in_r[126] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[127]$_DFFE_PP_  (.D(_00439_),
    .CLK(clknet_leaf_7_clk),
    .Q(\text_in_r[127] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[12]$_DFFE_PP_  (.D(_00440_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[13]$_DFFE_PP_  (.D(_00441_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[14]$_DFFE_PP_  (.D(_00442_),
    .CLK(clknet_leaf_23_clk),
    .Q(\text_in_r[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[15]$_DFFE_PP_  (.D(_00443_),
    .CLK(clknet_leaf_23_clk),
    .Q(\text_in_r[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[16]$_DFFE_PP_  (.D(_00444_),
    .CLK(clknet_leaf_20_clk),
    .Q(\text_in_r[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[17]$_DFFE_PP_  (.D(_00445_),
    .CLK(clknet_leaf_20_clk),
    .Q(\text_in_r[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[18]$_DFFE_PP_  (.D(_00446_),
    .CLK(clknet_leaf_20_clk),
    .Q(\text_in_r[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[19]$_DFFE_PP_  (.D(_00447_),
    .CLK(clknet_leaf_20_clk),
    .Q(\text_in_r[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[1]$_DFFE_PP_  (.D(_00448_),
    .CLK(clknet_leaf_18_clk),
    .Q(\text_in_r[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[20]$_DFFE_PP_  (.D(_00449_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[21]$_DFFE_PP_  (.D(_00450_),
    .CLK(clknet_leaf_18_clk),
    .Q(\text_in_r[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[22]$_DFFE_PP_  (.D(_00451_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[23]$_DFFE_PP_  (.D(_00452_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[24]$_DFFE_PP_  (.D(_00453_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[25]$_DFFE_PP_  (.D(_00454_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[26]$_DFFE_PP_  (.D(_00455_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[27]$_DFFE_PP_  (.D(_00456_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[28]$_DFFE_PP_  (.D(_00457_),
    .CLK(clknet_leaf_18_clk),
    .Q(\text_in_r[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[29]$_DFFE_PP_  (.D(_00458_),
    .CLK(clknet_leaf_18_clk),
    .Q(\text_in_r[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[2]$_DFFE_PP_  (.D(_00459_),
    .CLK(clknet_leaf_22_clk),
    .Q(\text_in_r[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[30]$_DFFE_PP_  (.D(_00460_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[31]$_DFFE_PP_  (.D(_00461_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[32]$_DFFE_PP_  (.D(_00462_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[33]$_DFFE_PP_  (.D(_00463_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[34]$_DFFE_PP_  (.D(_00464_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[35]$_DFFE_PP_  (.D(_00465_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[36]$_DFFE_PP_  (.D(_00466_),
    .CLK(clknet_leaf_16_clk),
    .Q(\text_in_r[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[37]$_DFFE_PP_  (.D(_00467_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[38]$_DFFE_PP_  (.D(_00468_),
    .CLK(clknet_leaf_16_clk),
    .Q(\text_in_r[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[39]$_DFFE_PP_  (.D(_00469_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[3]$_DFFE_PP_  (.D(_00470_),
    .CLK(clknet_leaf_20_clk),
    .Q(\text_in_r[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[40]$_DFFE_PP_  (.D(_00471_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[41]$_DFFE_PP_  (.D(_00472_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[42]$_DFFE_PP_  (.D(_00473_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[43]$_DFFE_PP_  (.D(_00474_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[44]$_DFFE_PP_  (.D(_00475_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[45]$_DFFE_PP_  (.D(_00476_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[46]$_DFFE_PP_  (.D(_00477_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[47]$_DFFE_PP_  (.D(_00478_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[48]$_DFFE_PP_  (.D(_00479_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[49]$_DFFE_PP_  (.D(_00480_),
    .CLK(clknet_leaf_16_clk),
    .Q(\text_in_r[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[4]$_DFFE_PP_  (.D(_00481_),
    .CLK(clknet_leaf_17_clk),
    .Q(\text_in_r[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[50]$_DFFE_PP_  (.D(_00482_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[51]$_DFFE_PP_  (.D(_00483_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[52]$_DFFE_PP_  (.D(_00484_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[53]$_DFFE_PP_  (.D(_00485_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[54]$_DFFE_PP_  (.D(_00486_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[55]$_DFFE_PP_  (.D(_00487_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[56]$_DFFE_PP_  (.D(_00488_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[57]$_DFFE_PP_  (.D(_00489_),
    .CLK(clknet_leaf_14_clk),
    .Q(\text_in_r[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[58]$_DFFE_PP_  (.D(_00490_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[59]$_DFFE_PP_  (.D(_00491_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[5]$_DFFE_PP_  (.D(_00492_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[60]$_DFFE_PP_  (.D(_00493_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[61]$_DFFE_PP_  (.D(_00494_),
    .CLK(clknet_leaf_12_clk),
    .Q(\text_in_r[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[62]$_DFFE_PP_  (.D(_00495_),
    .CLK(clknet_leaf_12_clk),
    .Q(\text_in_r[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[63]$_DFFE_PP_  (.D(_00496_),
    .CLK(clknet_leaf_15_clk),
    .Q(\text_in_r[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[64]$_DFFE_PP_  (.D(_00497_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[64] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[65]$_DFFE_PP_  (.D(_00498_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[65] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[66]$_DFFE_PP_  (.D(_00499_),
    .CLK(clknet_leaf_19_clk),
    .Q(\text_in_r[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[67]$_DFFE_PP_  (.D(_00500_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[68]$_DFFE_PP_  (.D(_00501_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[68] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[69]$_DFFE_PP_  (.D(_00502_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[69] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[6]$_DFFE_PP_  (.D(_00503_),
    .CLK(clknet_leaf_17_clk),
    .Q(\text_in_r[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[70]$_DFFE_PP_  (.D(_00504_),
    .CLK(clknet_leaf_11_clk),
    .Q(\text_in_r[70] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[71]$_DFFE_PP_  (.D(_00505_),
    .CLK(clknet_leaf_4_clk),
    .Q(\text_in_r[71] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[72]$_DFFE_PP_  (.D(_00506_),
    .CLK(clknet_leaf_24_clk),
    .Q(\text_in_r[72] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[73]$_DFFE_PP_  (.D(_00507_),
    .CLK(clknet_leaf_25_clk),
    .Q(\text_in_r[73] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[74]$_DFFE_PP_  (.D(_00508_),
    .CLK(clknet_leaf_24_clk),
    .Q(\text_in_r[74] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[75]$_DFFE_PP_  (.D(_00509_),
    .CLK(clknet_leaf_25_clk),
    .Q(\text_in_r[75] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[76]$_DFFE_PP_  (.D(_00510_),
    .CLK(clknet_leaf_17_clk),
    .Q(\text_in_r[76] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[77]$_DFFE_PP_  (.D(_00511_),
    .CLK(clknet_leaf_23_clk),
    .Q(\text_in_r[77] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[78]$_DFFE_PP_  (.D(_00512_),
    .CLK(clknet_leaf_4_clk),
    .Q(\text_in_r[78] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[79]$_DFFE_PP_  (.D(_00513_),
    .CLK(clknet_leaf_3_clk),
    .Q(\text_in_r[79] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[7]$_DFFE_PP_  (.D(_00514_),
    .CLK(clknet_leaf_17_clk),
    .Q(\text_in_r[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[80]$_DFFE_PP_  (.D(_00515_),
    .CLK(clknet_leaf_8_clk),
    .Q(\text_in_r[80] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[81]$_DFFE_PP_  (.D(_00516_),
    .CLK(clknet_leaf_8_clk),
    .Q(\text_in_r[81] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[82]$_DFFE_PP_  (.D(_00517_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[82] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[83]$_DFFE_PP_  (.D(_00518_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[83] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[84]$_DFFE_PP_  (.D(_00519_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[84] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[85]$_DFFE_PP_  (.D(_00520_),
    .CLK(clknet_leaf_7_clk),
    .Q(\text_in_r[85] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[86]$_DFFE_PP_  (.D(_00521_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[86] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[87]$_DFFE_PP_  (.D(_00522_),
    .CLK(clknet_leaf_7_clk),
    .Q(\text_in_r[87] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[88]$_DFFE_PP_  (.D(_00523_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[88] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[89]$_DFFE_PP_  (.D(_00524_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[89] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[8]$_DFFE_PP_  (.D(_00525_),
    .CLK(clknet_leaf_23_clk),
    .Q(\text_in_r[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[90]$_DFFE_PP_  (.D(_00526_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[90] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[91]$_DFFE_PP_  (.D(_00527_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[91] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[92]$_DFFE_PP_  (.D(_00528_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[92] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[93]$_DFFE_PP_  (.D(_00529_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[93] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[94]$_DFFE_PP_  (.D(_00530_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[94] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[95]$_DFFE_PP_  (.D(_00531_),
    .CLK(clknet_leaf_6_clk),
    .Q(\text_in_r[95] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[96]$_DFFE_PP_  (.D(_00532_),
    .CLK(clknet_leaf_12_clk),
    .Q(\text_in_r[96] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[97]$_DFFE_PP_  (.D(_00533_),
    .CLK(clknet_leaf_12_clk),
    .Q(\text_in_r[97] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[98]$_DFFE_PP_  (.D(_00534_),
    .CLK(clknet_leaf_12_clk),
    .Q(\text_in_r[98] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[99]$_DFFE_PP_  (.D(_00535_),
    .CLK(clknet_leaf_4_clk),
    .Q(\text_in_r[99] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[9]$_DFFE_PP_  (.D(_00536_),
    .CLK(clknet_leaf_23_clk),
    .Q(\text_in_r[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[0]$_DFF_P_  (.D(_00265_),
    .CLK(clknet_leaf_20_clk),
    .Q(net347));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[100]$_DFF_P_  (.D(_00165_),
    .CLK(clknet_leaf_13_clk),
    .Q(net348));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[101]$_DFF_P_  (.D(_00166_),
    .CLK(clknet_leaf_13_clk),
    .Q(net349));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[102]$_DFF_P_  (.D(_00167_),
    .CLK(clknet_leaf_13_clk),
    .Q(net350));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[103]$_DFF_P_  (.D(_00168_),
    .CLK(clknet_leaf_7_clk),
    .Q(net351));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[104]$_DFF_P_  (.D(_00169_),
    .CLK(clknet_leaf_9_clk),
    .Q(net352));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[105]$_DFF_P_  (.D(_00170_),
    .CLK(clknet_leaf_7_clk),
    .Q(net353));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[106]$_DFF_P_  (.D(_00171_),
    .CLK(clknet_leaf_4_clk),
    .Q(net354));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[107]$_DFF_P_  (.D(_00172_),
    .CLK(clknet_leaf_7_clk),
    .Q(net355));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[108]$_DFF_P_  (.D(_00173_),
    .CLK(clknet_leaf_7_clk),
    .Q(net356));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[109]$_DFF_P_  (.D(_00174_),
    .CLK(clknet_leaf_0_clk),
    .Q(net357));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[10]$_DFF_P_  (.D(_00195_),
    .CLK(clknet_leaf_22_clk),
    .Q(net358));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[110]$_DFF_P_  (.D(_00175_),
    .CLK(clknet_leaf_0_clk),
    .Q(net359));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[111]$_DFF_P_  (.D(_00176_),
    .CLK(clknet_leaf_0_clk),
    .Q(net360));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[112]$_DFF_P_  (.D(_00177_),
    .CLK(clknet_leaf_0_clk),
    .Q(net361));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[113]$_DFF_P_  (.D(_00178_),
    .CLK(clknet_leaf_0_clk),
    .Q(net362));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[114]$_DFF_P_  (.D(_00179_),
    .CLK(clknet_leaf_0_clk),
    .Q(net363));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[115]$_DFF_P_  (.D(_00180_),
    .CLK(clknet_leaf_0_clk),
    .Q(net364));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[116]$_DFF_P_  (.D(_00181_),
    .CLK(clknet_leaf_0_clk),
    .Q(net365));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[117]$_DFF_P_  (.D(_00182_),
    .CLK(clknet_leaf_0_clk),
    .Q(net366));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[118]$_DFF_P_  (.D(_00183_),
    .CLK(clknet_leaf_0_clk),
    .Q(net367));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[119]$_DFF_P_  (.D(_00184_),
    .CLK(clknet_leaf_0_clk),
    .Q(net368));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[11]$_DFF_P_  (.D(_00196_),
    .CLK(clknet_leaf_21_clk),
    .Q(net369));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[120]$_DFF_P_  (.D(_00185_),
    .CLK(clknet_leaf_6_clk),
    .Q(net370));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[121]$_DFF_P_  (.D(_00186_),
    .CLK(clknet_leaf_6_clk),
    .Q(net371));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[122]$_DFF_P_  (.D(_00187_),
    .CLK(clknet_leaf_6_clk),
    .Q(net372));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[123]$_DFF_P_  (.D(_00188_),
    .CLK(clknet_leaf_7_clk),
    .Q(net373));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[124]$_DFF_P_  (.D(_00189_),
    .CLK(clknet_leaf_7_clk),
    .Q(net374));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[125]$_DFF_P_  (.D(_00190_),
    .CLK(clknet_leaf_7_clk),
    .Q(net375));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[126]$_DFF_P_  (.D(_00191_),
    .CLK(clknet_leaf_7_clk),
    .Q(net376));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[127]$_DFF_P_  (.D(_00192_),
    .CLK(clknet_leaf_7_clk),
    .Q(net377));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[12]$_DFF_P_  (.D(_00197_),
    .CLK(clknet_leaf_21_clk),
    .Q(net378));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[13]$_DFF_P_  (.D(_00198_),
    .CLK(clknet_leaf_21_clk),
    .Q(net379));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[14]$_DFF_P_  (.D(_00199_),
    .CLK(clknet_leaf_21_clk),
    .Q(net380));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[15]$_DFF_P_  (.D(_00200_),
    .CLK(clknet_leaf_21_clk),
    .Q(net381));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[16]$_DFF_P_  (.D(_00201_),
    .CLK(clknet_leaf_21_clk),
    .Q(net382));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[17]$_DFF_P_  (.D(_00202_),
    .CLK(clknet_leaf_26_clk),
    .Q(net383));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[18]$_DFF_P_  (.D(_00203_),
    .CLK(clknet_leaf_21_clk),
    .Q(net384));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[19]$_DFF_P_  (.D(_00204_),
    .CLK(clknet_leaf_21_clk),
    .Q(net385));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[1]$_DFF_P_  (.D(_00266_),
    .CLK(clknet_leaf_20_clk),
    .Q(net386));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[20]$_DFF_P_  (.D(_00205_),
    .CLK(clknet_leaf_21_clk),
    .Q(net387));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[21]$_DFF_P_  (.D(_00206_),
    .CLK(clknet_leaf_21_clk),
    .Q(net388));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[22]$_DFF_P_  (.D(_00207_),
    .CLK(clknet_leaf_20_clk),
    .Q(net389));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[23]$_DFF_P_  (.D(_00208_),
    .CLK(clknet_leaf_20_clk),
    .Q(net390));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[24]$_DFF_P_  (.D(_00209_),
    .CLK(clknet_leaf_21_clk),
    .Q(net391));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[25]$_DFF_P_  (.D(_00210_),
    .CLK(clknet_leaf_20_clk),
    .Q(net392));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[26]$_DFF_P_  (.D(_00211_),
    .CLK(clknet_leaf_21_clk),
    .Q(net393));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[27]$_DFF_P_  (.D(_00212_),
    .CLK(clknet_leaf_21_clk),
    .Q(net394));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[28]$_DFF_P_  (.D(_00213_),
    .CLK(clknet_leaf_19_clk),
    .Q(net395));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[29]$_DFF_P_  (.D(_00214_),
    .CLK(clknet_leaf_19_clk),
    .Q(net396));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[2]$_DFF_P_  (.D(_00267_),
    .CLK(clknet_leaf_21_clk),
    .Q(net397));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[30]$_DFF_P_  (.D(_00215_),
    .CLK(clknet_leaf_19_clk),
    .Q(net398));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[31]$_DFF_P_  (.D(_00216_),
    .CLK(clknet_leaf_19_clk),
    .Q(net399));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[32]$_DFF_P_  (.D(_00217_),
    .CLK(clknet_leaf_14_clk),
    .Q(net400));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[33]$_DFF_P_  (.D(_00218_),
    .CLK(clknet_leaf_14_clk),
    .Q(net401));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[34]$_DFF_P_  (.D(_00219_),
    .CLK(clknet_leaf_14_clk),
    .Q(net402));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[35]$_DFF_P_  (.D(_00220_),
    .CLK(clknet_leaf_14_clk),
    .Q(net403));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[36]$_DFF_P_  (.D(_00221_),
    .CLK(clknet_leaf_14_clk),
    .Q(net404));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[37]$_DFF_P_  (.D(_00222_),
    .CLK(clknet_leaf_14_clk),
    .Q(net405));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[38]$_DFF_P_  (.D(_00223_),
    .CLK(clknet_leaf_13_clk),
    .Q(net406));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[39]$_DFF_P_  (.D(_00224_),
    .CLK(clknet_leaf_15_clk),
    .Q(net407));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[3]$_DFF_P_  (.D(_00268_),
    .CLK(clknet_leaf_20_clk),
    .Q(net408));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[40]$_DFF_P_  (.D(_00225_),
    .CLK(clknet_leaf_15_clk),
    .Q(net409));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[41]$_DFF_P_  (.D(_00226_),
    .CLK(clknet_leaf_19_clk),
    .Q(net410));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[42]$_DFF_P_  (.D(_00227_),
    .CLK(clknet_leaf_19_clk),
    .Q(net411));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[43]$_DFF_P_  (.D(_00228_),
    .CLK(clknet_leaf_19_clk),
    .Q(net412));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[44]$_DFF_P_  (.D(_00229_),
    .CLK(clknet_leaf_19_clk),
    .Q(net413));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[45]$_DFF_P_  (.D(_00230_),
    .CLK(clknet_leaf_19_clk),
    .Q(net414));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[46]$_DFF_P_  (.D(_00231_),
    .CLK(clknet_leaf_15_clk),
    .Q(net415));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[47]$_DFF_P_  (.D(_00232_),
    .CLK(clknet_leaf_19_clk),
    .Q(net416));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[48]$_DFF_P_  (.D(_00233_),
    .CLK(clknet_leaf_20_clk),
    .Q(net417));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[49]$_DFF_P_  (.D(_00234_),
    .CLK(clknet_leaf_19_clk),
    .Q(net418));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[4]$_DFF_P_  (.D(_00269_),
    .CLK(clknet_leaf_19_clk),
    .Q(net419));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[50]$_DFF_P_  (.D(_00235_),
    .CLK(clknet_leaf_19_clk),
    .Q(net420));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[51]$_DFF_P_  (.D(_00236_),
    .CLK(clknet_leaf_19_clk),
    .Q(net421));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[52]$_DFF_P_  (.D(_00237_),
    .CLK(clknet_leaf_19_clk),
    .Q(net422));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[53]$_DFF_P_  (.D(_00238_),
    .CLK(clknet_leaf_19_clk),
    .Q(net423));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[54]$_DFF_P_  (.D(_00239_),
    .CLK(clknet_leaf_19_clk),
    .Q(net424));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[55]$_DFF_P_  (.D(_00240_),
    .CLK(clknet_leaf_14_clk),
    .Q(net425));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[56]$_DFF_P_  (.D(_00241_),
    .CLK(clknet_leaf_14_clk),
    .Q(net426));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[57]$_DFF_P_  (.D(_00242_),
    .CLK(clknet_leaf_14_clk),
    .Q(net427));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[58]$_DFF_P_  (.D(_00243_),
    .CLK(clknet_leaf_14_clk),
    .Q(net428));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[59]$_DFF_P_  (.D(_00244_),
    .CLK(clknet_leaf_14_clk),
    .Q(net429));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[5]$_DFF_P_  (.D(_00270_),
    .CLK(clknet_leaf_19_clk),
    .Q(net430));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[60]$_DFF_P_  (.D(_00245_),
    .CLK(clknet_leaf_15_clk),
    .Q(net431));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[61]$_DFF_P_  (.D(_00246_),
    .CLK(clknet_leaf_13_clk),
    .Q(net432));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[62]$_DFF_P_  (.D(_00247_),
    .CLK(clknet_leaf_15_clk),
    .Q(net433));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[63]$_DFF_P_  (.D(_00248_),
    .CLK(clknet_leaf_15_clk),
    .Q(net434));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[64]$_DFF_P_  (.D(_00249_),
    .CLK(clknet_leaf_13_clk),
    .Q(net435));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[65]$_DFF_P_  (.D(_00250_),
    .CLK(clknet_leaf_13_clk),
    .Q(net436));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[66]$_DFF_P_  (.D(_00251_),
    .CLK(clknet_leaf_13_clk),
    .Q(net437));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[67]$_DFF_P_  (.D(_00252_),
    .CLK(clknet_leaf_13_clk),
    .Q(net438));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[68]$_DFF_P_  (.D(_00253_),
    .CLK(clknet_leaf_13_clk),
    .Q(net439));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[69]$_DFF_P_  (.D(_00254_),
    .CLK(clknet_leaf_9_clk),
    .Q(net440));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[6]$_DFF_P_  (.D(_00271_),
    .CLK(clknet_leaf_19_clk),
    .Q(net441));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[70]$_DFF_P_  (.D(_00255_),
    .CLK(clknet_leaf_9_clk),
    .Q(net442));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[71]$_DFF_P_  (.D(_00256_),
    .CLK(clknet_leaf_4_clk),
    .Q(net443));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[72]$_DFF_P_  (.D(_00257_),
    .CLK(clknet_leaf_19_clk),
    .Q(net444));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[73]$_DFF_P_  (.D(_00258_),
    .CLK(clknet_leaf_26_clk),
    .Q(net445));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[74]$_DFF_P_  (.D(_00259_),
    .CLK(clknet_leaf_0_clk),
    .Q(net446));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[75]$_DFF_P_  (.D(_00260_),
    .CLK(clknet_leaf_26_clk),
    .Q(net447));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[76]$_DFF_P_  (.D(_00261_),
    .CLK(clknet_leaf_21_clk),
    .Q(net448));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[77]$_DFF_P_  (.D(_00262_),
    .CLK(clknet_leaf_26_clk),
    .Q(net449));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[78]$_DFF_P_  (.D(_00263_),
    .CLK(clknet_leaf_26_clk),
    .Q(net450));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[79]$_DFF_P_  (.D(_00264_),
    .CLK(clknet_leaf_7_clk),
    .Q(net451));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[7]$_DFF_P_  (.D(_00272_),
    .CLK(clknet_leaf_19_clk),
    .Q(net452));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[80]$_DFF_P_  (.D(_00273_),
    .CLK(clknet_leaf_5_clk),
    .Q(net453));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[81]$_DFF_P_  (.D(_00274_),
    .CLK(clknet_leaf_8_clk),
    .Q(net454));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[82]$_DFF_P_  (.D(_00275_),
    .CLK(clknet_leaf_5_clk),
    .Q(net455));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[83]$_DFF_P_  (.D(_00276_),
    .CLK(clknet_leaf_5_clk),
    .Q(net456));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[84]$_DFF_P_  (.D(_00277_),
    .CLK(clknet_leaf_9_clk),
    .Q(net457));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[85]$_DFF_P_  (.D(_00278_),
    .CLK(clknet_leaf_8_clk),
    .Q(net458));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[86]$_DFF_P_  (.D(_00279_),
    .CLK(clknet_leaf_6_clk),
    .Q(net459));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[87]$_DFF_P_  (.D(_00280_),
    .CLK(clknet_leaf_7_clk),
    .Q(net460));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[88]$_DFF_P_  (.D(_00281_),
    .CLK(clknet_leaf_9_clk),
    .Q(net461));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[89]$_DFF_P_  (.D(_00282_),
    .CLK(clknet_leaf_9_clk),
    .Q(net462));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[8]$_DFF_P_  (.D(_00193_),
    .CLK(clknet_leaf_21_clk),
    .Q(net463));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[90]$_DFF_P_  (.D(_00283_),
    .CLK(clknet_leaf_9_clk),
    .Q(net464));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[91]$_DFF_P_  (.D(_00284_),
    .CLK(clknet_leaf_9_clk),
    .Q(net465));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[92]$_DFF_P_  (.D(_00285_),
    .CLK(clknet_leaf_6_clk),
    .Q(net466));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[93]$_DFF_P_  (.D(_00286_),
    .CLK(clknet_leaf_6_clk),
    .Q(net467));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[94]$_DFF_P_  (.D(_00287_),
    .CLK(clknet_leaf_7_clk),
    .Q(net468));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[95]$_DFF_P_  (.D(_00288_),
    .CLK(clknet_leaf_7_clk),
    .Q(net469));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[96]$_DFF_P_  (.D(_00161_),
    .CLK(clknet_leaf_13_clk),
    .Q(net470));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[97]$_DFF_P_  (.D(_00162_),
    .CLK(clknet_leaf_13_clk),
    .Q(net471));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[98]$_DFF_P_  (.D(_00163_),
    .CLK(clknet_leaf_13_clk),
    .Q(net472));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[99]$_DFF_P_  (.D(_00164_),
    .CLK(clknet_leaf_13_clk),
    .Q(net473));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[9]$_DFF_P_  (.D(_00194_),
    .CLK(clknet_leaf_21_clk),
    .Q(net474));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[24]$_SDFF_PP1_  (.D(_00537_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.out[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[25]$_SDFF_PP0_  (.D(_00538_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.out[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[26]$_SDFF_PP0_  (.D(_00539_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.out[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[27]$_SDFF_PP0_  (.D(_00540_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.out[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[28]$_SDFF_PP0_  (.D(_00541_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.out[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[29]$_SDFF_PP0_  (.D(_00542_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.r0.out[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[30]$_SDFF_PP0_  (.D(_00543_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.r0.out[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[31]$_SDFF_PP0_  (.D(_00544_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.r0.out[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[0]$_SDFF_PP0_  (.D(_00545_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.r0.rcnt[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[1]$_SDFF_PP0_  (.D(_00546_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.r0.rcnt[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[2]$_SDFF_PP0_  (.D(_00547_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.rcnt[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[3]$_SDFF_PP0_  (.D(_00548_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.r0.rcnt[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[0]$_DFF_P_  (.D(_00000_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.subword[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[1]$_DFF_P_  (.D(_00001_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[2]$_DFF_P_  (.D(_00002_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[3]$_DFF_P_  (.D(_00003_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[4]$_DFF_P_  (.D(_00004_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[5]$_DFF_P_  (.D(_00005_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[6]$_DFF_P_  (.D(_00006_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[7]$_DFF_P_  (.D(_00007_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[0]$_DFF_P_  (.D(_00008_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.subword[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.u1.d[1]$_DFF_P_  (.D(_00009_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.subword[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[2]$_DFF_P_  (.D(_00010_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[3]$_DFF_P_  (.D(_00011_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[4]$_DFF_P_  (.D(_00012_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[5]$_DFF_P_  (.D(_00013_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[6]$_DFF_P_  (.D(_00014_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.subword[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[7]$_DFF_P_  (.D(_00015_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.subword[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[0]$_DFF_P_  (.D(_00016_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.subword[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[1]$_DFF_P_  (.D(_00017_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.subword[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[2]$_DFF_P_  (.D(_00018_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.subword[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[3]$_DFF_P_  (.D(_00019_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.subword[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[4]$_DFF_P_  (.D(_00020_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.subword[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[5]$_DFF_P_  (.D(_00021_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.subword[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[6]$_DFF_P_  (.D(_00022_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.subword[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[7]$_DFF_P_  (.D(_00023_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.subword[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[0]$_DFF_P_  (.D(_00024_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.subword[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.u3.d[1]$_DFF_P_  (.D(_00025_),
    .CLK(clknet_leaf_4_clk),
    .Q(\u0.subword[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[2]$_DFF_P_  (.D(_00026_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.subword[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[3]$_DFF_P_  (.D(_00027_),
    .CLK(clknet_leaf_4_clk),
    .Q(\u0.subword[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[4]$_DFF_P_  (.D(_00028_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.subword[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[5]$_DFF_P_  (.D(_00029_),
    .CLK(clknet_leaf_4_clk),
    .Q(\u0.subword[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[6]$_DFF_P_  (.D(_00030_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.subword[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[7]$_DFF_P_  (.D(_00031_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.subword[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][0]$_DFF_P_  (.D(_00289_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][10]$_DFF_P_  (.D(_00290_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][11]$_DFF_P_  (.D(_00291_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][12]$_DFF_P_  (.D(_00292_),
    .CLK(clknet_leaf_23_clk),
    .Q(\u0.w[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][13]$_DFF_P_  (.D(_00293_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][14]$_DFF_P_  (.D(_00294_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][15]$_DFF_P_  (.D(_00295_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][16]$_DFF_P_  (.D(_00296_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][17]$_DFF_P_  (.D(_00297_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][18]$_DFF_P_  (.D(_00298_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][19]$_DFF_P_  (.D(_00299_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][1]$_DFF_P_  (.D(_00300_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][20]$_DFF_P_  (.D(_00301_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][21]$_DFF_P_  (.D(_00302_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][22]$_DFF_P_  (.D(_00303_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][23]$_DFF_P_  (.D(_00304_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][24]$_DFF_P_  (.D(_00305_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][25]$_DFF_P_  (.D(_00306_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][26]$_DFF_P_  (.D(_00307_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][27]$_DFF_P_  (.D(_00308_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][28]$_DFF_P_  (.D(_00309_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][29]$_DFF_P_  (.D(_00310_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][2]$_DFF_P_  (.D(_00311_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][30]$_DFF_P_  (.D(_00312_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.w[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][31]$_DFF_P_  (.D(_00313_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.w[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][3]$_DFF_P_  (.D(_00314_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][4]$_DFF_P_  (.D(_00315_),
    .CLK(clknet_leaf_17_clk),
    .Q(\u0.w[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][5]$_DFF_P_  (.D(_00316_),
    .CLK(clknet_leaf_4_clk),
    .Q(\u0.w[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][6]$_DFF_P_  (.D(_00317_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][7]$_DFF_P_  (.D(_00318_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][8]$_DFF_P_  (.D(_00319_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[0][9]$_DFF_P_  (.D(_00320_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][0]$_DFF_P_  (.D(_00321_),
    .CLK(clknet_leaf_12_clk),
    .Q(\u0.w[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][10]$_DFF_P_  (.D(_00322_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][11]$_DFF_P_  (.D(_00323_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][12]$_DFF_P_  (.D(_00324_),
    .CLK(clknet_leaf_23_clk),
    .Q(\u0.w[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][13]$_DFF_P_  (.D(_00325_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][14]$_DFF_P_  (.D(_00326_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][15]$_DFF_P_  (.D(_00327_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][16]$_DFF_P_  (.D(_00328_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][17]$_DFF_P_  (.D(_00329_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][18]$_DFF_P_  (.D(_00330_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][19]$_DFF_P_  (.D(_00331_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][1]$_DFF_P_  (.D(_00332_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][20]$_DFF_P_  (.D(_00333_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][21]$_DFF_P_  (.D(_00334_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][22]$_DFF_P_  (.D(_00335_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][23]$_DFF_P_  (.D(_00336_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][24]$_DFF_P_  (.D(_00337_),
    .CLK(clknet_leaf_5_clk),
    .Q(\u0.w[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][25]$_DFF_P_  (.D(_00338_),
    .CLK(clknet_leaf_5_clk),
    .Q(\u0.w[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][26]$_DFF_P_  (.D(_00339_),
    .CLK(clknet_leaf_5_clk),
    .Q(\u0.w[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][27]$_DFF_P_  (.D(_00340_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][28]$_DFF_P_  (.D(_00341_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][29]$_DFF_P_  (.D(_00342_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.w[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][2]$_DFF_P_  (.D(_00343_),
    .CLK(clknet_leaf_12_clk),
    .Q(\u0.w[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][30]$_DFF_P_  (.D(_00344_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.w[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][31]$_DFF_P_  (.D(_00345_),
    .CLK(clknet_leaf_7_clk),
    .Q(\u0.w[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][3]$_DFF_P_  (.D(_00346_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][4]$_DFF_P_  (.D(_00347_),
    .CLK(clknet_leaf_17_clk),
    .Q(\u0.w[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][5]$_DFF_P_  (.D(_00348_),
    .CLK(clknet_leaf_4_clk),
    .Q(\u0.w[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][6]$_DFF_P_  (.D(_00349_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][7]$_DFF_P_  (.D(_00350_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][8]$_DFF_P_  (.D(_00351_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[1][9]$_DFF_P_  (.D(_00352_),
    .CLK(clknet_leaf_25_clk),
    .Q(\u0.w[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][0]$_DFF_P_  (.D(_00353_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][10]$_DFF_P_  (.D(_00354_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][11]$_DFF_P_  (.D(_00355_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.w[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][12]$_DFF_P_  (.D(_00356_),
    .CLK(clknet_leaf_17_clk),
    .Q(\u0.w[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][13]$_DFF_P_  (.D(_00357_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][14]$_DFF_P_  (.D(_00358_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][15]$_DFF_P_  (.D(_00359_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][16]$_DFF_P_  (.D(_00360_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][17]$_DFF_P_  (.D(_00361_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][18]$_DFF_P_  (.D(_00362_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][19]$_DFF_P_  (.D(_00363_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][1]$_DFF_P_  (.D(_00364_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][20]$_DFF_P_  (.D(_00365_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][21]$_DFF_P_  (.D(_00366_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][22]$_DFF_P_  (.D(_00367_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][23]$_DFF_P_  (.D(_00368_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][24]$_DFF_P_  (.D(_00369_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][25]$_DFF_P_  (.D(_00370_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][26]$_DFF_P_  (.D(_00371_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][27]$_DFF_P_  (.D(_00372_),
    .CLK(clknet_leaf_6_clk),
    .Q(\u0.w[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][28]$_DFF_P_  (.D(_00373_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.w[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][29]$_DFF_P_  (.D(_00374_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][2]$_DFF_P_  (.D(_00375_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][30]$_DFF_P_  (.D(_00376_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.w[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][31]$_DFF_P_  (.D(_00377_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][3]$_DFF_P_  (.D(_00378_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][4]$_DFF_P_  (.D(_00379_),
    .CLK(clknet_leaf_17_clk),
    .Q(\u0.w[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][5]$_DFF_P_  (.D(_00380_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][6]$_DFF_P_  (.D(_00381_),
    .CLK(clknet_leaf_17_clk),
    .Q(\u0.w[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][7]$_DFF_P_  (.D(_00382_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.w[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][8]$_DFF_P_  (.D(_00383_),
    .CLK(clknet_leaf_17_clk),
    .Q(\u0.w[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[2][9]$_DFF_P_  (.D(_00384_),
    .CLK(clknet_leaf_25_clk),
    .Q(\u0.w[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][0]$_DFF_P_  (.D(net87),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.tmp_w[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][10]$_DFF_P_  (.D(_15596_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][11]$_DFF_P_  (.D(_00385_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][12]$_DFF_P_  (.D(_00386_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][13]$_DFF_P_  (.D(_00387_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][14]$_DFF_P_  (.D(_00388_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][15]$_DFF_P_  (.D(_00389_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][16]$_DFF_P_  (.D(net5),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][17]$_DFF_P_  (.D(net6),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][18]$_DFF_P_  (.D(_15562_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][19]$_DFF_P_  (.D(_00390_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][1]$_DFF_P_  (.D(net86),
    .CLK(clknet_leaf_23_clk),
    .Q(\u0.tmp_w[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][20]$_DFF_P_  (.D(_00391_),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][21]$_DFF_P_  (.D(_00392_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.tmp_w[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][22]$_DFF_P_  (.D(_00393_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.tmp_w[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][23]$_DFF_P_  (.D(_00394_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.tmp_w[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][24]$_DFF_P_  (.D(net25),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][25]$_DFF_P_  (.D(net37),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][26]$_DFF_P_  (.D(_15659_),
    .CLK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][27]$_DFF_P_  (.D(_00395_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][28]$_DFF_P_  (.D(_00396_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][29]$_DFF_P_  (.D(_00397_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][2]$_DFF_P_  (.D(_15630_),
    .CLK(clknet_leaf_23_clk),
    .Q(\u0.tmp_w[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][30]$_DFF_P_  (.D(_00398_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][31]$_DFF_P_  (.D(_00399_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][3]$_DFF_P_  (.D(_00400_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.tmp_w[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][4]$_DFF_P_  (.D(_00401_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.tmp_w[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][5]$_DFF_P_  (.D(_00402_),
    .CLK(clknet_leaf_24_clk),
    .Q(\u0.tmp_w[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][6]$_DFF_P_  (.D(_00403_),
    .CLK(clknet_leaf_23_clk),
    .Q(\u0.tmp_w[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][7]$_DFF_P_  (.D(_00404_),
    .CLK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][8]$_DFF_P_  (.D(net77),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \u0.w[3][9]$_DFF_P_  (.D(net30),
    .CLK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[9] ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone1 (.A1(_11322_),
    .A2(_11321_),
    .ZN(net1));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone2 (.A1(_14445_),
    .A2(net526),
    .ZN(net2));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone3 (.A1(_05267_),
    .A2(_05262_),
    .ZN(net3));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone4 (.A1(_12916_),
    .A2(net780),
    .ZN(net4));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone5 (.A1(_07468_),
    .A2(_07394_),
    .B(_07448_),
    .ZN(net5));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone6 (.A1(net534),
    .A2(_07468_),
    .B(_07471_),
    .ZN(net6));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone7 (.A1(_05390_),
    .A2(_05389_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone8 (.A1(_15079_),
    .A2(_15078_),
    .ZN(net8));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone9 (.A1(_03835_),
    .A2(_03834_),
    .ZN(net9));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone10 (.A1(_15294_),
    .A2(_15293_),
    .ZN(net10));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone11 (.A1(_07688_),
    .A2(_07687_),
    .ZN(net11));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone12 (.A1(net963),
    .A2(_12857_),
    .ZN(net12));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone13 (.A1(_12226_),
    .A2(_12052_),
    .ZN(net13));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone14 (.A1(_14338_),
    .A2(_14337_),
    .ZN(net14));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone15 (.A1(net641),
    .A2(net635),
    .ZN(net15));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone16 (.A1(_00830_),
    .A2(_00829_),
    .ZN(net16));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone17 (.A1(net1171),
    .A2(_12131_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone18 (.A1(net909),
    .A2(net908),
    .ZN(net18));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone19 (.A1(net1134),
    .A2(_13717_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone20 (.I(net1153),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone21 (.A1(net1228),
    .A2(net1230),
    .ZN(net21));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone22 (.A1(_04531_),
    .A2(_04526_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone23 (.I(_06085_),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone24 (.A1(_06060_),
    .A2(_06059_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone25 (.A1(_09736_),
    .A2(_09735_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone26 (.I(net948),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone27 (.A1(_01616_),
    .A2(net862),
    .ZN(net27));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone28 (.A1(_13601_),
    .A2(net1135),
    .ZN(net28));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone29 (.A1(_03061_),
    .A2(_03056_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone30 (.A1(_07404_),
    .A2(_07609_),
    .B(_07612_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone31 (.A1(net813),
    .A2(net804),
    .ZN(net31));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone32 (.A1(_10386_),
    .A2(_10385_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone33 (.A1(net616),
    .A2(_10442_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone34 (.A1(_00875_),
    .A2(_00874_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split35 (.I(\sa01_sr[7] ),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone36 (.A1(net1261),
    .A2(net831),
    .ZN(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 clone37 (.I(_15650_),
    .ZN(net37));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split38 (.I(\sa32_sub[1] ),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 split39 (.I(\sa03_sr[7] ),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer431 (.I(net4),
    .Z(net928));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone41 (.A1(_12806_),
    .A2(_12805_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone42 (.I(net980),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone43 (.I(net520),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone44 (.I(_03156_),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone46 (.I(net678),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone47 (.I(\sa20_sr[7] ),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone48 (.A1(_03043_),
    .A2(_03038_),
    .ZN(net48));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone49 (.I(\sa20_sub[7] ),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split50 (.I(net744),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone51 (.A1(_03880_),
    .A2(_03832_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 clone52 (.A1(_03826_),
    .A2(_03824_),
    .B(\u0.tmp_w[10] ),
    .ZN(net52));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 clone53 (.A1(_03830_),
    .A2(_07615_),
    .A3(_03829_),
    .ZN(net53));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clone54 (.I(\sa32_sub[7] ),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 split57 (.I(net1172),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone58 (.I(net1182),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone59 (.A1(_03811_),
    .A2(_03816_),
    .ZN(net59));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone60 (.A1(_03799_),
    .A2(_03794_),
    .ZN(net60));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone61 (.A1(net1034),
    .A2(_07536_),
    .ZN(net61));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split62 (.I(net817),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer188 (.I(_03122_),
    .Z(net647));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone64 (.A1(_03877_),
    .A2(_03875_),
    .ZN(net64));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clone66 (.I(_02425_),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 clone68 (.I(\sa30_sr[7] ),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clone69 (.I(_02367_),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone70 (.A1(_02390_),
    .A2(_02389_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone71 (.A1(_12049_),
    .A2(_12048_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 split72 (.I(\sa12_sr[7] ),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone73 (.A1(net1082),
    .A2(net1081),
    .ZN(net73));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone74 (.I(_04571_),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split75 (.I(\sa00_sr[0] ),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 split76 (.I(\sa00_sr[7] ),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone77 (.A1(_07467_),
    .A2(_07601_),
    .B(_07604_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone78 (.A1(_07613_),
    .A2(_07610_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone79 (.I(_08603_),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone80 (.A1(_10413_),
    .A2(_10407_),
    .ZN(net80));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone81 (.I(_06726_),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone82 (.A1(_07472_),
    .A2(_07469_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone83 (.A1(_13643_),
    .A2(net692),
    .ZN(net83));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone84 (.I(_08564_),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone85 (.A1(_06799_),
    .A2(_06797_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone86 (.A1(_07542_),
    .A2(_07550_),
    .B(_07553_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone87 (.A1(_07468_),
    .A2(_07541_),
    .B(_07545_),
    .ZN(net87));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone88 (.A1(_07546_),
    .A2(_07543_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone89 (.A1(_07554_),
    .A2(_07551_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone90 (.I(_03833_),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone91 (.I(_03832_),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone92 (.A1(_02301_),
    .A2(_02305_),
    .ZN(net92));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_469 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_470 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_471 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_472 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_473 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_474 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_475 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_476 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_477 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_478 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_479 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_480 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_481 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_482 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_483 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_484 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_485 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_486 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_487 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_488 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_489 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_490 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(key[0]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input2 (.I(key[100]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input3 (.I(key[101]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input4 (.I(key[102]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input5 (.I(key[103]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input6 (.I(key[104]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(key[105]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(key[106]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(key[107]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input10 (.I(key[108]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(key[109]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(key[10]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(key[110]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(key[111]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(key[112]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(key[113]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(key[114]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(key[115]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(key[116]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(key[117]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(key[118]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(key[119]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(key[11]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(key[120]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(key[121]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(key[122]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(key[123]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(key[124]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(key[125]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(key[126]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(key[127]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(key[12]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input33 (.I(key[13]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(key[14]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(key[15]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(key[16]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(key[17]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(key[18]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(key[19]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(key[1]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(key[20]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(key[21]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(key[22]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(key[23]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(key[24]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input46 (.I(key[25]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input47 (.I(key[26]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(key[27]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(key[28]),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(key[29]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input51 (.I(key[2]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(key[30]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(key[31]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input54 (.I(key[32]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input55 (.I(key[33]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input56 (.I(key[34]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input57 (.I(key[35]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input58 (.I(key[36]),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input59 (.I(key[37]),
    .Z(net146));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input60 (.I(key[38]),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input61 (.I(key[39]),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input62 (.I(key[3]),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(key[40]),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input64 (.I(key[41]),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input65 (.I(key[42]),
    .Z(net152));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input66 (.I(key[43]),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input67 (.I(key[44]),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input68 (.I(key[45]),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input69 (.I(key[46]),
    .Z(net156));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input70 (.I(key[47]),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input71 (.I(key[48]),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input72 (.I(key[49]),
    .Z(net159));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input73 (.I(key[4]),
    .Z(net160));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input74 (.I(key[50]),
    .Z(net161));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input75 (.I(key[51]),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input76 (.I(key[52]),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input77 (.I(key[53]),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input78 (.I(key[54]),
    .Z(net165));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input79 (.I(key[55]),
    .Z(net166));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input80 (.I(key[56]),
    .Z(net167));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input81 (.I(key[57]),
    .Z(net168));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input82 (.I(key[58]),
    .Z(net169));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input83 (.I(key[59]),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input84 (.I(key[5]),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input85 (.I(key[60]),
    .Z(net172));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input86 (.I(key[61]),
    .Z(net173));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input87 (.I(key[62]),
    .Z(net174));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input88 (.I(key[63]),
    .Z(net175));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input89 (.I(key[64]),
    .Z(net176));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input90 (.I(key[65]),
    .Z(net177));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input91 (.I(key[66]),
    .Z(net178));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input92 (.I(key[67]),
    .Z(net179));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input93 (.I(key[68]),
    .Z(net180));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input94 (.I(key[69]),
    .Z(net181));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input95 (.I(key[6]),
    .Z(net182));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input96 (.I(key[70]),
    .Z(net183));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input97 (.I(key[71]),
    .Z(net184));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input98 (.I(key[72]),
    .Z(net185));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input99 (.I(key[73]),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input100 (.I(key[74]),
    .Z(net187));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input101 (.I(key[75]),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input102 (.I(key[76]),
    .Z(net189));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input103 (.I(key[77]),
    .Z(net190));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input104 (.I(key[78]),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input105 (.I(key[79]),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input106 (.I(key[7]),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input107 (.I(key[80]),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input108 (.I(key[81]),
    .Z(net195));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input109 (.I(key[82]),
    .Z(net196));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input110 (.I(key[83]),
    .Z(net197));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input111 (.I(key[84]),
    .Z(net198));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input112 (.I(key[85]),
    .Z(net199));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input113 (.I(key[86]),
    .Z(net200));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input114 (.I(key[87]),
    .Z(net201));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input115 (.I(key[88]),
    .Z(net202));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input116 (.I(key[89]),
    .Z(net203));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input117 (.I(key[8]),
    .Z(net204));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input118 (.I(key[90]),
    .Z(net205));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input119 (.I(key[91]),
    .Z(net206));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input120 (.I(key[92]),
    .Z(net207));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input121 (.I(key[93]),
    .Z(net208));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input122 (.I(key[94]),
    .Z(net209));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input123 (.I(key[95]),
    .Z(net210));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input124 (.I(key[96]),
    .Z(net211));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input125 (.I(key[97]),
    .Z(net212));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input126 (.I(key[98]),
    .Z(net213));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input127 (.I(key[99]),
    .Z(net214));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input128 (.I(key[9]),
    .Z(net215));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input129 (.I(ld),
    .Z(net216));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input130 (.I(rst),
    .Z(net217));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input131 (.I(text_in[0]),
    .Z(net218));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input132 (.I(text_in[100]),
    .Z(net219));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input133 (.I(text_in[101]),
    .Z(net220));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input134 (.I(text_in[102]),
    .Z(net221));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input135 (.I(text_in[103]),
    .Z(net222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input136 (.I(text_in[104]),
    .Z(net223));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input137 (.I(text_in[105]),
    .Z(net224));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input138 (.I(text_in[106]),
    .Z(net225));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input139 (.I(text_in[107]),
    .Z(net226));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input140 (.I(text_in[108]),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input141 (.I(text_in[109]),
    .Z(net228));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input142 (.I(text_in[10]),
    .Z(net229));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input143 (.I(text_in[110]),
    .Z(net230));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input144 (.I(text_in[111]),
    .Z(net231));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input145 (.I(text_in[112]),
    .Z(net232));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input146 (.I(text_in[113]),
    .Z(net233));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input147 (.I(text_in[114]),
    .Z(net234));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input148 (.I(text_in[115]),
    .Z(net235));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input149 (.I(text_in[116]),
    .Z(net236));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input150 (.I(text_in[117]),
    .Z(net237));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input151 (.I(text_in[118]),
    .Z(net238));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input152 (.I(text_in[119]),
    .Z(net239));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input153 (.I(text_in[11]),
    .Z(net240));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input154 (.I(text_in[120]),
    .Z(net241));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input155 (.I(text_in[121]),
    .Z(net242));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input156 (.I(text_in[122]),
    .Z(net243));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input157 (.I(text_in[123]),
    .Z(net244));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input158 (.I(text_in[124]),
    .Z(net245));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input159 (.I(text_in[125]),
    .Z(net246));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input160 (.I(text_in[126]),
    .Z(net247));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input161 (.I(text_in[127]),
    .Z(net248));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input162 (.I(text_in[12]),
    .Z(net249));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input163 (.I(text_in[13]),
    .Z(net250));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input164 (.I(text_in[14]),
    .Z(net251));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input165 (.I(text_in[15]),
    .Z(net252));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input166 (.I(text_in[16]),
    .Z(net253));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input167 (.I(text_in[17]),
    .Z(net254));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input168 (.I(text_in[18]),
    .Z(net255));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input169 (.I(text_in[19]),
    .Z(net256));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input170 (.I(text_in[1]),
    .Z(net257));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input171 (.I(text_in[20]),
    .Z(net258));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input172 (.I(text_in[21]),
    .Z(net259));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input173 (.I(text_in[22]),
    .Z(net260));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input174 (.I(text_in[23]),
    .Z(net261));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input175 (.I(text_in[24]),
    .Z(net262));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input176 (.I(text_in[25]),
    .Z(net263));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input177 (.I(text_in[26]),
    .Z(net264));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input178 (.I(text_in[27]),
    .Z(net265));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input179 (.I(text_in[28]),
    .Z(net266));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input180 (.I(text_in[29]),
    .Z(net267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input181 (.I(text_in[2]),
    .Z(net268));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input182 (.I(text_in[30]),
    .Z(net269));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input183 (.I(text_in[31]),
    .Z(net270));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input184 (.I(text_in[32]),
    .Z(net271));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input185 (.I(text_in[33]),
    .Z(net272));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input186 (.I(text_in[34]),
    .Z(net273));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input187 (.I(text_in[35]),
    .Z(net274));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input188 (.I(text_in[36]),
    .Z(net275));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input189 (.I(text_in[37]),
    .Z(net276));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input190 (.I(text_in[38]),
    .Z(net277));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input191 (.I(text_in[39]),
    .Z(net278));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input192 (.I(text_in[3]),
    .Z(net279));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input193 (.I(text_in[40]),
    .Z(net280));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input194 (.I(text_in[41]),
    .Z(net281));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input195 (.I(text_in[42]),
    .Z(net282));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input196 (.I(text_in[43]),
    .Z(net283));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input197 (.I(text_in[44]),
    .Z(net284));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input198 (.I(text_in[45]),
    .Z(net285));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input199 (.I(text_in[46]),
    .Z(net286));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input200 (.I(text_in[47]),
    .Z(net287));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input201 (.I(text_in[48]),
    .Z(net288));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input202 (.I(text_in[49]),
    .Z(net289));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input203 (.I(text_in[4]),
    .Z(net290));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input204 (.I(text_in[50]),
    .Z(net291));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input205 (.I(text_in[51]),
    .Z(net292));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input206 (.I(text_in[52]),
    .Z(net293));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input207 (.I(text_in[53]),
    .Z(net294));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input208 (.I(text_in[54]),
    .Z(net295));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input209 (.I(text_in[55]),
    .Z(net296));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input210 (.I(text_in[56]),
    .Z(net297));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input211 (.I(text_in[57]),
    .Z(net298));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input212 (.I(text_in[58]),
    .Z(net299));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input213 (.I(text_in[59]),
    .Z(net300));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input214 (.I(text_in[5]),
    .Z(net301));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input215 (.I(text_in[60]),
    .Z(net302));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input216 (.I(text_in[61]),
    .Z(net303));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input217 (.I(text_in[62]),
    .Z(net304));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input218 (.I(text_in[63]),
    .Z(net305));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input219 (.I(text_in[64]),
    .Z(net306));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input220 (.I(text_in[65]),
    .Z(net307));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input221 (.I(text_in[66]),
    .Z(net308));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input222 (.I(text_in[67]),
    .Z(net309));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input223 (.I(text_in[68]),
    .Z(net310));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input224 (.I(text_in[69]),
    .Z(net311));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input225 (.I(text_in[6]),
    .Z(net312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input226 (.I(text_in[70]),
    .Z(net313));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input227 (.I(text_in[71]),
    .Z(net314));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input228 (.I(text_in[72]),
    .Z(net315));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input229 (.I(text_in[73]),
    .Z(net316));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input230 (.I(text_in[74]),
    .Z(net317));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input231 (.I(text_in[75]),
    .Z(net318));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input232 (.I(text_in[76]),
    .Z(net319));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input233 (.I(text_in[77]),
    .Z(net320));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input234 (.I(text_in[78]),
    .Z(net321));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input235 (.I(text_in[79]),
    .Z(net322));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input236 (.I(text_in[7]),
    .Z(net323));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input237 (.I(text_in[80]),
    .Z(net324));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input238 (.I(text_in[81]),
    .Z(net325));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input239 (.I(text_in[82]),
    .Z(net326));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input240 (.I(text_in[83]),
    .Z(net327));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input241 (.I(text_in[84]),
    .Z(net328));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input242 (.I(text_in[85]),
    .Z(net329));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input243 (.I(text_in[86]),
    .Z(net330));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input244 (.I(text_in[87]),
    .Z(net331));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input245 (.I(text_in[88]),
    .Z(net332));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input246 (.I(text_in[89]),
    .Z(net333));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input247 (.I(text_in[8]),
    .Z(net334));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input248 (.I(text_in[90]),
    .Z(net335));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input249 (.I(text_in[91]),
    .Z(net336));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input250 (.I(text_in[92]),
    .Z(net337));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input251 (.I(text_in[93]),
    .Z(net338));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input252 (.I(text_in[94]),
    .Z(net339));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input253 (.I(text_in[95]),
    .Z(net340));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input254 (.I(text_in[96]),
    .Z(net341));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input255 (.I(text_in[97]),
    .Z(net342));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input256 (.I(text_in[98]),
    .Z(net343));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input257 (.I(text_in[99]),
    .Z(net344));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input258 (.I(text_in[9]),
    .Z(net345));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output259 (.I(net346),
    .Z(done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output260 (.I(net347),
    .Z(text_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output261 (.I(net348),
    .Z(text_out[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output262 (.I(net349),
    .Z(text_out[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output263 (.I(net350),
    .Z(text_out[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output264 (.I(net351),
    .Z(text_out[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output265 (.I(net352),
    .Z(text_out[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output266 (.I(net353),
    .Z(text_out[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output267 (.I(net354),
    .Z(text_out[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output268 (.I(net355),
    .Z(text_out[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output269 (.I(net356),
    .Z(text_out[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output270 (.I(net357),
    .Z(text_out[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output271 (.I(net358),
    .Z(text_out[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output272 (.I(net359),
    .Z(text_out[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output273 (.I(net360),
    .Z(text_out[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output274 (.I(net361),
    .Z(text_out[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output275 (.I(net362),
    .Z(text_out[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output276 (.I(net363),
    .Z(text_out[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output277 (.I(net364),
    .Z(text_out[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output278 (.I(net365),
    .Z(text_out[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output279 (.I(net366),
    .Z(text_out[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output280 (.I(net367),
    .Z(text_out[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output281 (.I(net368),
    .Z(text_out[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output282 (.I(net369),
    .Z(text_out[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output283 (.I(net370),
    .Z(text_out[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output284 (.I(net371),
    .Z(text_out[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output285 (.I(net372),
    .Z(text_out[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output286 (.I(net373),
    .Z(text_out[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output287 (.I(net374),
    .Z(text_out[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output288 (.I(net375),
    .Z(text_out[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output289 (.I(net376),
    .Z(text_out[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output290 (.I(net377),
    .Z(text_out[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output291 (.I(net378),
    .Z(text_out[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output292 (.I(net379),
    .Z(text_out[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output293 (.I(net380),
    .Z(text_out[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output294 (.I(net381),
    .Z(text_out[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output295 (.I(net382),
    .Z(text_out[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output296 (.I(net383),
    .Z(text_out[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output297 (.I(net384),
    .Z(text_out[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output298 (.I(net385),
    .Z(text_out[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output299 (.I(net386),
    .Z(text_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output300 (.I(net387),
    .Z(text_out[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output301 (.I(net388),
    .Z(text_out[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output302 (.I(net389),
    .Z(text_out[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output303 (.I(net390),
    .Z(text_out[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output304 (.I(net391),
    .Z(text_out[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output305 (.I(net392),
    .Z(text_out[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output306 (.I(net393),
    .Z(text_out[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output307 (.I(net394),
    .Z(text_out[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output308 (.I(net395),
    .Z(text_out[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output309 (.I(net396),
    .Z(text_out[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output310 (.I(net397),
    .Z(text_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output311 (.I(net398),
    .Z(text_out[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output312 (.I(net399),
    .Z(text_out[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output313 (.I(net400),
    .Z(text_out[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output314 (.I(net401),
    .Z(text_out[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output315 (.I(net402),
    .Z(text_out[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output316 (.I(net403),
    .Z(text_out[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output317 (.I(net404),
    .Z(text_out[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output318 (.I(net405),
    .Z(text_out[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output319 (.I(net406),
    .Z(text_out[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output320 (.I(net407),
    .Z(text_out[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output321 (.I(net408),
    .Z(text_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output322 (.I(net409),
    .Z(text_out[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output323 (.I(net410),
    .Z(text_out[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output324 (.I(net411),
    .Z(text_out[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output325 (.I(net412),
    .Z(text_out[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output326 (.I(net413),
    .Z(text_out[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output327 (.I(net414),
    .Z(text_out[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output328 (.I(net415),
    .Z(text_out[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output329 (.I(net416),
    .Z(text_out[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output330 (.I(net417),
    .Z(text_out[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output331 (.I(net418),
    .Z(text_out[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output332 (.I(net419),
    .Z(text_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output333 (.I(net420),
    .Z(text_out[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output334 (.I(net421),
    .Z(text_out[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output335 (.I(net422),
    .Z(text_out[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output336 (.I(net423),
    .Z(text_out[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output337 (.I(net424),
    .Z(text_out[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output338 (.I(net425),
    .Z(text_out[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output339 (.I(net426),
    .Z(text_out[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output340 (.I(net427),
    .Z(text_out[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output341 (.I(net428),
    .Z(text_out[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output342 (.I(net429),
    .Z(text_out[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output343 (.I(net430),
    .Z(text_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output344 (.I(net431),
    .Z(text_out[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output345 (.I(net432),
    .Z(text_out[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output346 (.I(net433),
    .Z(text_out[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output347 (.I(net434),
    .Z(text_out[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output348 (.I(net435),
    .Z(text_out[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output349 (.I(net436),
    .Z(text_out[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output350 (.I(net437),
    .Z(text_out[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output351 (.I(net438),
    .Z(text_out[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output352 (.I(net439),
    .Z(text_out[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output353 (.I(net440),
    .Z(text_out[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output354 (.I(net441),
    .Z(text_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output355 (.I(net442),
    .Z(text_out[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output356 (.I(net443),
    .Z(text_out[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output357 (.I(net444),
    .Z(text_out[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output358 (.I(net445),
    .Z(text_out[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output359 (.I(net446),
    .Z(text_out[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output360 (.I(net447),
    .Z(text_out[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output361 (.I(net448),
    .Z(text_out[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output362 (.I(net449),
    .Z(text_out[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output363 (.I(net450),
    .Z(text_out[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output364 (.I(net451),
    .Z(text_out[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output365 (.I(net452),
    .Z(text_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output366 (.I(net453),
    .Z(text_out[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output367 (.I(net454),
    .Z(text_out[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output368 (.I(net455),
    .Z(text_out[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output369 (.I(net456),
    .Z(text_out[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output370 (.I(net457),
    .Z(text_out[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output371 (.I(net458),
    .Z(text_out[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output372 (.I(net459),
    .Z(text_out[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output373 (.I(net460),
    .Z(text_out[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output374 (.I(net461),
    .Z(text_out[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output375 (.I(net462),
    .Z(text_out[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output376 (.I(net463),
    .Z(text_out[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output377 (.I(net464),
    .Z(text_out[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output378 (.I(net465),
    .Z(text_out[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output379 (.I(net466),
    .Z(text_out[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output380 (.I(net467),
    .Z(text_out[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output381 (.I(net468),
    .Z(text_out[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output382 (.I(net469),
    .Z(text_out[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output383 (.I(net470),
    .Z(text_out[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output384 (.I(net471),
    .Z(text_out[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output385 (.I(net472),
    .Z(text_out[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output386 (.I(net473),
    .Z(text_out[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output387 (.I(net474),
    .Z(text_out[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 clkload1 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload2 (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload3 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload4 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload5 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload6 (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkload7 (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload8 (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload9 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload10 (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload11 (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload12 (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload13 (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload14 (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload15 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload16 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload17 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload18 (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload19 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload20 (.I(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload21 (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload22 (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload23 (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload24 (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload25 (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload26 (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer1 (.I(ld_r),
    .Z(net475));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer2 (.I(net475),
    .Z(net476));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer3 (.I(ld_r),
    .Z(net477));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer4 (.I(net477),
    .Z(net478));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer41 (.I(_15834_),
    .Z(net503));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer42 (.I(_15834_),
    .Z(net504));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer43 (.I(net504),
    .Z(net505));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer44 (.I(net505),
    .Z(net506));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer45 (.I(_15836_),
    .Z(net507));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer46 (.I(_15836_),
    .Z(net508));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone50 (.A1(_14384_),
    .A2(net503),
    .ZN(net509));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer51 (.I(_14438_),
    .Z(net510));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer52 (.I(net555),
    .Z(net511));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer53 (.I(_14334_),
    .Z(net512));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer54 (.I(net1273),
    .Z(net513));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer55 (.I(_14551_),
    .Z(net514));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer56 (.I(_14551_),
    .Z(net515));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer57 (.I(\sa30_sub[0] ),
    .Z(net516));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer58 (.I(net516),
    .Z(net517));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer59 (.I(\sa30_sub[0] ),
    .Z(net518));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer60 (.I(net518),
    .Z(net519));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer61 (.I(\sa11_sr[7] ),
    .Z(net520));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer62 (.I(_14351_),
    .Z(net521));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer63 (.I(_15833_),
    .Z(net522));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer64 (.I(net43),
    .Z(net523));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer65 (.I(net523),
    .Z(net524));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer66 (.I(net524),
    .Z(net525));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer67 (.I(_14444_),
    .Z(net526));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer92 (.I(_14317_),
    .Z(net551));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer93 (.I(_15839_),
    .Z(net552));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer94 (.I(net552),
    .Z(net553));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer95 (.I(net553),
    .Z(net554));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer96 (.I(net552),
    .Z(net555));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer114 (.I(\sa20_sr[0] ),
    .Z(net573));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer115 (.I(\sa20_sr[0] ),
    .Z(net574));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer116 (.I(\sa10_sr[0] ),
    .Z(net575));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer117 (.I(\sa10_sr[0] ),
    .Z(net576));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer118 (.I(\sa20_sr[0] ),
    .Z(net577));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer119 (.I(_16076_),
    .Z(net578));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer120 (.I(_04663_),
    .Z(net579));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer121 (.I(\sa30_sr[0] ),
    .Z(net580));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer122 (.I(net617),
    .Z(net581));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer123 (.I(\sa30_sr[0] ),
    .Z(net582));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer124 (.I(\sa30_sr[0] ),
    .Z(net583));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer125 (.I(\sa30_sr[0] ),
    .Z(net584));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer132 (.I(_10622_),
    .Z(net591));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer133 (.I(net591),
    .Z(net592));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer134 (.I(net591),
    .Z(net593));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer135 (.I(_10409_),
    .Z(net594));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer136 (.I(net594),
    .Z(net595));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer137 (.I(_10409_),
    .Z(net596));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer138 (.I(_15673_),
    .Z(net597));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer139 (.I(_15673_),
    .Z(net598));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer140 (.I(_15679_),
    .Z(net599));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer141 (.I(net599),
    .Z(net600));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer142 (.I(net599),
    .Z(net601));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer143 (.I(net601),
    .Z(net602));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer144 (.I(_10444_),
    .Z(net603));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer145 (.I(_10444_),
    .Z(net604));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer146 (.I(net1079),
    .Z(net605));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer147 (.I(\sa30_sr[1] ),
    .Z(net606));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer148 (.I(net690),
    .Z(net607));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer149 (.I(_15676_),
    .Z(net608));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 rebuffer150 (.I(_10536_),
    .Z(net609));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer151 (.I(_15674_),
    .Z(net610));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer152 (.I(net610),
    .Z(net611));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer153 (.I(_15674_),
    .Z(net612));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer154 (.I(\sa20_sr[1] ),
    .Z(net613));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer155 (.I(\sa20_sr[1] ),
    .Z(net614));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer156 (.I(\sa20_sr[1] ),
    .Z(net615));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer157 (.I(_10441_),
    .Z(net616));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer173 (.I(_16012_),
    .Z(net632));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer174 (.I(_15064_),
    .Z(net633));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer175 (.I(_16004_),
    .Z(net634));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer176 (.I(_03080_),
    .Z(net635));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer177 (.I(_16002_),
    .Z(net636));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer178 (.I(net636),
    .Z(net637));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer179 (.I(_16001_),
    .Z(net638));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer180 (.I(net638),
    .Z(net639));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer181 (.I(net638),
    .Z(net640));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer182 (.I(_03079_),
    .Z(net641));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer183 (.I(net649),
    .Z(net642));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer184 (.I(\sa31_sub[7] ),
    .Z(net643));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer185 (.I(_03174_),
    .Z(net644));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone186 (.I(_03174_),
    .Z(net645));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone187 (.I(_03174_),
    .Z(net646));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer189 (.I(_03122_),
    .Z(net648));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer190 (.I(net650),
    .Z(net649));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer191 (.I(net651),
    .Z(net650));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer192 (.I(\sa31_sub[7] ),
    .Z(net651));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer197 (.I(net1136),
    .Z(net656));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer198 (.I(net676),
    .Z(net657));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer199 (.I(net657),
    .Z(net658));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer200 (.I(_13706_),
    .Z(net659));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer201 (.I(_15810_),
    .Z(net660));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer202 (.I(net660),
    .Z(net661));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer203 (.I(net661),
    .Z(net662));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer204 (.I(net662),
    .Z(net663));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer205 (.I(_15810_),
    .Z(net664));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer206 (.I(net664),
    .Z(net665));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer207 (.I(net665),
    .Z(net666));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer208 (.I(net665),
    .Z(net667));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer209 (.I(_15804_),
    .Z(net668));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer210 (.I(_15804_),
    .Z(net669));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer211 (.I(_15801_),
    .Z(net670));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer212 (.I(_15801_),
    .Z(net671));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer213 (.I(_13642_),
    .Z(net672));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer214 (.I(_13597_),
    .Z(net673));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer215 (.I(_13647_),
    .Z(net674));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer216 (.I(_13647_),
    .Z(net675));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer217 (.I(_15807_),
    .Z(net676));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer218 (.I(net676),
    .Z(net677));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer219 (.I(\sa10_sr[7] ),
    .Z(net678));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer220 (.I(\sa10_sr[0] ),
    .Z(net679));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer221 (.I(_13836_),
    .Z(net680));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer222 (.I(_10360_),
    .Z(net681));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer223 (.I(net681),
    .Z(net682));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer224 (.I(net682),
    .Z(net683));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer225 (.I(_13714_),
    .Z(net684));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer226 (.I(_13714_),
    .Z(net685));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer227 (.I(_13647_),
    .Z(net686));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer228 (.I(\sa30_sr[1] ),
    .Z(net687));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer229 (.I(\sa30_sr[1] ),
    .Z(net688));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer230 (.I(_10354_),
    .Z(net689));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer231 (.I(\sa30_sr[1] ),
    .Z(net690));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer232 (.I(_10347_),
    .Z(net691));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer233 (.I(_13644_),
    .Z(net692));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer234 (.I(net83),
    .Z(net693));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer235 (.I(net693),
    .Z(net694));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer236 (.I(\sa00_sr[0] ),
    .Z(net695));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer242 (.I(_03087_),
    .Z(net701));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone243 (.I(_03151_),
    .Z(net702));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone244 (.I(_03122_),
    .Z(net703));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone245 (.I(_03152_),
    .Z(net704));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer246 (.I(_03252_),
    .Z(net705));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer253 (.I(_03903_),
    .Z(net712));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer254 (.I(_16037_),
    .Z(net713));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer255 (.I(net713),
    .Z(net714));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer256 (.I(\sa03_sr[0] ),
    .Z(net715));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer257 (.I(net717),
    .Z(net716));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer258 (.I(net723),
    .Z(net717));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer259 (.I(net748),
    .Z(net718));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer260 (.I(net725),
    .Z(net719));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer261 (.I(\sa03_sr[0] ),
    .Z(net720));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer262 (.I(\sa03_sr[0] ),
    .Z(net721));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer263 (.I(\sa10_sub[0] ),
    .Z(net722));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer264 (.I(\sa03_sr[0] ),
    .Z(net723));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer265 (.I(_16037_),
    .Z(net724));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer266 (.I(_16037_),
    .Z(net725));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer267 (.I(\sa03_sr[0] ),
    .Z(net726));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer268 (.I(\sa03_sr[0] ),
    .Z(net727));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer269 (.I(_03831_),
    .Z(net728));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer270 (.I(net728),
    .Z(net729));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer271 (.I(_04024_),
    .Z(net730));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer272 (.I(net730),
    .Z(net731));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer273 (.I(_16040_),
    .Z(net732));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer274 (.I(\sa10_sub[1] ),
    .Z(net733));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer275 (.I(\sa10_sub[1] ),
    .Z(net734));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer276 (.I(net734),
    .Z(net735));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer277 (.I(\sa10_sub[1] ),
    .Z(net736));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer278 (.I(\sa03_sr[1] ),
    .Z(net737));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer279 (.I(\sa03_sr[1] ),
    .Z(net738));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer280 (.I(\sa03_sr[1] ),
    .Z(net739));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer281 (.I(_16038_),
    .Z(net740));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer282 (.I(net740),
    .Z(net741));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer283 (.I(_03827_),
    .Z(net742));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer284 (.I(_16040_),
    .Z(net743));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer285 (.I(\sa21_sub[7] ),
    .Z(net744));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer286 (.I(net744),
    .Z(net745));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer287 (.I(\sa32_sub[0] ),
    .Z(net746));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer288 (.I(_04233_),
    .Z(net747));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer289 (.I(_16037_),
    .Z(net748));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer290 (.I(_03813_),
    .Z(net749));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer291 (.I(_16048_),
    .Z(net750));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer292 (.I(net754),
    .Z(net751));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer293 (.I(_03891_),
    .Z(net752));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer294 (.I(_03891_),
    .Z(net753));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer295 (.I(_03891_),
    .Z(net754));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer296 (.I(_00881_),
    .Z(net755));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer297 (.I(_03783_),
    .Z(net756));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer328 (.I(\sa31_sub[0] ),
    .Z(net787));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer329 (.I(net789),
    .Z(net788));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer330 (.I(\sa31_sub[0] ),
    .Z(net789));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer335 (.I(_15965_),
    .Z(net794));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer336 (.I(\sa11_sr[0] ),
    .Z(net795));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer337 (.I(\sa11_sr[0] ),
    .Z(net796));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer338 (.I(_15966_),
    .Z(net797));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer339 (.I(\sa01_sr[0] ),
    .Z(net798));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer340 (.I(\sa01_sr[0] ),
    .Z(net799));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer341 (.I(\sa01_sr[0] ),
    .Z(net800));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer342 (.I(_15968_),
    .Z(net801));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer343 (.I(_15968_),
    .Z(net802));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer344 (.I(_02388_),
    .Z(net803));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer345 (.I(net821),
    .Z(net804));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer346 (.I(\sa11_sr[1] ),
    .Z(net805));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer347 (.I(net805),
    .Z(net806));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer348 (.I(\sa11_sr[1] ),
    .Z(net807));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer349 (.I(\sa11_sr[1] ),
    .Z(net808));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer350 (.I(_02303_),
    .Z(net809));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone351 (.I(_02401_),
    .Z(net810));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone352 (.I(_10378_),
    .Z(net811));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer353 (.I(\sa01_sr[0] ),
    .Z(net812));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer354 (.I(_02338_),
    .Z(net813));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer355 (.I(\sa21_sr[0] ),
    .Z(net814));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer356 (.I(\sa21_sr[0] ),
    .Z(net815));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer357 (.I(\sa30_sub[7] ),
    .Z(net816));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer358 (.I(net816),
    .Z(net817));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer359 (.I(net817),
    .Z(net818));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer360 (.I(net62),
    .Z(net819));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer361 (.I(_02391_),
    .Z(net820));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer362 (.I(_02339_),
    .Z(net821));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer367 (.I(_10613_),
    .Z(net826));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer368 (.I(_10380_),
    .Z(net827));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer369 (.I(_15682_),
    .Z(net828));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer370 (.I(net828),
    .Z(net829));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer371 (.I(net828),
    .Z(net830));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer372 (.I(_10665_),
    .Z(net831));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer375 (.I(_15871_),
    .Z(net834));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer376 (.I(_15871_),
    .Z(net835));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer377 (.I(net835),
    .Z(net836));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer378 (.I(_15175_),
    .Z(net837));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer407 (.I(_10362_),
    .Z(net866));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer408 (.I(_13753_),
    .Z(net867));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer409 (.I(_13615_),
    .Z(net868));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer410 (.I(_13615_),
    .Z(net869));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer411 (.I(_13801_),
    .Z(net870));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer412 (.I(_13845_),
    .Z(net871));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone413 (.I(net873),
    .Z(net872));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer414 (.I(_13642_),
    .Z(net873));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer415 (.I(\sa20_sr[1] ),
    .Z(net874));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer416 (.I(\sa20_sr[1] ),
    .Z(net875));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer417 (.I(_10345_),
    .Z(net876));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer418 (.I(_03162_),
    .Z(net877));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer419 (.I(net877),
    .Z(net878));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer420 (.I(_03169_),
    .Z(net879));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer421 (.I(_03169_),
    .Z(net880));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer422 (.I(_03367_),
    .Z(net881));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer423 (.I(net881),
    .Z(net882));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer424 (.I(_03276_),
    .Z(net883));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer425 (.I(_16002_),
    .Z(net884));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer441 (.I(_16170_),
    .Z(net900));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer442 (.I(_06762_),
    .Z(net901));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer443 (.I(_06762_),
    .Z(net902));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer444 (.I(_06762_),
    .Z(net903));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer445 (.I(net903),
    .Z(net904));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer446 (.I(_06896_),
    .Z(net905));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer447 (.I(_16172_),
    .Z(net906));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer448 (.I(_06713_),
    .Z(net907));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer449 (.I(_06918_),
    .Z(net908));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer450 (.I(_06917_),
    .Z(net909));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer451 (.I(_06757_),
    .Z(net910));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer452 (.I(\sa32_sub[1] ),
    .Z(net911));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer453 (.I(_06726_),
    .Z(net912));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone454 (.A1(_16169_),
    .A2(net912),
    .ZN(net913));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer455 (.I(_12774_),
    .Z(net914));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone484 (.I(_02384_),
    .Z(net943));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer485 (.I(_02549_),
    .Z(net944));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer487 (.I(net533),
    .Z(net946));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer488 (.I(\sa21_sr[1] ),
    .Z(net947));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer489 (.I(\sa21_sr[7] ),
    .Z(net948));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer490 (.I(_14414_),
    .Z(net949));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer491 (.I(net949),
    .Z(net950));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer492 (.I(_14414_),
    .Z(net951));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer493 (.I(net951),
    .Z(net952));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold494 (.I(net216),
    .Z(net953));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer5 (.I(net1115),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer6 (.I(net588),
    .Z(net479));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer7 (.I(_15650_),
    .Z(net480));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer8 (.I(net480),
    .Z(net481));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer9 (.I(_15650_),
    .Z(net482));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer10 (.I(_15897_),
    .Z(net483));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer11 (.I(net483),
    .Z(net484));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer12 (.I(_15897_),
    .Z(net485));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer13 (.I(net968),
    .Z(net486));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer14 (.I(net486),
    .Z(net487));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer15 (.I(\u0.w[2][24] ),
    .Z(net488));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer16 (.I(net488),
    .Z(net489));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer17 (.I(net489),
    .Z(net490));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer18 (.I(\sa10_sub[0] ),
    .Z(net491));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer19 (.I(\sa10_sr[1] ),
    .Z(net492));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer20 (.I(\sa10_sr[1] ),
    .Z(net493));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer21 (.I(_15929_),
    .Z(net494));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer22 (.I(net557),
    .Z(net495));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer23 (.I(net1269),
    .Z(net496));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer24 (.I(net1269),
    .Z(net497));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer25 (.I(_01057_),
    .Z(net498));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer26 (.I(net1269),
    .Z(net499));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer27 (.I(_15903_),
    .Z(net500));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer28 (.I(net500),
    .Z(net501));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer29 (.I(net1270),
    .Z(net502));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer30 (.I(net1270),
    .Z(net527));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer31 (.I(\sa21_sub[1] ),
    .Z(net528));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer32 (.I(\sa21_sub[1] ),
    .Z(net529));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer33 (.I(net529),
    .Z(net530));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer34 (.I(\sa03_sr[1] ),
    .Z(net531));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer35 (.I(\sa21_sub[0] ),
    .Z(net532));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer36 (.I(net918),
    .Z(net533));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer37 (.I(_07466_),
    .Z(net534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer38 (.I(_15906_),
    .Z(net535));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer39 (.I(_15906_),
    .Z(net536));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer40 (.I(net536),
    .Z(net537));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer47 (.I(_15778_),
    .Z(net538));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer48 (.I(net538),
    .Z(net539));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer49 (.I(net542),
    .Z(net540));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer50 (.I(net542),
    .Z(net541));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer68 (.I(_15778_),
    .Z(net542));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer69 (.I(_15866_),
    .Z(net543));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer70 (.I(_15866_),
    .Z(net544));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer71 (.I(_15866_),
    .Z(net545));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer72 (.I(net545),
    .Z(net546));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer73 (.I(_15802_),
    .Z(net547));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer74 (.I(_15203_),
    .Z(net548));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer75 (.I(_15769_),
    .Z(net549));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer76 (.I(net549),
    .Z(net550));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer77 (.I(_15769_),
    .Z(net556));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer78 (.I(_15929_),
    .Z(net557));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer100 (.I(net865),
    .Z(net586));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer101 (.I(net586),
    .Z(net587));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone102 (.A1(_01574_),
    .A2(_01579_),
    .ZN(net588));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer103 (.I(_01993_),
    .Z(net589));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer104 (.I(_01993_),
    .Z(net590));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer105 (.I(\sa30_sr[0] ),
    .Z(net617));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer106 (.I(\sa00_sr[1] ),
    .Z(net618));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer107 (.I(net618),
    .Z(net619));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer108 (.I(\sa00_sr[1] ),
    .Z(net620));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer109 (.I(_15932_),
    .Z(net621));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer110 (.I(\u0.w[2][25] ),
    .Z(net622));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer111 (.I(net622),
    .Z(net623));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer112 (.I(_09752_),
    .Z(net624));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer113 (.I(_15640_),
    .Z(net625));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer126 (.I(\u0.tmp_w[25] ),
    .Z(net626));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer127 (.I(net626),
    .Z(net627));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer128 (.I(net626),
    .Z(net628));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer129 (.I(\u0.w[0][25] ),
    .Z(net629));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer130 (.I(\u0.w[0][25] ),
    .Z(net630));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer131 (.I(net630),
    .Z(net631));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer158 (.I(\u0.w[1][25] ),
    .Z(net652));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer159 (.I(net652),
    .Z(net653));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer160 (.I(net652),
    .Z(net654));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer161 (.I(net654),
    .Z(net655));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer162 (.I(\u0.w[1][24] ),
    .Z(net696));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer163 (.I(\u0.w[1][24] ),
    .Z(net697));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer164 (.I(net697),
    .Z(net698));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer165 (.I(net698),
    .Z(net699));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer166 (.I(net699),
    .Z(net700));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer167 (.I(_07697_),
    .Z(net706));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer168 (.I(_07697_),
    .Z(net707));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer169 (.I(_07674_),
    .Z(net708));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer170 (.I(\u0.w[2][26] ),
    .Z(net709));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer171 (.I(_07682_),
    .Z(net710));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer172 (.I(_15642_),
    .Z(net711));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer186 (.I(net962),
    .Z(net757));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer187 (.I(net757),
    .Z(net758));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer193 (.I(net962),
    .Z(net759));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer194 (.I(_09753_),
    .Z(net760));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer195 (.I(_09809_),
    .Z(net761));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer196 (.I(_15639_),
    .Z(net762));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer237 (.I(net762),
    .Z(net763));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer238 (.I(_07679_),
    .Z(net764));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer239 (.I(_09779_),
    .Z(net765));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer240 (.I(\u0.w[1][26] ),
    .Z(net766));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer241 (.I(net766),
    .Z(net767));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer243 (.I(net767),
    .Z(net768));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer244 (.I(_15775_),
    .Z(net769));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer245 (.I(_15775_),
    .Z(net770));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer247 (.I(_12801_),
    .Z(net771));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer248 (.I(\sa10_sub[7] ),
    .Z(net772));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer249 (.I(_12998_),
    .Z(net773));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer250 (.I(_15772_),
    .Z(net774));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer251 (.I(_13034_),
    .Z(net775));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone252 (.I(_12912_),
    .Z(net776));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer298 (.I(\sa21_sub[1] ),
    .Z(net777));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer299 (.I(_12768_),
    .Z(net778));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer300 (.I(_12801_),
    .Z(net779));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer301 (.I(_12917_),
    .Z(net780));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer312 (.I(_09912_),
    .Z(net822));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer313 (.I(net822),
    .Z(net823));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer314 (.I(_07706_),
    .Z(net824));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer315 (.I(_07706_),
    .Z(net825));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer316 (.I(_09734_),
    .Z(net832));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer317 (.I(net832),
    .Z(net833));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer318 (.I(net832),
    .Z(net838));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer319 (.I(net838),
    .Z(net839));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer320 (.I(_09842_),
    .Z(net840));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer321 (.I(_15708_),
    .Z(net841));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer322 (.I(_15705_),
    .Z(net842));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer323 (.I(net842),
    .Z(net843));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer324 (.I(net843),
    .Z(net844));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer325 (.I(_15705_),
    .Z(net845));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer366 (.I(_01614_),
    .Z(net857));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer373 (.I(net857),
    .Z(net858));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer374 (.I(\sa10_sr[2] ),
    .Z(net859));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer379 (.I(\sa10_sr[2] ),
    .Z(net860));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer380 (.I(\sa10_sr[2] ),
    .Z(net861));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer381 (.I(_01615_),
    .Z(net862));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer382 (.I(_15940_),
    .Z(net863));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer383 (.I(net863),
    .Z(net864));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer384 (.I(net863),
    .Z(net865));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer385 (.I(_01591_),
    .Z(net885));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 rebuffer386 (.I(_01620_),
    .Z(net886));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer392 (.I(_16175_),
    .Z(net892));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer395 (.I(_15537_),
    .Z(net895));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer396 (.I(_08011_),
    .Z(net896));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer403 (.I(\sa21_sr[1] ),
    .Z(net918));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer404 (.I(_15840_),
    .Z(net919));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer405 (.I(net919),
    .Z(net920));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer429 (.I(_13139_),
    .Z(net926));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer430 (.I(_13139_),
    .Z(net927));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer432 (.I(net4),
    .Z(net929));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer433 (.I(_13403_),
    .Z(net930));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer434 (.I(_12783_),
    .Z(net931));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer435 (.I(_12783_),
    .Z(net932));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer436 (.I(_13174_),
    .Z(net933));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer457 (.I(_00873_),
    .Z(net940));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer458 (.I(_00873_),
    .Z(net941));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer469 (.I(_15645_),
    .Z(net962));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer470 (.I(_12858_),
    .Z(net963));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer471 (.I(_12826_),
    .Z(net964));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer472 (.I(_13000_),
    .Z(net965));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer473 (.I(_12982_),
    .Z(net966));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer474 (.I(_12981_),
    .Z(net967));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer475 (.I(_15770_),
    .Z(net968));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer476 (.I(_12918_),
    .Z(net969));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone477 (.A1(_12861_),
    .A2(net487),
    .ZN(net970));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer478 (.I(_12807_),
    .Z(net971));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer479 (.I(_12996_),
    .Z(net972));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer480 (.I(_13101_),
    .Z(net973));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer481 (.I(_12810_),
    .Z(net974));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer482 (.I(_12809_),
    .Z(net975));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer483 (.I(net975),
    .Z(net976));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer494 (.I(_15712_),
    .Z(net979));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer495 (.I(net1147),
    .Z(net980));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer508 (.I(_00811_),
    .Z(net993));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer526 (.I(_00907_),
    .Z(net1011));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer537 (.I(\sa01_sr[7] ),
    .Z(net1022));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer538 (.I(_15706_),
    .Z(net1023));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer539 (.I(_15706_),
    .Z(net1024));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer543 (.I(_11161_),
    .Z(net1028));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer544 (.I(\sa30_sub[1] ),
    .Z(net1029));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer545 (.I(\u0.w[1][17] ),
    .Z(net1030));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer546 (.I(net1030),
    .Z(net1031));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer547 (.I(net1031),
    .Z(net1032));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer548 (.I(\u0.w[1][17] ),
    .Z(net1033));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer549 (.I(_07987_),
    .Z(net1034));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer550 (.I(\u0.subword[17] ),
    .Z(net1035));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer551 (.I(_15543_),
    .Z(net1036));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer552 (.I(net1036),
    .Z(net1037));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer553 (.I(_15543_),
    .Z(net1038));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer554 (.I(net18),
    .Z(net1039));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone555 (.I(net910),
    .Z(net1040));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer556 (.I(_06902_),
    .Z(net1041));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer557 (.I(_06902_),
    .Z(net1042));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer562 (.I(_15176_),
    .Z(net1047));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer563 (.I(_15865_),
    .Z(net1048));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer564 (.I(_15865_),
    .Z(net1049));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer565 (.I(net1258),
    .Z(net1050));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 clone566 (.A1(net8),
    .A2(_15883_),
    .A3(net1048),
    .ZN(net1051));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer567 (.I(_03963_),
    .Z(net1052));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer568 (.I(net1052),
    .Z(net1053));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer569 (.I(net1052),
    .Z(net1054));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer570 (.I(_03963_),
    .Z(net1055));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer571 (.I(_03973_),
    .Z(net1056));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer572 (.I(_03982_),
    .Z(net1057));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer573 (.I(net1057),
    .Z(net1058));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer574 (.I(net1057),
    .Z(net1059));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer575 (.I(_16046_),
    .Z(net1060));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer580 (.I(_16073_),
    .Z(net1065));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer581 (.I(net1065),
    .Z(net1066));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer582 (.I(\sa00_sr[0] ),
    .Z(net1067));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer583 (.I(_16074_),
    .Z(net1068));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer584 (.I(_04534_),
    .Z(net1069));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer585 (.I(_04655_),
    .Z(net1070));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer586 (.I(_04767_),
    .Z(net1071));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer587 (.I(_04767_),
    .Z(net1072));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer588 (.I(\sa20_sr[0] ),
    .Z(net1073));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone589 (.I(_04574_),
    .Z(net1074));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer590 (.I(_04571_),
    .Z(net1075));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone591 (.I(_04574_),
    .Z(net1076));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer592 (.I(_04656_),
    .Z(net1077));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer593 (.I(\sa30_sr[1] ),
    .Z(net1078));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer594 (.I(\sa30_sr[1] ),
    .Z(net1079));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer595 (.I(_04568_),
    .Z(net1080));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer596 (.I(_04594_),
    .Z(net1081));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer597 (.I(_04595_),
    .Z(net1082));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer598 (.I(_04662_),
    .Z(net1083));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer599 (.I(_04630_),
    .Z(net1084));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer600 (.I(_01588_),
    .Z(net1085));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer603 (.I(_15898_),
    .Z(net1088));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer604 (.I(_15898_),
    .Z(net1089));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer605 (.I(_00876_),
    .Z(net1090));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer606 (.I(net1090),
    .Z(net1091));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone607 (.I(net1093),
    .Z(net1092));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer608 (.I(_00946_),
    .Z(net1093));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone609 (.I(_00946_),
    .Z(net1094));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer610 (.I(_01064_),
    .Z(net1095));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer611 (.I(_01064_),
    .Z(net1096));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer612 (.I(_00906_),
    .Z(net1097));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer613 (.I(_05302_),
    .Z(net1098));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer628 (.I(_01790_),
    .Z(net1113));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer629 (.I(_01722_),
    .Z(net1114));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer630 (.I(_15935_),
    .Z(net1115));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer631 (.I(_15935_),
    .Z(net1116));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer632 (.I(_01562_),
    .Z(net1117));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer633 (.I(_15930_),
    .Z(net1118));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer634 (.I(_01596_),
    .Z(net1119));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer635 (.I(net27),
    .Z(net1120));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer636 (.I(_16105_),
    .Z(net1121));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer637 (.I(net1121),
    .Z(net1122));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer638 (.I(_16108_),
    .Z(net1123));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer647 (.I(_13796_),
    .Z(net1132));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer648 (.I(_13782_),
    .Z(net1133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer649 (.I(_13718_),
    .Z(net1134));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer650 (.I(_13602_),
    .Z(net1135));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer651 (.I(_15807_),
    .Z(net1136));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone652 (.I(_01725_),
    .Z(net1137));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer653 (.I(_13583_),
    .Z(net1138));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer654 (.I(_01743_),
    .Z(net1139));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer657 (.I(_16079_),
    .Z(net1142));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer658 (.I(_16079_),
    .Z(net1143));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer659 (.I(_04724_),
    .Z(net1144));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer661 (.I(_11147_),
    .Z(net1146));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer662 (.I(_11186_),
    .Z(net1147));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer664 (.I(_12138_),
    .Z(net1149));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 rebuffer665 (.I(_15746_),
    .Z(net1150));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer666 (.I(net1150),
    .Z(net1151));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer667 (.I(_11997_),
    .Z(net1152));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer668 (.I(_11997_),
    .Z(net1153));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer669 (.I(net1153),
    .Z(net1154));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 clone670 (.A1(_15755_),
    .A2(net71),
    .A3(net20),
    .ZN(net1155));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer671 (.I(_15737_),
    .Z(net1156));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer672 (.I(\sa12_sr[7] ),
    .Z(net1157));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer673 (.I(_12225_),
    .Z(net1158));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer674 (.I(_15744_),
    .Z(net1159));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer675 (.I(_15744_),
    .Z(net1160));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer676 (.I(_15740_),
    .Z(net1161));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer677 (.I(_15738_),
    .Z(net1162));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer678 (.I(_12279_),
    .Z(net1163));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer679 (.I(_12279_),
    .Z(net1164));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer680 (.I(\sa12_sr[7] ),
    .Z(net1165));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer681 (.I(_11991_),
    .Z(net1166));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer682 (.I(_11960_),
    .Z(net1167));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer683 (.I(_11960_),
    .Z(net1168));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer684 (.I(\sa20_sub[1] ),
    .Z(net1169));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer685 (.I(\sa20_sub[1] ),
    .Z(net1170));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer686 (.I(_12132_),
    .Z(net1171));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer687 (.I(\sa02_sr[7] ),
    .Z(net1172));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer688 (.I(net1172),
    .Z(net1173));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer689 (.I(_12000_),
    .Z(net1174));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer690 (.I(_11963_),
    .Z(net1175));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer691 (.I(\sa02_sr[0] ),
    .Z(net1176));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer692 (.I(\sa02_sr[0] ),
    .Z(net1177));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer693 (.I(\sa12_sr[0] ),
    .Z(net1178));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer694 (.I(\sa12_sr[0] ),
    .Z(net1179));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split695 (.I(\sa12_sr[0] ),
    .Z(net1180));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer696 (.I(_06024_),
    .Z(net1181));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer697 (.I(_05987_),
    .Z(net1182));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer698 (.I(net1182),
    .Z(net1183));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer699 (.I(_16137_),
    .Z(net1184));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer700 (.I(net1184),
    .Z(net1185));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer701 (.I(_06123_),
    .Z(net1186));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer702 (.I(net1207),
    .Z(net1187));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer703 (.I(_16137_),
    .Z(net1188));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer704 (.I(_16146_),
    .Z(net1189));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer705 (.I(\sa12_sr[1] ),
    .Z(net1190));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer706 (.I(_06053_),
    .Z(net1191));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer707 (.I(_03026_),
    .Z(net1192));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer708 (.I(_06025_),
    .Z(net1193));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer709 (.I(_06000_),
    .Z(net1194));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer710 (.I(_06116_),
    .Z(net1195));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer711 (.I(net1195),
    .Z(net1196));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer712 (.I(_06303_),
    .Z(net1197));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer713 (.I(\sa02_sr[1] ),
    .Z(net1198));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer714 (.I(_06050_),
    .Z(net1199));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer715 (.I(_06050_),
    .Z(net1200));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone716 (.I(_06090_),
    .Z(net1201));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer717 (.I(_16143_),
    .Z(net1202));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer720 (.I(_16144_),
    .Z(net1205));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 rebuffer721 (.I(_06031_),
    .Z(net1206));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer722 (.I(_16144_),
    .Z(net1207));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer723 (.I(_16144_),
    .Z(net1208));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone724 (.I(_06071_),
    .Z(net1209));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer725 (.I(_16138_),
    .Z(net1210));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer726 (.I(_05994_),
    .Z(net1211));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer727 (.I(_01646_),
    .Z(net1212));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer728 (.I(_01646_),
    .Z(net1213));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer729 (.I(net1213),
    .Z(net1214));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer730 (.I(_01730_),
    .Z(net1215));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 rebuffer731 (.I(_01643_),
    .Z(net1216));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer732 (.I(_15874_),
    .Z(net1217));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer733 (.I(net1217),
    .Z(net1218));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer734 (.I(net1217),
    .Z(net1219));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer735 (.I(net1217),
    .Z(net1220));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer736 (.I(net1220),
    .Z(net1221));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer737 (.I(_00868_),
    .Z(net1222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer738 (.I(_00906_),
    .Z(net1223));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer739 (.I(_00877_),
    .Z(net1224));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer740 (.I(net1224),
    .Z(net1225));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer741 (.I(_00872_),
    .Z(net1226));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer742 (.I(_00807_),
    .Z(net1227));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer743 (.I(net1234),
    .Z(net1228));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone744 (.A1(net21),
    .A2(_00909_),
    .ZN(net1229));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer745 (.I(_01070_),
    .Z(net1230));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer746 (.I(_15904_),
    .Z(net1231));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer747 (.I(_15904_),
    .Z(net1232));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer748 (.I(_01109_),
    .Z(net1233));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer749 (.I(_01071_),
    .Z(net1234));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer754 (.I(_11215_),
    .Z(net1239));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer755 (.I(_05297_),
    .Z(net1240));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer756 (.I(net1240),
    .Z(net1241));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer773 (.I(_15865_),
    .Z(net1258));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer774 (.I(_15679_),
    .Z(net1259));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer775 (.I(_15679_),
    .Z(net1260));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer776 (.I(_10664_),
    .Z(net1261));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer777 (.I(net36),
    .Z(net1262));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer778 (.I(net36),
    .Z(net1263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer779 (.I(net1263),
    .Z(net1264));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer781 (.I(_01106_),
    .Z(net1266));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer782 (.I(_01106_),
    .Z(net1267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer783 (.I(_00827_),
    .Z(net1268));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer784 (.I(_15903_),
    .Z(net1269));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer785 (.I(_00825_),
    .Z(net1270));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer786 (.I(_00995_),
    .Z(net1271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer788 (.I(_15833_),
    .Z(net1273));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net216));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_241_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_241_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_241_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2220 ();
endmodule
