module skid_buffer (clk,
    m_ready,
    m_valid,
    rst_n,
    s_ready,
    s_valid,
    m_data,
    s_data);
 input clk;
 input m_ready;
 output m_valid;
 input rst_n;
 output s_ready;
 input s_valid;
 output [7:0] m_data;
 input [7:0] s_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire \skid_reg[0] ;
 wire \skid_reg[1] ;
 wire \skid_reg[2] ;
 wire \skid_reg[3] ;
 wire \skid_reg[4] ;
 wire \skid_reg[5] ;
 wire \skid_reg[6] ;
 wire \skid_reg[7] ;
 wire skid_valid_reg;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X4 _087_ (.A(net18),
    .Z(_030_));
 CLKBUF_X3 _088_ (.A(_030_),
    .Z(_031_));
 CLKBUF_X3 _089_ (.A(m_ready),
    .Z(_032_));
 CLKBUF_X3 _090_ (.A(_032_),
    .Z(_033_));
 AOI21_X1 _091_ (.A(_000_),
    .B1(_031_),
    .B2(_033_),
    .ZN(_034_));
 INV_X1 _092_ (.A(_034_),
    .ZN(net19));
 BUF_X2 _093_ (.A(rst_n),
    .Z(_035_));
 BUF_X4 _094_ (.A(skid_valid_reg),
    .Z(_036_));
 NAND3_X4 _095_ (.A1(_032_),
    .A2(_030_),
    .A3(_036_),
    .ZN(_037_));
 MUX2_X1 _096_ (.A(\skid_reg[0] ),
    .B(net1),
    .S(_037_),
    .Z(_038_));
 MUX2_X1 _097_ (.A(_030_),
    .B(net9),
    .S(_000_),
    .Z(_039_));
 INV_X2 _098_ (.A(_030_),
    .ZN(_040_));
 OAI21_X4 _099_ (.A(_039_),
    .B1(_040_),
    .B2(_032_),
    .ZN(_041_));
 BUF_X8 _100_ (.A(_041_),
    .Z(_042_));
 MUX2_X1 _101_ (.A(_038_),
    .B(net10),
    .S(_042_),
    .Z(_043_));
 AND2_X1 _102_ (.A1(_035_),
    .A2(_043_),
    .ZN(_001_));
 INV_X2 _103_ (.A(_035_),
    .ZN(_044_));
 NAND4_X1 _104_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[1] ),
    .ZN(_045_));
 AOI21_X1 _105_ (.A(_042_),
    .B1(_037_),
    .B2(net2),
    .ZN(_046_));
 INV_X1 _106_ (.A(net11),
    .ZN(_047_));
 AOI221_X1 _107_ (.A(_044_),
    .B1(_045_),
    .B2(_046_),
    .C1(_042_),
    .C2(_047_),
    .ZN(_002_));
 NAND4_X1 _108_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[2] ),
    .ZN(_048_));
 AOI21_X1 _109_ (.A(_042_),
    .B1(_037_),
    .B2(net3),
    .ZN(_049_));
 INV_X1 _110_ (.A(net12),
    .ZN(_050_));
 AOI221_X1 _111_ (.A(_044_),
    .B1(_048_),
    .B2(_049_),
    .C1(_042_),
    .C2(_050_),
    .ZN(_003_));
 NAND4_X1 _112_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[3] ),
    .ZN(_051_));
 AOI21_X1 _113_ (.A(_041_),
    .B1(_037_),
    .B2(net4),
    .ZN(_052_));
 INV_X1 _114_ (.A(net13),
    .ZN(_053_));
 AOI221_X1 _115_ (.A(_044_),
    .B1(_051_),
    .B2(_052_),
    .C1(_042_),
    .C2(_053_),
    .ZN(_004_));
 NAND4_X1 _116_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[4] ),
    .ZN(_054_));
 AOI21_X1 _117_ (.A(_041_),
    .B1(_037_),
    .B2(net5),
    .ZN(_055_));
 INV_X1 _118_ (.A(net14),
    .ZN(_056_));
 AOI221_X1 _119_ (.A(_044_),
    .B1(_054_),
    .B2(_055_),
    .C1(_042_),
    .C2(_056_),
    .ZN(_005_));
 NAND4_X1 _120_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[5] ),
    .ZN(_057_));
 AOI21_X1 _121_ (.A(_041_),
    .B1(_037_),
    .B2(net6),
    .ZN(_058_));
 INV_X1 _122_ (.A(net15),
    .ZN(_059_));
 AOI221_X1 _123_ (.A(_044_),
    .B1(_057_),
    .B2(_058_),
    .C1(_042_),
    .C2(_059_),
    .ZN(_006_));
 NAND4_X1 _124_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[6] ),
    .ZN(_060_));
 AOI21_X1 _125_ (.A(_041_),
    .B1(_037_),
    .B2(net7),
    .ZN(_061_));
 INV_X1 _126_ (.A(net16),
    .ZN(_062_));
 AOI221_X1 _127_ (.A(_044_),
    .B1(_060_),
    .B2(_061_),
    .C1(_042_),
    .C2(_062_),
    .ZN(_007_));
 NAND4_X1 _128_ (.A1(_033_),
    .A2(_031_),
    .A3(_036_),
    .A4(\skid_reg[7] ),
    .ZN(_063_));
 AOI21_X1 _129_ (.A(_041_),
    .B1(_037_),
    .B2(net8),
    .ZN(_064_));
 INV_X1 _130_ (.A(net17),
    .ZN(_065_));
 AOI221_X1 _131_ (.A(_044_),
    .B1(_063_),
    .B2(_064_),
    .C1(_042_),
    .C2(_065_),
    .ZN(_008_));
 NAND2_X1 _132_ (.A1(net9),
    .A2(_000_),
    .ZN(_066_));
 NOR3_X4 _133_ (.A1(_032_),
    .A2(_040_),
    .A3(_066_),
    .ZN(_067_));
 MUX2_X1 _134_ (.A(\skid_reg[0] ),
    .B(net1),
    .S(_067_),
    .Z(_068_));
 AND2_X1 _135_ (.A1(_035_),
    .A2(_068_),
    .ZN(_009_));
 MUX2_X1 _136_ (.A(\skid_reg[1] ),
    .B(net2),
    .S(_067_),
    .Z(_069_));
 AND2_X1 _137_ (.A1(_035_),
    .A2(_069_),
    .ZN(_010_));
 MUX2_X1 _138_ (.A(\skid_reg[2] ),
    .B(net3),
    .S(_067_),
    .Z(_019_));
 AND2_X1 _139_ (.A1(_035_),
    .A2(_019_),
    .ZN(_011_));
 MUX2_X1 _140_ (.A(\skid_reg[3] ),
    .B(net4),
    .S(_067_),
    .Z(_020_));
 AND2_X1 _141_ (.A1(_035_),
    .A2(_020_),
    .ZN(_012_));
 MUX2_X1 _142_ (.A(\skid_reg[4] ),
    .B(net5),
    .S(_067_),
    .Z(_021_));
 AND2_X1 _143_ (.A1(_035_),
    .A2(_021_),
    .ZN(_013_));
 MUX2_X1 _144_ (.A(\skid_reg[5] ),
    .B(net6),
    .S(_067_),
    .Z(_022_));
 AND2_X1 _145_ (.A1(_035_),
    .A2(_022_),
    .ZN(_014_));
 MUX2_X1 _146_ (.A(\skid_reg[6] ),
    .B(net7),
    .S(_067_),
    .Z(_023_));
 AND2_X1 _147_ (.A1(_035_),
    .A2(_023_),
    .ZN(_015_));
 MUX2_X1 _148_ (.A(\skid_reg[7] ),
    .B(net8),
    .S(_067_),
    .Z(_024_));
 AND2_X1 _149_ (.A1(_035_),
    .A2(_024_),
    .ZN(_016_));
 NAND2_X1 _150_ (.A1(_033_),
    .A2(_031_),
    .ZN(_025_));
 AOI21_X1 _151_ (.A(_067_),
    .B1(_025_),
    .B2(_036_),
    .ZN(_026_));
 NOR2_X1 _152_ (.A1(_044_),
    .A2(_026_),
    .ZN(_017_));
 INV_X1 _153_ (.A(net9),
    .ZN(_027_));
 NAND2_X1 _154_ (.A1(_033_),
    .A2(_027_),
    .ZN(_028_));
 OAI21_X1 _155_ (.A(_031_),
    .B1(_036_),
    .B2(_028_),
    .ZN(_029_));
 AOI21_X1 _156_ (.A(_044_),
    .B1(_066_),
    .B2(_029_),
    .ZN(_018_));
 DFF_X2 \data_reg[0]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net10),
    .QN(_086_));
 DFF_X2 \data_reg[1]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net11),
    .QN(_085_));
 DFF_X2 \data_reg[2]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net12),
    .QN(_084_));
 DFF_X2 \data_reg[3]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_083_));
 DFF_X2 \data_reg[4]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net14),
    .QN(_082_));
 DFF_X2 \data_reg[5]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net15),
    .QN(_081_));
 DFF_X2 \data_reg[6]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_080_));
 DFF_X2 \data_reg[7]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_079_));
 DFF_X1 \skid_reg[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\skid_reg[0] ),
    .QN(_078_));
 DFF_X1 \skid_reg[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\skid_reg[1] ),
    .QN(_077_));
 DFF_X1 \skid_reg[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\skid_reg[2] ),
    .QN(_076_));
 DFF_X1 \skid_reg[3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\skid_reg[3] ),
    .QN(_075_));
 DFF_X1 \skid_reg[4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\skid_reg[4] ),
    .QN(_074_));
 DFF_X1 \skid_reg[5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\skid_reg[5] ),
    .QN(_073_));
 DFF_X1 \skid_reg[6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\skid_reg[6] ),
    .QN(_072_));
 DFF_X1 \skid_reg[7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\skid_reg[7] ),
    .QN(_071_));
 DFF_X1 \skid_valid_reg$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_1_0__leaf_clk),
    .Q(skid_valid_reg),
    .QN(_000_));
 DFF_X2 \valid_reg$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net18),
    .QN(_070_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_292 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_293 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_294 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_295 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_296 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_297 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_298 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_299 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_300 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_301 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_302 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_303 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_304 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_305 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_306 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_307 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_308 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_330 ();
 BUF_X1 input1 (.A(s_data[0]),
    .Z(net1));
 CLKBUF_X2 input2 (.A(s_data[1]),
    .Z(net2));
 BUF_X1 input3 (.A(s_data[2]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(s_data[3]),
    .Z(net4));
 CLKBUF_X2 input5 (.A(s_data[4]),
    .Z(net5));
 CLKBUF_X2 input6 (.A(s_data[5]),
    .Z(net6));
 CLKBUF_X2 input7 (.A(s_data[6]),
    .Z(net7));
 CLKBUF_X2 input8 (.A(s_data[7]),
    .Z(net8));
 CLKBUF_X2 input9 (.A(s_valid),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(m_data[0]));
 BUF_X1 output11 (.A(net11),
    .Z(m_data[1]));
 BUF_X1 output12 (.A(net12),
    .Z(m_data[2]));
 BUF_X1 output13 (.A(net13),
    .Z(m_data[3]));
 BUF_X1 output14 (.A(net14),
    .Z(m_data[4]));
 BUF_X1 output15 (.A(net15),
    .Z(m_data[5]));
 BUF_X1 output16 (.A(net16),
    .Z(m_data[6]));
 BUF_X1 output17 (.A(net17),
    .Z(m_data[7]));
 BUF_X1 output18 (.A(net18),
    .Z(m_valid));
 BUF_X1 output19 (.A(net19),
    .Z(s_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X8 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_464 ();
 FILLCELL_X32 FILLER_0_496 ();
 FILLCELL_X32 FILLER_0_528 ();
 FILLCELL_X32 FILLER_0_560 ();
 FILLCELL_X32 FILLER_0_592 ();
 FILLCELL_X4 FILLER_0_624 ();
 FILLCELL_X2 FILLER_0_628 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X32 FILLER_0_856 ();
 FILLCELL_X32 FILLER_0_888 ();
 FILLCELL_X32 FILLER_0_920 ();
 FILLCELL_X16 FILLER_0_952 ();
 FILLCELL_X8 FILLER_0_968 ();
 FILLCELL_X2 FILLER_0_976 ();
 FILLCELL_X1 FILLER_0_978 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X16 FILLER_1_449 ();
 FILLCELL_X8 FILLER_1_465 ();
 FILLCELL_X2 FILLER_1_473 ();
 FILLCELL_X1 FILLER_1_475 ();
 FILLCELL_X32 FILLER_1_480 ();
 FILLCELL_X32 FILLER_1_512 ();
 FILLCELL_X32 FILLER_1_544 ();
 FILLCELL_X32 FILLER_1_576 ();
 FILLCELL_X32 FILLER_1_608 ();
 FILLCELL_X32 FILLER_1_640 ();
 FILLCELL_X32 FILLER_1_672 ();
 FILLCELL_X32 FILLER_1_704 ();
 FILLCELL_X32 FILLER_1_736 ();
 FILLCELL_X32 FILLER_1_768 ();
 FILLCELL_X32 FILLER_1_800 ();
 FILLCELL_X32 FILLER_1_832 ();
 FILLCELL_X32 FILLER_1_864 ();
 FILLCELL_X32 FILLER_1_896 ();
 FILLCELL_X32 FILLER_1_928 ();
 FILLCELL_X16 FILLER_1_960 ();
 FILLCELL_X2 FILLER_1_976 ();
 FILLCELL_X1 FILLER_1_978 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X16 FILLER_2_952 ();
 FILLCELL_X8 FILLER_2_968 ();
 FILLCELL_X2 FILLER_2_976 ();
 FILLCELL_X1 FILLER_2_978 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X16 FILLER_3_961 ();
 FILLCELL_X2 FILLER_3_977 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X16 FILLER_4_952 ();
 FILLCELL_X8 FILLER_4_968 ();
 FILLCELL_X2 FILLER_4_976 ();
 FILLCELL_X1 FILLER_4_978 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X16 FILLER_5_961 ();
 FILLCELL_X2 FILLER_5_977 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X16 FILLER_6_952 ();
 FILLCELL_X8 FILLER_6_968 ();
 FILLCELL_X2 FILLER_6_976 ();
 FILLCELL_X1 FILLER_6_978 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X16 FILLER_7_961 ();
 FILLCELL_X2 FILLER_7_977 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X16 FILLER_8_952 ();
 FILLCELL_X8 FILLER_8_968 ();
 FILLCELL_X2 FILLER_8_976 ();
 FILLCELL_X1 FILLER_8_978 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X16 FILLER_9_961 ();
 FILLCELL_X2 FILLER_9_977 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X16 FILLER_10_952 ();
 FILLCELL_X8 FILLER_10_968 ();
 FILLCELL_X2 FILLER_10_976 ();
 FILLCELL_X1 FILLER_10_978 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X16 FILLER_11_961 ();
 FILLCELL_X2 FILLER_11_977 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X16 FILLER_12_952 ();
 FILLCELL_X8 FILLER_12_968 ();
 FILLCELL_X2 FILLER_12_976 ();
 FILLCELL_X1 FILLER_12_978 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X16 FILLER_13_961 ();
 FILLCELL_X2 FILLER_13_977 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X16 FILLER_14_952 ();
 FILLCELL_X8 FILLER_14_968 ();
 FILLCELL_X2 FILLER_14_976 ();
 FILLCELL_X1 FILLER_14_978 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X16 FILLER_15_961 ();
 FILLCELL_X2 FILLER_15_977 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X16 FILLER_16_952 ();
 FILLCELL_X8 FILLER_16_968 ();
 FILLCELL_X2 FILLER_16_976 ();
 FILLCELL_X1 FILLER_16_978 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X16 FILLER_17_961 ();
 FILLCELL_X2 FILLER_17_977 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X16 FILLER_18_952 ();
 FILLCELL_X8 FILLER_18_968 ();
 FILLCELL_X2 FILLER_18_976 ();
 FILLCELL_X1 FILLER_18_978 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X16 FILLER_19_961 ();
 FILLCELL_X2 FILLER_19_977 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X16 FILLER_20_952 ();
 FILLCELL_X8 FILLER_20_968 ();
 FILLCELL_X2 FILLER_20_976 ();
 FILLCELL_X1 FILLER_20_978 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X16 FILLER_21_961 ();
 FILLCELL_X2 FILLER_21_977 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X16 FILLER_22_952 ();
 FILLCELL_X8 FILLER_22_968 ();
 FILLCELL_X2 FILLER_22_976 ();
 FILLCELL_X1 FILLER_22_978 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X16 FILLER_23_961 ();
 FILLCELL_X2 FILLER_23_977 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X16 FILLER_24_952 ();
 FILLCELL_X8 FILLER_24_968 ();
 FILLCELL_X2 FILLER_24_976 ();
 FILLCELL_X1 FILLER_24_978 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X16 FILLER_25_961 ();
 FILLCELL_X2 FILLER_25_977 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X16 FILLER_26_952 ();
 FILLCELL_X8 FILLER_26_968 ();
 FILLCELL_X2 FILLER_26_976 ();
 FILLCELL_X1 FILLER_26_978 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X16 FILLER_27_961 ();
 FILLCELL_X2 FILLER_27_977 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X16 FILLER_28_952 ();
 FILLCELL_X8 FILLER_28_968 ();
 FILLCELL_X2 FILLER_28_976 ();
 FILLCELL_X1 FILLER_28_978 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X16 FILLER_29_961 ();
 FILLCELL_X2 FILLER_29_977 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X16 FILLER_30_952 ();
 FILLCELL_X8 FILLER_30_968 ();
 FILLCELL_X2 FILLER_30_976 ();
 FILLCELL_X1 FILLER_30_978 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X16 FILLER_31_961 ();
 FILLCELL_X2 FILLER_31_977 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X16 FILLER_32_952 ();
 FILLCELL_X8 FILLER_32_968 ();
 FILLCELL_X2 FILLER_32_976 ();
 FILLCELL_X1 FILLER_32_978 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X16 FILLER_33_961 ();
 FILLCELL_X2 FILLER_33_977 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X16 FILLER_34_952 ();
 FILLCELL_X8 FILLER_34_968 ();
 FILLCELL_X2 FILLER_34_976 ();
 FILLCELL_X1 FILLER_34_978 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X16 FILLER_35_961 ();
 FILLCELL_X2 FILLER_35_977 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X16 FILLER_36_952 ();
 FILLCELL_X8 FILLER_36_968 ();
 FILLCELL_X2 FILLER_36_976 ();
 FILLCELL_X1 FILLER_36_978 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X16 FILLER_37_961 ();
 FILLCELL_X2 FILLER_37_977 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X16 FILLER_38_952 ();
 FILLCELL_X8 FILLER_38_968 ();
 FILLCELL_X2 FILLER_38_976 ();
 FILLCELL_X1 FILLER_38_978 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X16 FILLER_39_961 ();
 FILLCELL_X2 FILLER_39_977 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X16 FILLER_40_952 ();
 FILLCELL_X8 FILLER_40_968 ();
 FILLCELL_X2 FILLER_40_976 ();
 FILLCELL_X1 FILLER_40_978 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X16 FILLER_41_961 ();
 FILLCELL_X2 FILLER_41_977 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X16 FILLER_42_952 ();
 FILLCELL_X8 FILLER_42_968 ();
 FILLCELL_X2 FILLER_42_976 ();
 FILLCELL_X1 FILLER_42_978 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X16 FILLER_43_961 ();
 FILLCELL_X2 FILLER_43_977 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X16 FILLER_44_952 ();
 FILLCELL_X8 FILLER_44_968 ();
 FILLCELL_X2 FILLER_44_976 ();
 FILLCELL_X1 FILLER_44_978 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X16 FILLER_45_961 ();
 FILLCELL_X2 FILLER_45_977 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X16 FILLER_46_952 ();
 FILLCELL_X8 FILLER_46_968 ();
 FILLCELL_X2 FILLER_46_976 ();
 FILLCELL_X1 FILLER_46_978 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X16 FILLER_47_961 ();
 FILLCELL_X2 FILLER_47_977 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X16 FILLER_48_952 ();
 FILLCELL_X8 FILLER_48_968 ();
 FILLCELL_X2 FILLER_48_976 ();
 FILLCELL_X1 FILLER_48_978 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X16 FILLER_49_961 ();
 FILLCELL_X2 FILLER_49_977 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X16 FILLER_50_952 ();
 FILLCELL_X8 FILLER_50_968 ();
 FILLCELL_X2 FILLER_50_976 ();
 FILLCELL_X1 FILLER_50_978 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X16 FILLER_51_961 ();
 FILLCELL_X2 FILLER_51_977 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X16 FILLER_52_952 ();
 FILLCELL_X8 FILLER_52_968 ();
 FILLCELL_X2 FILLER_52_976 ();
 FILLCELL_X1 FILLER_52_978 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X16 FILLER_53_961 ();
 FILLCELL_X2 FILLER_53_977 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X16 FILLER_54_952 ();
 FILLCELL_X8 FILLER_54_968 ();
 FILLCELL_X2 FILLER_54_976 ();
 FILLCELL_X1 FILLER_54_978 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X16 FILLER_55_961 ();
 FILLCELL_X2 FILLER_55_977 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X16 FILLER_56_513 ();
 FILLCELL_X8 FILLER_56_529 ();
 FILLCELL_X1 FILLER_56_537 ();
 FILLCELL_X32 FILLER_56_543 ();
 FILLCELL_X32 FILLER_56_575 ();
 FILLCELL_X16 FILLER_56_607 ();
 FILLCELL_X8 FILLER_56_623 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X16 FILLER_56_952 ();
 FILLCELL_X8 FILLER_56_968 ();
 FILLCELL_X2 FILLER_56_976 ();
 FILLCELL_X1 FILLER_56_978 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X8 FILLER_57_513 ();
 FILLCELL_X2 FILLER_57_521 ();
 FILLCELL_X1 FILLER_57_523 ();
 FILLCELL_X4 FILLER_57_540 ();
 FILLCELL_X1 FILLER_57_544 ();
 FILLCELL_X32 FILLER_57_552 ();
 FILLCELL_X32 FILLER_57_584 ();
 FILLCELL_X32 FILLER_57_616 ();
 FILLCELL_X32 FILLER_57_648 ();
 FILLCELL_X32 FILLER_57_680 ();
 FILLCELL_X32 FILLER_57_712 ();
 FILLCELL_X32 FILLER_57_744 ();
 FILLCELL_X32 FILLER_57_776 ();
 FILLCELL_X32 FILLER_57_808 ();
 FILLCELL_X32 FILLER_57_840 ();
 FILLCELL_X32 FILLER_57_872 ();
 FILLCELL_X32 FILLER_57_904 ();
 FILLCELL_X4 FILLER_57_936 ();
 FILLCELL_X32 FILLER_57_944 ();
 FILLCELL_X2 FILLER_57_976 ();
 FILLCELL_X1 FILLER_57_978 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X16 FILLER_58_513 ();
 FILLCELL_X2 FILLER_58_529 ();
 FILLCELL_X2 FILLER_58_545 ();
 FILLCELL_X2 FILLER_58_550 ();
 FILLCELL_X1 FILLER_58_552 ();
 FILLCELL_X4 FILLER_58_555 ();
 FILLCELL_X32 FILLER_58_566 ();
 FILLCELL_X32 FILLER_58_598 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X16 FILLER_58_952 ();
 FILLCELL_X1 FILLER_58_968 ();
 FILLCELL_X4 FILLER_58_972 ();
 FILLCELL_X2 FILLER_58_976 ();
 FILLCELL_X1 FILLER_58_978 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X16 FILLER_59_449 ();
 FILLCELL_X8 FILLER_59_465 ();
 FILLCELL_X2 FILLER_59_473 ();
 FILLCELL_X1 FILLER_59_479 ();
 FILLCELL_X32 FILLER_59_488 ();
 FILLCELL_X4 FILLER_59_520 ();
 FILLCELL_X2 FILLER_59_524 ();
 FILLCELL_X2 FILLER_59_556 ();
 FILLCELL_X2 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_581 ();
 FILLCELL_X32 FILLER_59_613 ();
 FILLCELL_X32 FILLER_59_645 ();
 FILLCELL_X32 FILLER_59_677 ();
 FILLCELL_X32 FILLER_59_709 ();
 FILLCELL_X32 FILLER_59_741 ();
 FILLCELL_X32 FILLER_59_773 ();
 FILLCELL_X32 FILLER_59_805 ();
 FILLCELL_X32 FILLER_59_837 ();
 FILLCELL_X32 FILLER_59_869 ();
 FILLCELL_X32 FILLER_59_901 ();
 FILLCELL_X16 FILLER_59_933 ();
 FILLCELL_X8 FILLER_59_949 ();
 FILLCELL_X1 FILLER_59_957 ();
 FILLCELL_X16 FILLER_59_961 ();
 FILLCELL_X2 FILLER_59_977 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X4 FILLER_60_449 ();
 FILLCELL_X2 FILLER_60_453 ();
 FILLCELL_X1 FILLER_60_455 ();
 FILLCELL_X4 FILLER_60_463 ();
 FILLCELL_X2 FILLER_60_467 ();
 FILLCELL_X2 FILLER_60_488 ();
 FILLCELL_X32 FILLER_60_495 ();
 FILLCELL_X16 FILLER_60_527 ();
 FILLCELL_X4 FILLER_60_543 ();
 FILLCELL_X1 FILLER_60_547 ();
 FILLCELL_X1 FILLER_60_552 ();
 FILLCELL_X32 FILLER_60_557 ();
 FILLCELL_X32 FILLER_60_589 ();
 FILLCELL_X8 FILLER_60_621 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X16 FILLER_60_952 ();
 FILLCELL_X8 FILLER_60_968 ();
 FILLCELL_X2 FILLER_60_976 ();
 FILLCELL_X1 FILLER_60_978 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_470 ();
 FILLCELL_X32 FILLER_61_502 ();
 FILLCELL_X32 FILLER_61_534 ();
 FILLCELL_X32 FILLER_61_566 ();
 FILLCELL_X32 FILLER_61_598 ();
 FILLCELL_X32 FILLER_61_630 ();
 FILLCELL_X32 FILLER_61_662 ();
 FILLCELL_X32 FILLER_61_694 ();
 FILLCELL_X32 FILLER_61_726 ();
 FILLCELL_X32 FILLER_61_758 ();
 FILLCELL_X32 FILLER_61_790 ();
 FILLCELL_X32 FILLER_61_822 ();
 FILLCELL_X32 FILLER_61_854 ();
 FILLCELL_X32 FILLER_61_886 ();
 FILLCELL_X32 FILLER_61_918 ();
 FILLCELL_X16 FILLER_61_950 ();
 FILLCELL_X8 FILLER_61_966 ();
 FILLCELL_X4 FILLER_61_974 ();
 FILLCELL_X1 FILLER_61_978 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X16 FILLER_62_449 ();
 FILLCELL_X4 FILLER_62_465 ();
 FILLCELL_X1 FILLER_62_469 ();
 FILLCELL_X4 FILLER_62_481 ();
 FILLCELL_X2 FILLER_62_485 ();
 FILLCELL_X1 FILLER_62_491 ();
 FILLCELL_X1 FILLER_62_497 ();
 FILLCELL_X8 FILLER_62_525 ();
 FILLCELL_X2 FILLER_62_533 ();
 FILLCELL_X1 FILLER_62_535 ();
 FILLCELL_X32 FILLER_62_560 ();
 FILLCELL_X32 FILLER_62_592 ();
 FILLCELL_X4 FILLER_62_624 ();
 FILLCELL_X2 FILLER_62_628 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X8 FILLER_62_952 ();
 FILLCELL_X4 FILLER_62_960 ();
 FILLCELL_X2 FILLER_62_964 ();
 FILLCELL_X1 FILLER_62_966 ();
 FILLCELL_X8 FILLER_62_970 ();
 FILLCELL_X1 FILLER_62_978 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X16 FILLER_63_449 ();
 FILLCELL_X4 FILLER_63_465 ();
 FILLCELL_X1 FILLER_63_469 ();
 FILLCELL_X32 FILLER_63_487 ();
 FILLCELL_X8 FILLER_63_519 ();
 FILLCELL_X2 FILLER_63_527 ();
 FILLCELL_X2 FILLER_63_536 ();
 FILLCELL_X32 FILLER_63_541 ();
 FILLCELL_X32 FILLER_63_573 ();
 FILLCELL_X32 FILLER_63_605 ();
 FILLCELL_X32 FILLER_63_637 ();
 FILLCELL_X32 FILLER_63_669 ();
 FILLCELL_X32 FILLER_63_701 ();
 FILLCELL_X32 FILLER_63_733 ();
 FILLCELL_X32 FILLER_63_765 ();
 FILLCELL_X32 FILLER_63_797 ();
 FILLCELL_X32 FILLER_63_829 ();
 FILLCELL_X32 FILLER_63_861 ();
 FILLCELL_X32 FILLER_63_893 ();
 FILLCELL_X32 FILLER_63_925 ();
 FILLCELL_X16 FILLER_63_957 ();
 FILLCELL_X4 FILLER_63_973 ();
 FILLCELL_X2 FILLER_63_977 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X16 FILLER_64_481 ();
 FILLCELL_X8 FILLER_64_497 ();
 FILLCELL_X1 FILLER_64_505 ();
 FILLCELL_X32 FILLER_64_511 ();
 FILLCELL_X32 FILLER_64_543 ();
 FILLCELL_X32 FILLER_64_575 ();
 FILLCELL_X16 FILLER_64_607 ();
 FILLCELL_X8 FILLER_64_623 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X16 FILLER_64_952 ();
 FILLCELL_X8 FILLER_64_968 ();
 FILLCELL_X2 FILLER_64_976 ();
 FILLCELL_X1 FILLER_64_978 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X2 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_455 ();
 FILLCELL_X16 FILLER_65_487 ();
 FILLCELL_X4 FILLER_65_503 ();
 FILLCELL_X1 FILLER_65_507 ();
 FILLCELL_X8 FILLER_65_512 ();
 FILLCELL_X1 FILLER_65_520 ();
 FILLCELL_X2 FILLER_65_528 ();
 FILLCELL_X1 FILLER_65_534 ();
 FILLCELL_X4 FILLER_65_541 ();
 FILLCELL_X2 FILLER_65_545 ();
 FILLCELL_X1 FILLER_65_547 ();
 FILLCELL_X4 FILLER_65_550 ();
 FILLCELL_X2 FILLER_65_554 ();
 FILLCELL_X1 FILLER_65_556 ();
 FILLCELL_X32 FILLER_65_576 ();
 FILLCELL_X32 FILLER_65_608 ();
 FILLCELL_X32 FILLER_65_640 ();
 FILLCELL_X32 FILLER_65_672 ();
 FILLCELL_X32 FILLER_65_704 ();
 FILLCELL_X32 FILLER_65_736 ();
 FILLCELL_X32 FILLER_65_768 ();
 FILLCELL_X32 FILLER_65_800 ();
 FILLCELL_X32 FILLER_65_832 ();
 FILLCELL_X32 FILLER_65_864 ();
 FILLCELL_X32 FILLER_65_896 ();
 FILLCELL_X8 FILLER_65_928 ();
 FILLCELL_X2 FILLER_65_936 ();
 FILLCELL_X1 FILLER_65_938 ();
 FILLCELL_X8 FILLER_65_943 ();
 FILLCELL_X4 FILLER_65_951 ();
 FILLCELL_X16 FILLER_65_958 ();
 FILLCELL_X4 FILLER_65_974 ();
 FILLCELL_X1 FILLER_65_978 ();
 FILLCELL_X8 FILLER_66_1 ();
 FILLCELL_X4 FILLER_66_9 ();
 FILLCELL_X1 FILLER_66_13 ();
 FILLCELL_X32 FILLER_66_17 ();
 FILLCELL_X32 FILLER_66_49 ();
 FILLCELL_X32 FILLER_66_81 ();
 FILLCELL_X32 FILLER_66_113 ();
 FILLCELL_X32 FILLER_66_145 ();
 FILLCELL_X32 FILLER_66_177 ();
 FILLCELL_X32 FILLER_66_209 ();
 FILLCELL_X32 FILLER_66_241 ();
 FILLCELL_X32 FILLER_66_273 ();
 FILLCELL_X32 FILLER_66_305 ();
 FILLCELL_X32 FILLER_66_337 ();
 FILLCELL_X32 FILLER_66_369 ();
 FILLCELL_X32 FILLER_66_401 ();
 FILLCELL_X8 FILLER_66_433 ();
 FILLCELL_X4 FILLER_66_441 ();
 FILLCELL_X1 FILLER_66_445 ();
 FILLCELL_X4 FILLER_66_463 ();
 FILLCELL_X2 FILLER_66_467 ();
 FILLCELL_X1 FILLER_66_469 ();
 FILLCELL_X8 FILLER_66_491 ();
 FILLCELL_X1 FILLER_66_499 ();
 FILLCELL_X4 FILLER_66_520 ();
 FILLCELL_X1 FILLER_66_524 ();
 FILLCELL_X32 FILLER_66_530 ();
 FILLCELL_X32 FILLER_66_562 ();
 FILLCELL_X32 FILLER_66_594 ();
 FILLCELL_X4 FILLER_66_626 ();
 FILLCELL_X1 FILLER_66_630 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X16 FILLER_66_952 ();
 FILLCELL_X8 FILLER_66_968 ();
 FILLCELL_X2 FILLER_66_976 ();
 FILLCELL_X1 FILLER_66_978 ();
 FILLCELL_X16 FILLER_67_1 ();
 FILLCELL_X4 FILLER_67_17 ();
 FILLCELL_X1 FILLER_67_21 ();
 FILLCELL_X32 FILLER_67_26 ();
 FILLCELL_X32 FILLER_67_58 ();
 FILLCELL_X32 FILLER_67_90 ();
 FILLCELL_X32 FILLER_67_122 ();
 FILLCELL_X32 FILLER_67_154 ();
 FILLCELL_X32 FILLER_67_186 ();
 FILLCELL_X32 FILLER_67_218 ();
 FILLCELL_X32 FILLER_67_250 ();
 FILLCELL_X32 FILLER_67_282 ();
 FILLCELL_X32 FILLER_67_314 ();
 FILLCELL_X32 FILLER_67_346 ();
 FILLCELL_X32 FILLER_67_378 ();
 FILLCELL_X32 FILLER_67_410 ();
 FILLCELL_X8 FILLER_67_442 ();
 FILLCELL_X2 FILLER_67_450 ();
 FILLCELL_X1 FILLER_67_452 ();
 FILLCELL_X16 FILLER_67_460 ();
 FILLCELL_X2 FILLER_67_476 ();
 FILLCELL_X1 FILLER_67_478 ();
 FILLCELL_X32 FILLER_67_494 ();
 FILLCELL_X32 FILLER_67_526 ();
 FILLCELL_X32 FILLER_67_558 ();
 FILLCELL_X32 FILLER_67_590 ();
 FILLCELL_X32 FILLER_67_622 ();
 FILLCELL_X32 FILLER_67_654 ();
 FILLCELL_X32 FILLER_67_686 ();
 FILLCELL_X32 FILLER_67_718 ();
 FILLCELL_X32 FILLER_67_750 ();
 FILLCELL_X32 FILLER_67_782 ();
 FILLCELL_X32 FILLER_67_814 ();
 FILLCELL_X32 FILLER_67_846 ();
 FILLCELL_X32 FILLER_67_878 ();
 FILLCELL_X32 FILLER_67_910 ();
 FILLCELL_X32 FILLER_67_942 ();
 FILLCELL_X4 FILLER_67_974 ();
 FILLCELL_X1 FILLER_67_978 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X16 FILLER_68_481 ();
 FILLCELL_X8 FILLER_68_497 ();
 FILLCELL_X4 FILLER_68_505 ();
 FILLCELL_X1 FILLER_68_509 ();
 FILLCELL_X32 FILLER_68_515 ();
 FILLCELL_X32 FILLER_68_547 ();
 FILLCELL_X32 FILLER_68_579 ();
 FILLCELL_X16 FILLER_68_611 ();
 FILLCELL_X4 FILLER_68_627 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X16 FILLER_68_952 ();
 FILLCELL_X8 FILLER_68_968 ();
 FILLCELL_X2 FILLER_68_976 ();
 FILLCELL_X1 FILLER_68_978 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X4 FILLER_69_449 ();
 FILLCELL_X2 FILLER_69_453 ();
 FILLCELL_X1 FILLER_69_455 ();
 FILLCELL_X32 FILLER_69_460 ();
 FILLCELL_X8 FILLER_69_492 ();
 FILLCELL_X2 FILLER_69_500 ();
 FILLCELL_X1 FILLER_69_502 ();
 FILLCELL_X8 FILLER_69_507 ();
 FILLCELL_X2 FILLER_69_515 ();
 FILLCELL_X32 FILLER_69_530 ();
 FILLCELL_X32 FILLER_69_562 ();
 FILLCELL_X32 FILLER_69_594 ();
 FILLCELL_X32 FILLER_69_626 ();
 FILLCELL_X32 FILLER_69_658 ();
 FILLCELL_X32 FILLER_69_690 ();
 FILLCELL_X32 FILLER_69_722 ();
 FILLCELL_X32 FILLER_69_754 ();
 FILLCELL_X32 FILLER_69_786 ();
 FILLCELL_X32 FILLER_69_818 ();
 FILLCELL_X32 FILLER_69_850 ();
 FILLCELL_X32 FILLER_69_882 ();
 FILLCELL_X32 FILLER_69_914 ();
 FILLCELL_X32 FILLER_69_946 ();
 FILLCELL_X1 FILLER_69_978 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X16 FILLER_70_417 ();
 FILLCELL_X8 FILLER_70_433 ();
 FILLCELL_X4 FILLER_70_441 ();
 FILLCELL_X2 FILLER_70_445 ();
 FILLCELL_X8 FILLER_70_464 ();
 FILLCELL_X2 FILLER_70_472 ();
 FILLCELL_X8 FILLER_70_491 ();
 FILLCELL_X2 FILLER_70_499 ();
 FILLCELL_X32 FILLER_70_534 ();
 FILLCELL_X32 FILLER_70_566 ();
 FILLCELL_X32 FILLER_70_598 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X16 FILLER_70_952 ();
 FILLCELL_X8 FILLER_70_968 ();
 FILLCELL_X2 FILLER_70_976 ();
 FILLCELL_X1 FILLER_70_978 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X4 FILLER_71_449 ();
 FILLCELL_X8 FILLER_71_460 ();
 FILLCELL_X4 FILLER_71_468 ();
 FILLCELL_X2 FILLER_71_472 ();
 FILLCELL_X4 FILLER_71_485 ();
 FILLCELL_X16 FILLER_71_494 ();
 FILLCELL_X8 FILLER_71_510 ();
 FILLCELL_X4 FILLER_71_518 ();
 FILLCELL_X2 FILLER_71_522 ();
 FILLCELL_X1 FILLER_71_524 ();
 FILLCELL_X2 FILLER_71_530 ();
 FILLCELL_X32 FILLER_71_538 ();
 FILLCELL_X32 FILLER_71_570 ();
 FILLCELL_X32 FILLER_71_602 ();
 FILLCELL_X32 FILLER_71_634 ();
 FILLCELL_X32 FILLER_71_666 ();
 FILLCELL_X32 FILLER_71_698 ();
 FILLCELL_X32 FILLER_71_730 ();
 FILLCELL_X32 FILLER_71_762 ();
 FILLCELL_X32 FILLER_71_794 ();
 FILLCELL_X32 FILLER_71_826 ();
 FILLCELL_X32 FILLER_71_858 ();
 FILLCELL_X32 FILLER_71_890 ();
 FILLCELL_X32 FILLER_71_922 ();
 FILLCELL_X16 FILLER_71_954 ();
 FILLCELL_X8 FILLER_71_970 ();
 FILLCELL_X1 FILLER_71_978 ();
 FILLCELL_X4 FILLER_72_1 ();
 FILLCELL_X2 FILLER_72_5 ();
 FILLCELL_X1 FILLER_72_7 ();
 FILLCELL_X32 FILLER_72_11 ();
 FILLCELL_X32 FILLER_72_43 ();
 FILLCELL_X32 FILLER_72_75 ();
 FILLCELL_X32 FILLER_72_107 ();
 FILLCELL_X32 FILLER_72_139 ();
 FILLCELL_X32 FILLER_72_171 ();
 FILLCELL_X32 FILLER_72_203 ();
 FILLCELL_X32 FILLER_72_235 ();
 FILLCELL_X32 FILLER_72_267 ();
 FILLCELL_X32 FILLER_72_299 ();
 FILLCELL_X32 FILLER_72_331 ();
 FILLCELL_X32 FILLER_72_363 ();
 FILLCELL_X32 FILLER_72_395 ();
 FILLCELL_X16 FILLER_72_427 ();
 FILLCELL_X8 FILLER_72_443 ();
 FILLCELL_X4 FILLER_72_451 ();
 FILLCELL_X1 FILLER_72_455 ();
 FILLCELL_X32 FILLER_72_463 ();
 FILLCELL_X4 FILLER_72_495 ();
 FILLCELL_X1 FILLER_72_499 ();
 FILLCELL_X8 FILLER_72_507 ();
 FILLCELL_X4 FILLER_72_515 ();
 FILLCELL_X2 FILLER_72_519 ();
 FILLCELL_X32 FILLER_72_542 ();
 FILLCELL_X32 FILLER_72_574 ();
 FILLCELL_X16 FILLER_72_606 ();
 FILLCELL_X8 FILLER_72_622 ();
 FILLCELL_X1 FILLER_72_630 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X16 FILLER_72_952 ();
 FILLCELL_X8 FILLER_72_968 ();
 FILLCELL_X2 FILLER_72_976 ();
 FILLCELL_X1 FILLER_72_978 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X2 FILLER_73_33 ();
 FILLCELL_X1 FILLER_73_35 ();
 FILLCELL_X32 FILLER_73_40 ();
 FILLCELL_X32 FILLER_73_72 ();
 FILLCELL_X32 FILLER_73_104 ();
 FILLCELL_X32 FILLER_73_136 ();
 FILLCELL_X32 FILLER_73_168 ();
 FILLCELL_X32 FILLER_73_200 ();
 FILLCELL_X32 FILLER_73_232 ();
 FILLCELL_X32 FILLER_73_264 ();
 FILLCELL_X32 FILLER_73_296 ();
 FILLCELL_X32 FILLER_73_328 ();
 FILLCELL_X32 FILLER_73_360 ();
 FILLCELL_X32 FILLER_73_392 ();
 FILLCELL_X8 FILLER_73_424 ();
 FILLCELL_X2 FILLER_73_432 ();
 FILLCELL_X16 FILLER_73_438 ();
 FILLCELL_X2 FILLER_73_454 ();
 FILLCELL_X8 FILLER_73_467 ();
 FILLCELL_X4 FILLER_73_475 ();
 FILLCELL_X2 FILLER_73_479 ();
 FILLCELL_X16 FILLER_73_485 ();
 FILLCELL_X4 FILLER_73_501 ();
 FILLCELL_X2 FILLER_73_505 ();
 FILLCELL_X1 FILLER_73_507 ();
 FILLCELL_X8 FILLER_73_512 ();
 FILLCELL_X32 FILLER_73_531 ();
 FILLCELL_X32 FILLER_73_563 ();
 FILLCELL_X32 FILLER_73_595 ();
 FILLCELL_X32 FILLER_73_627 ();
 FILLCELL_X32 FILLER_73_659 ();
 FILLCELL_X32 FILLER_73_691 ();
 FILLCELL_X32 FILLER_73_723 ();
 FILLCELL_X32 FILLER_73_755 ();
 FILLCELL_X32 FILLER_73_787 ();
 FILLCELL_X32 FILLER_73_819 ();
 FILLCELL_X32 FILLER_73_851 ();
 FILLCELL_X32 FILLER_73_883 ();
 FILLCELL_X32 FILLER_73_915 ();
 FILLCELL_X32 FILLER_73_947 ();
 FILLCELL_X4 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_8 ();
 FILLCELL_X32 FILLER_74_40 ();
 FILLCELL_X32 FILLER_74_72 ();
 FILLCELL_X32 FILLER_74_104 ();
 FILLCELL_X32 FILLER_74_136 ();
 FILLCELL_X32 FILLER_74_168 ();
 FILLCELL_X32 FILLER_74_200 ();
 FILLCELL_X32 FILLER_74_232 ();
 FILLCELL_X32 FILLER_74_264 ();
 FILLCELL_X32 FILLER_74_296 ();
 FILLCELL_X32 FILLER_74_328 ();
 FILLCELL_X32 FILLER_74_360 ();
 FILLCELL_X32 FILLER_74_392 ();
 FILLCELL_X16 FILLER_74_424 ();
 FILLCELL_X8 FILLER_74_440 ();
 FILLCELL_X1 FILLER_74_448 ();
 FILLCELL_X16 FILLER_74_468 ();
 FILLCELL_X1 FILLER_74_484 ();
 FILLCELL_X8 FILLER_74_491 ();
 FILLCELL_X4 FILLER_74_499 ();
 FILLCELL_X8 FILLER_74_520 ();
 FILLCELL_X4 FILLER_74_528 ();
 FILLCELL_X32 FILLER_74_538 ();
 FILLCELL_X32 FILLER_74_570 ();
 FILLCELL_X16 FILLER_74_602 ();
 FILLCELL_X8 FILLER_74_618 ();
 FILLCELL_X4 FILLER_74_626 ();
 FILLCELL_X1 FILLER_74_630 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X16 FILLER_74_952 ();
 FILLCELL_X8 FILLER_74_968 ();
 FILLCELL_X2 FILLER_74_976 ();
 FILLCELL_X1 FILLER_74_978 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X8 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_491 ();
 FILLCELL_X8 FILLER_75_523 ();
 FILLCELL_X4 FILLER_75_531 ();
 FILLCELL_X1 FILLER_75_535 ();
 FILLCELL_X32 FILLER_75_538 ();
 FILLCELL_X32 FILLER_75_570 ();
 FILLCELL_X32 FILLER_75_602 ();
 FILLCELL_X32 FILLER_75_634 ();
 FILLCELL_X32 FILLER_75_666 ();
 FILLCELL_X32 FILLER_75_698 ();
 FILLCELL_X32 FILLER_75_730 ();
 FILLCELL_X32 FILLER_75_762 ();
 FILLCELL_X32 FILLER_75_794 ();
 FILLCELL_X32 FILLER_75_826 ();
 FILLCELL_X32 FILLER_75_858 ();
 FILLCELL_X32 FILLER_75_890 ();
 FILLCELL_X32 FILLER_75_922 ();
 FILLCELL_X16 FILLER_75_954 ();
 FILLCELL_X8 FILLER_75_970 ();
 FILLCELL_X1 FILLER_75_978 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X16 FILLER_76_449 ();
 FILLCELL_X8 FILLER_76_465 ();
 FILLCELL_X2 FILLER_76_473 ();
 FILLCELL_X1 FILLER_76_475 ();
 FILLCELL_X32 FILLER_76_495 ();
 FILLCELL_X2 FILLER_76_527 ();
 FILLCELL_X32 FILLER_76_548 ();
 FILLCELL_X32 FILLER_76_580 ();
 FILLCELL_X16 FILLER_76_612 ();
 FILLCELL_X2 FILLER_76_628 ();
 FILLCELL_X1 FILLER_76_630 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X16 FILLER_76_952 ();
 FILLCELL_X8 FILLER_76_968 ();
 FILLCELL_X2 FILLER_76_976 ();
 FILLCELL_X1 FILLER_76_978 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X16 FILLER_77_961 ();
 FILLCELL_X2 FILLER_77_977 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X16 FILLER_78_952 ();
 FILLCELL_X8 FILLER_78_968 ();
 FILLCELL_X2 FILLER_78_976 ();
 FILLCELL_X1 FILLER_78_978 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X16 FILLER_79_961 ();
 FILLCELL_X2 FILLER_79_977 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X16 FILLER_80_952 ();
 FILLCELL_X8 FILLER_80_968 ();
 FILLCELL_X2 FILLER_80_976 ();
 FILLCELL_X1 FILLER_80_978 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X16 FILLER_81_961 ();
 FILLCELL_X2 FILLER_81_977 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X16 FILLER_82_952 ();
 FILLCELL_X8 FILLER_82_968 ();
 FILLCELL_X2 FILLER_82_976 ();
 FILLCELL_X1 FILLER_82_978 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X16 FILLER_83_961 ();
 FILLCELL_X2 FILLER_83_977 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X16 FILLER_84_952 ();
 FILLCELL_X8 FILLER_84_968 ();
 FILLCELL_X2 FILLER_84_976 ();
 FILLCELL_X1 FILLER_84_978 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X16 FILLER_85_961 ();
 FILLCELL_X2 FILLER_85_977 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X16 FILLER_86_952 ();
 FILLCELL_X8 FILLER_86_968 ();
 FILLCELL_X2 FILLER_86_976 ();
 FILLCELL_X1 FILLER_86_978 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X16 FILLER_87_961 ();
 FILLCELL_X2 FILLER_87_977 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X16 FILLER_88_952 ();
 FILLCELL_X8 FILLER_88_968 ();
 FILLCELL_X2 FILLER_88_976 ();
 FILLCELL_X1 FILLER_88_978 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X16 FILLER_89_961 ();
 FILLCELL_X2 FILLER_89_977 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X16 FILLER_90_952 ();
 FILLCELL_X8 FILLER_90_968 ();
 FILLCELL_X2 FILLER_90_976 ();
 FILLCELL_X1 FILLER_90_978 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X16 FILLER_91_961 ();
 FILLCELL_X2 FILLER_91_977 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X16 FILLER_92_952 ();
 FILLCELL_X8 FILLER_92_968 ();
 FILLCELL_X2 FILLER_92_976 ();
 FILLCELL_X1 FILLER_92_978 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X16 FILLER_93_961 ();
 FILLCELL_X2 FILLER_93_977 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X16 FILLER_94_952 ();
 FILLCELL_X8 FILLER_94_968 ();
 FILLCELL_X2 FILLER_94_976 ();
 FILLCELL_X1 FILLER_94_978 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X16 FILLER_95_961 ();
 FILLCELL_X2 FILLER_95_977 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X16 FILLER_96_952 ();
 FILLCELL_X8 FILLER_96_968 ();
 FILLCELL_X2 FILLER_96_976 ();
 FILLCELL_X1 FILLER_96_978 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X16 FILLER_97_961 ();
 FILLCELL_X2 FILLER_97_977 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X16 FILLER_98_952 ();
 FILLCELL_X8 FILLER_98_968 ();
 FILLCELL_X2 FILLER_98_976 ();
 FILLCELL_X1 FILLER_98_978 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X16 FILLER_99_961 ();
 FILLCELL_X2 FILLER_99_977 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X16 FILLER_100_952 ();
 FILLCELL_X8 FILLER_100_968 ();
 FILLCELL_X2 FILLER_100_976 ();
 FILLCELL_X1 FILLER_100_978 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X16 FILLER_101_961 ();
 FILLCELL_X2 FILLER_101_977 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X16 FILLER_102_952 ();
 FILLCELL_X8 FILLER_102_968 ();
 FILLCELL_X2 FILLER_102_976 ();
 FILLCELL_X1 FILLER_102_978 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X16 FILLER_103_961 ();
 FILLCELL_X2 FILLER_103_977 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X16 FILLER_104_952 ();
 FILLCELL_X8 FILLER_104_968 ();
 FILLCELL_X2 FILLER_104_976 ();
 FILLCELL_X1 FILLER_104_978 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X16 FILLER_105_961 ();
 FILLCELL_X2 FILLER_105_977 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X16 FILLER_106_952 ();
 FILLCELL_X8 FILLER_106_968 ();
 FILLCELL_X2 FILLER_106_976 ();
 FILLCELL_X1 FILLER_106_978 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X16 FILLER_107_961 ();
 FILLCELL_X2 FILLER_107_977 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X32 FILLER_108_856 ();
 FILLCELL_X32 FILLER_108_888 ();
 FILLCELL_X32 FILLER_108_920 ();
 FILLCELL_X16 FILLER_108_952 ();
 FILLCELL_X8 FILLER_108_968 ();
 FILLCELL_X2 FILLER_108_976 ();
 FILLCELL_X1 FILLER_108_978 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X16 FILLER_109_961 ();
 FILLCELL_X2 FILLER_109_977 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X16 FILLER_110_952 ();
 FILLCELL_X8 FILLER_110_968 ();
 FILLCELL_X2 FILLER_110_976 ();
 FILLCELL_X1 FILLER_110_978 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X16 FILLER_111_961 ();
 FILLCELL_X2 FILLER_111_977 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X16 FILLER_112_952 ();
 FILLCELL_X8 FILLER_112_968 ();
 FILLCELL_X2 FILLER_112_976 ();
 FILLCELL_X1 FILLER_112_978 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X32 FILLER_113_833 ();
 FILLCELL_X32 FILLER_113_865 ();
 FILLCELL_X32 FILLER_113_897 ();
 FILLCELL_X32 FILLER_113_929 ();
 FILLCELL_X16 FILLER_113_961 ();
 FILLCELL_X2 FILLER_113_977 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X16 FILLER_114_952 ();
 FILLCELL_X8 FILLER_114_968 ();
 FILLCELL_X2 FILLER_114_976 ();
 FILLCELL_X1 FILLER_114_978 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X32 FILLER_115_801 ();
 FILLCELL_X32 FILLER_115_833 ();
 FILLCELL_X32 FILLER_115_865 ();
 FILLCELL_X32 FILLER_115_897 ();
 FILLCELL_X32 FILLER_115_929 ();
 FILLCELL_X16 FILLER_115_961 ();
 FILLCELL_X2 FILLER_115_977 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X32 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_888 ();
 FILLCELL_X32 FILLER_116_920 ();
 FILLCELL_X16 FILLER_116_952 ();
 FILLCELL_X8 FILLER_116_968 ();
 FILLCELL_X2 FILLER_116_976 ();
 FILLCELL_X1 FILLER_116_978 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X32 FILLER_117_801 ();
 FILLCELL_X32 FILLER_117_833 ();
 FILLCELL_X32 FILLER_117_865 ();
 FILLCELL_X32 FILLER_117_897 ();
 FILLCELL_X32 FILLER_117_929 ();
 FILLCELL_X16 FILLER_117_961 ();
 FILLCELL_X2 FILLER_117_977 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X16 FILLER_118_952 ();
 FILLCELL_X8 FILLER_118_968 ();
 FILLCELL_X2 FILLER_118_976 ();
 FILLCELL_X1 FILLER_118_978 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X16 FILLER_119_961 ();
 FILLCELL_X2 FILLER_119_977 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X16 FILLER_120_952 ();
 FILLCELL_X8 FILLER_120_968 ();
 FILLCELL_X2 FILLER_120_976 ();
 FILLCELL_X1 FILLER_120_978 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X16 FILLER_121_961 ();
 FILLCELL_X2 FILLER_121_977 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X16 FILLER_122_952 ();
 FILLCELL_X8 FILLER_122_968 ();
 FILLCELL_X2 FILLER_122_976 ();
 FILLCELL_X1 FILLER_122_978 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X16 FILLER_123_961 ();
 FILLCELL_X2 FILLER_123_977 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X16 FILLER_124_952 ();
 FILLCELL_X8 FILLER_124_968 ();
 FILLCELL_X2 FILLER_124_976 ();
 FILLCELL_X1 FILLER_124_978 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X16 FILLER_125_961 ();
 FILLCELL_X2 FILLER_125_977 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X16 FILLER_126_952 ();
 FILLCELL_X8 FILLER_126_968 ();
 FILLCELL_X2 FILLER_126_976 ();
 FILLCELL_X1 FILLER_126_978 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X16 FILLER_127_961 ();
 FILLCELL_X2 FILLER_127_977 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X16 FILLER_128_952 ();
 FILLCELL_X8 FILLER_128_968 ();
 FILLCELL_X2 FILLER_128_976 ();
 FILLCELL_X1 FILLER_128_978 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X16 FILLER_129_961 ();
 FILLCELL_X2 FILLER_129_977 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X16 FILLER_130_952 ();
 FILLCELL_X8 FILLER_130_968 ();
 FILLCELL_X2 FILLER_130_976 ();
 FILLCELL_X1 FILLER_130_978 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X8 FILLER_131_481 ();
 FILLCELL_X4 FILLER_131_489 ();
 FILLCELL_X16 FILLER_131_496 ();
 FILLCELL_X4 FILLER_131_512 ();
 FILLCELL_X2 FILLER_131_516 ();
 FILLCELL_X1 FILLER_131_518 ();
 FILLCELL_X2 FILLER_131_523 ();
 FILLCELL_X1 FILLER_131_525 ();
 FILLCELL_X8 FILLER_131_529 ();
 FILLCELL_X4 FILLER_131_537 ();
 FILLCELL_X2 FILLER_131_544 ();
 FILLCELL_X1 FILLER_131_546 ();
 FILLCELL_X32 FILLER_131_550 ();
 FILLCELL_X32 FILLER_131_582 ();
 FILLCELL_X16 FILLER_131_614 ();
 FILLCELL_X1 FILLER_131_630 ();
 FILLCELL_X32 FILLER_131_632 ();
 FILLCELL_X32 FILLER_131_664 ();
 FILLCELL_X32 FILLER_131_696 ();
 FILLCELL_X32 FILLER_131_728 ();
 FILLCELL_X32 FILLER_131_760 ();
 FILLCELL_X32 FILLER_131_792 ();
 FILLCELL_X32 FILLER_131_824 ();
 FILLCELL_X32 FILLER_131_856 ();
 FILLCELL_X32 FILLER_131_888 ();
 FILLCELL_X32 FILLER_131_920 ();
 FILLCELL_X16 FILLER_131_952 ();
 FILLCELL_X8 FILLER_131_968 ();
 FILLCELL_X2 FILLER_131_976 ();
 FILLCELL_X1 FILLER_131_978 ();
endmodule
