module parameterized_decade_counter (clk,
    enable,
    rst_n,
    tc,
    count);
 input clk;
 input enable;
 input rst_n;
 output tc;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net8;

 sky130_fd_sc_hd__nand2_1 _19_ (.A(net6),
    .B(_15_),
    .Y(_04_));
 sky130_fd_sc_hd__nor2_1 _20_ (.A(net5),
    .B(_04_),
    .Y(net7));
 sky130_fd_sc_hd__inv_1 _21_ (.A(net4),
    .Y(_14_));
 sky130_fd_sc_hd__nand2b_1 _22_ (.A_N(net3),
    .B(net2),
    .Y(_05_));
 sky130_fd_sc_hd__nand2b_1 _23_ (.A_N(net2),
    .B(net3),
    .Y(_06_));
 sky130_fd_sc_hd__o21ai_0 _24_ (.A1(net7),
    .A2(_05_),
    .B1(_06_),
    .Y(_00_));
 sky130_fd_sc_hd__nand2b_1 _25_ (.A_N(_16_),
    .B(net2),
    .Y(_07_));
 sky130_fd_sc_hd__o22ai_1 _26_ (.A1(net2),
    .A2(_14_),
    .B1(net7),
    .B2(_07_),
    .Y(_01_));
 sky130_fd_sc_hd__nand2_1 _27_ (.A(net2),
    .B(_17_),
    .Y(_08_));
 sky130_fd_sc_hd__nor3b_1 _28_ (.A(net5),
    .B(_08_),
    .C_N(_04_),
    .Y(_09_));
 sky130_fd_sc_hd__a21o_1 _29_ (.A1(net5),
    .A2(_08_),
    .B1(_09_),
    .X(_02_));
 sky130_fd_sc_hd__nand3_1 _30_ (.A(net2),
    .B(net4),
    .C(net3),
    .Y(_10_));
 sky130_fd_sc_hd__a21bo_1 _31_ (.A1(net4),
    .A2(net3),
    .B1_N(net6),
    .X(_11_));
 sky130_fd_sc_hd__o21ai_0 _32_ (.A1(net6),
    .A2(_10_),
    .B1(_11_),
    .Y(_12_));
 sky130_fd_sc_hd__o21ai_0 _33_ (.A1(net5),
    .A2(_15_),
    .B1(net2),
    .Y(_13_));
 sky130_fd_sc_hd__a22o_1 _34_ (.A1(net5),
    .A2(_12_),
    .B1(_13_),
    .B2(net6),
    .X(_03_));
 sky130_fd_sc_hd__ha_1 _35_ (.A(net3),
    .B(_14_),
    .COUT(_15_),
    .SUM(_16_));
 sky130_fd_sc_hd__ha_1 _36_ (.A(net3),
    .B(net4),
    .COUT(_17_),
    .SUM(_18_));
 sky130_fd_sc_hd__dfrtp_2 \count[0]$_DFFE_PN0P_  (.D(_00_),
    .Q(net3),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \count[1]$_DFFE_PN0P_  (.D(_01_),
    .Q(net4),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \count[2]$_DFFE_PN0P_  (.D(_02_),
    .Q(net5),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \count[3]$_DFFE_PN0P_  (.D(_03_),
    .Q(net6),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1 (.A(net8),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_26 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(enable),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 output2 (.A(net3),
    .X(count[0]));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net4),
    .X(count[1]));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net5),
    .X(count[2]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net6),
    .X(count[3]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net7),
    .X(tc));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net8));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_101 ();
endmodule
