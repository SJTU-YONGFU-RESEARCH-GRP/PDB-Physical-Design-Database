module siso_register (clk,
    enable,
    rst_n,
    serial_in,
    serial_out);
 input clk;
 input enable;
 input rst_n;
 input serial_in;
 output serial_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire \shift_reg[1] ;
 wire \shift_reg[2] ;
 wire \shift_reg[3] ;
 wire \shift_reg[4] ;
 wire \shift_reg[5] ;
 wire \shift_reg[6] ;
 wire \shift_reg[7] ;
 wire net1;
 wire net2;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X1 _26_ (.A(rst_n),
    .Z(_08_));
 BUF_X4 _27_ (.A(enable),
    .Z(_09_));
 MUX2_X1 _28_ (.A(net2),
    .B(\shift_reg[1] ),
    .S(_09_),
    .Z(_10_));
 AND2_X1 _29_ (.A1(_08_),
    .A2(_10_),
    .ZN(_00_));
 MUX2_X1 _30_ (.A(\shift_reg[1] ),
    .B(\shift_reg[2] ),
    .S(_09_),
    .Z(_11_));
 AND2_X1 _31_ (.A1(_08_),
    .A2(_11_),
    .ZN(_01_));
 MUX2_X1 _32_ (.A(\shift_reg[2] ),
    .B(\shift_reg[3] ),
    .S(_09_),
    .Z(_12_));
 AND2_X1 _33_ (.A1(_08_),
    .A2(_12_),
    .ZN(_02_));
 MUX2_X1 _34_ (.A(\shift_reg[3] ),
    .B(\shift_reg[4] ),
    .S(_09_),
    .Z(_13_));
 AND2_X1 _35_ (.A1(_08_),
    .A2(_13_),
    .ZN(_03_));
 MUX2_X1 _36_ (.A(\shift_reg[4] ),
    .B(\shift_reg[5] ),
    .S(_09_),
    .Z(_14_));
 AND2_X1 _37_ (.A1(_08_),
    .A2(_14_),
    .ZN(_04_));
 MUX2_X1 _38_ (.A(\shift_reg[5] ),
    .B(\shift_reg[6] ),
    .S(_09_),
    .Z(_15_));
 AND2_X1 _39_ (.A1(_08_),
    .A2(_15_),
    .ZN(_05_));
 MUX2_X1 _40_ (.A(\shift_reg[6] ),
    .B(\shift_reg[7] ),
    .S(_09_),
    .Z(_16_));
 AND2_X1 _41_ (.A1(_08_),
    .A2(_16_),
    .ZN(_06_));
 MUX2_X1 _42_ (.A(\shift_reg[7] ),
    .B(net1),
    .S(_09_),
    .Z(_17_));
 AND2_X1 _43_ (.A1(_08_),
    .A2(_17_),
    .ZN(_07_));
 DFF_X1 \shift_reg[0]$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net2),
    .QN(_25_));
 DFF_X1 \shift_reg[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[1] ),
    .QN(_24_));
 DFF_X1 \shift_reg[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[2] ),
    .QN(_23_));
 DFF_X1 \shift_reg[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[3] ),
    .QN(_22_));
 DFF_X1 \shift_reg[4]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[4] ),
    .QN(_21_));
 DFF_X1 \shift_reg[5]$_SDFFE_PN0P_  (.D(_05_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[5] ),
    .QN(_20_));
 DFF_X1 \shift_reg[6]$_SDFFE_PN0P_  (.D(_06_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[6] ),
    .QN(_19_));
 DFF_X1 \shift_reg[7]$_SDFFE_PN0P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[7] ),
    .QN(_18_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_49 ();
 BUF_X1 input1 (.A(serial_in),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(serial_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X16 FILLER_0_161 ();
 FILLCELL_X8 FILLER_0_177 ();
 FILLCELL_X2 FILLER_0_185 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X16 FILLER_1_161 ();
 FILLCELL_X8 FILLER_1_177 ();
 FILLCELL_X2 FILLER_1_185 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X16 FILLER_2_161 ();
 FILLCELL_X8 FILLER_2_177 ();
 FILLCELL_X2 FILLER_2_185 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X16 FILLER_3_161 ();
 FILLCELL_X8 FILLER_3_177 ();
 FILLCELL_X2 FILLER_3_185 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X16 FILLER_4_161 ();
 FILLCELL_X8 FILLER_4_177 ();
 FILLCELL_X2 FILLER_4_185 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X16 FILLER_5_161 ();
 FILLCELL_X8 FILLER_5_177 ();
 FILLCELL_X2 FILLER_5_185 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X8 FILLER_6_177 ();
 FILLCELL_X2 FILLER_6_185 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_40 ();
 FILLCELL_X32 FILLER_7_72 ();
 FILLCELL_X32 FILLER_7_104 ();
 FILLCELL_X32 FILLER_7_136 ();
 FILLCELL_X16 FILLER_7_168 ();
 FILLCELL_X2 FILLER_7_184 ();
 FILLCELL_X1 FILLER_7_186 ();
 FILLCELL_X4 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_5 ();
 FILLCELL_X1 FILLER_8_7 ();
 FILLCELL_X8 FILLER_8_25 ();
 FILLCELL_X2 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_52 ();
 FILLCELL_X32 FILLER_8_84 ();
 FILLCELL_X32 FILLER_8_116 ();
 FILLCELL_X32 FILLER_8_148 ();
 FILLCELL_X4 FILLER_8_180 ();
 FILLCELL_X2 FILLER_8_184 ();
 FILLCELL_X1 FILLER_8_186 ();
 FILLCELL_X1 FILLER_9_1 ();
 FILLCELL_X1 FILLER_9_5 ();
 FILLCELL_X1 FILLER_9_13 ();
 FILLCELL_X4 FILLER_9_29 ();
 FILLCELL_X32 FILLER_9_57 ();
 FILLCELL_X32 FILLER_9_89 ();
 FILLCELL_X32 FILLER_9_121 ();
 FILLCELL_X32 FILLER_9_153 ();
 FILLCELL_X2 FILLER_9_185 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_17 ();
 FILLCELL_X2 FILLER_10_35 ();
 FILLCELL_X1 FILLER_10_37 ();
 FILLCELL_X32 FILLER_10_53 ();
 FILLCELL_X32 FILLER_10_85 ();
 FILLCELL_X32 FILLER_10_117 ();
 FILLCELL_X32 FILLER_10_149 ();
 FILLCELL_X4 FILLER_10_181 ();
 FILLCELL_X2 FILLER_10_185 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X16 FILLER_11_161 ();
 FILLCELL_X8 FILLER_11_177 ();
 FILLCELL_X2 FILLER_11_185 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_17 ();
 FILLCELL_X4 FILLER_12_25 ();
 FILLCELL_X2 FILLER_12_29 ();
 FILLCELL_X1 FILLER_12_31 ();
 FILLCELL_X32 FILLER_12_37 ();
 FILLCELL_X32 FILLER_12_69 ();
 FILLCELL_X32 FILLER_12_101 ();
 FILLCELL_X32 FILLER_12_133 ();
 FILLCELL_X16 FILLER_12_165 ();
 FILLCELL_X4 FILLER_12_181 ();
 FILLCELL_X2 FILLER_12_185 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X8 FILLER_13_17 ();
 FILLCELL_X2 FILLER_13_25 ();
 FILLCELL_X32 FILLER_13_55 ();
 FILLCELL_X32 FILLER_13_87 ();
 FILLCELL_X32 FILLER_13_119 ();
 FILLCELL_X32 FILLER_13_151 ();
 FILLCELL_X4 FILLER_13_183 ();
 FILLCELL_X1 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X4 FILLER_14_36 ();
 FILLCELL_X1 FILLER_14_40 ();
 FILLCELL_X32 FILLER_14_48 ();
 FILLCELL_X32 FILLER_14_80 ();
 FILLCELL_X32 FILLER_14_112 ();
 FILLCELL_X32 FILLER_14_144 ();
 FILLCELL_X8 FILLER_14_176 ();
 FILLCELL_X2 FILLER_14_184 ();
 FILLCELL_X1 FILLER_14_186 ();
 FILLCELL_X2 FILLER_15_11 ();
 FILLCELL_X2 FILLER_15_30 ();
 FILLCELL_X32 FILLER_15_53 ();
 FILLCELL_X32 FILLER_15_85 ();
 FILLCELL_X32 FILLER_15_117 ();
 FILLCELL_X32 FILLER_15_149 ();
 FILLCELL_X4 FILLER_15_181 ();
 FILLCELL_X2 FILLER_15_185 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X4 FILLER_16_24 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X16 FILLER_16_161 ();
 FILLCELL_X8 FILLER_16_177 ();
 FILLCELL_X2 FILLER_16_185 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X16 FILLER_17_161 ();
 FILLCELL_X8 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_185 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X16 FILLER_18_161 ();
 FILLCELL_X8 FILLER_18_177 ();
 FILLCELL_X2 FILLER_18_185 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X8 FILLER_19_177 ();
 FILLCELL_X2 FILLER_19_185 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X16 FILLER_20_161 ();
 FILLCELL_X8 FILLER_20_177 ();
 FILLCELL_X2 FILLER_20_185 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X8 FILLER_21_177 ();
 FILLCELL_X2 FILLER_21_185 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X8 FILLER_22_177 ();
 FILLCELL_X2 FILLER_22_185 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X16 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_177 ();
 FILLCELL_X2 FILLER_23_185 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X16 FILLER_24_161 ();
 FILLCELL_X8 FILLER_24_177 ();
 FILLCELL_X2 FILLER_24_185 ();
endmodule
