module multi_phase_pwm_controller (clk,
    enable,
    rst_n,
    deadtime,
    duty,
    pwm_n_out,
    pwm_p_out);
 input clk;
 input enable;
 input rst_n;
 input [5:0] deadtime;
 input [7:0] duty;
 output [2:0] pwm_n_out;
 output [2:0] pwm_p_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire _494_;
 wire _495_;
 wire _496_;
 wire _497_;
 wire _498_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _499_ (.I(net13),
    .ZN(_464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _500_ (.I(_327_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _501_ (.I(net14),
    .ZN(_461_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _502_ (.I(\counter[4] ),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _503_ (.I(\counter[6] ),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _504_ (.I(\counter[2] ),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _505_ (.I(\counter[7] ),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _506_ (.I(\counter[3] ),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _507_ (.A1(\counter[0] ),
    .A2(_411_),
    .B(\counter[2] ),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _508_ (.A1(_274_),
    .A2(_014_),
    .B(_270_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _509_ (.A1(\counter[5] ),
    .A2(_015_),
    .B(\counter[6] ),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _510_ (.A1(_258_),
    .A2(_016_),
    .ZN(_347_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _511_ (.A1(\counter[2] ),
    .A2(_365_),
    .B(\counter[3] ),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _512_ (.A1(_270_),
    .A2(_017_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _513_ (.A1(\counter[5] ),
    .A2(_018_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _514_ (.A1(_262_),
    .A2(_019_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _515_ (.I(_020_),
    .ZN(_350_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _516_ (.A1(\counter[5] ),
    .A2(_015_),
    .ZN(_353_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _517_ (.A1(\counter[4] ),
    .A2(_017_),
    .ZN(_356_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _518_ (.A1(_274_),
    .A2(_014_),
    .ZN(_359_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _519_ (.A1(\counter[2] ),
    .A2(_365_),
    .Z(_362_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _520_ (.I(_413_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _521_ (.A1(_274_),
    .A2(_021_),
    .B(_270_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _522_ (.A1(\counter[5] ),
    .A2(_022_),
    .B(\counter[6] ),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _523_ (.A1(\counter[7] ),
    .A2(_023_),
    .ZN(_396_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _524_ (.I(\counter[5] ),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _525_ (.A1(\counter[2] ),
    .A2(\counter[1] ),
    .B(\counter[3] ),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _526_ (.A1(_270_),
    .A2(_024_),
    .B(_266_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _527_ (.A1(\counter[6] ),
    .A2(_025_),
    .ZN(_399_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _528_ (.A1(_266_),
    .A2(_022_),
    .ZN(_402_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _529_ (.A1(_270_),
    .A2(_024_),
    .ZN(_405_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _530_ (.A1(\counter[3] ),
    .A2(_413_),
    .Z(_408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _531_ (.I(\counter[0] ),
    .ZN(_330_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _532_ (.I(net2),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _533_ (.I(\counter[1] ),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _534_ (.I(net6),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _535_ (.I(net5),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _536_ (.I(net4),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _537_ (.I(net3),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _538_ (.I(_297_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _539_ (.A1(_026_),
    .A2(_256_),
    .B(_298_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _540_ (.I(_282_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _541_ (.A1(_028_),
    .A2(_250_),
    .B(_301_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _542_ (.A1(_255_),
    .A2(_292_),
    .A3(_297_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _543_ (.A1(_292_),
    .A2(_027_),
    .B1(_029_),
    .B2(_030_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _544_ (.A1(net13),
    .A2(_461_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _545_ (.A1(_287_),
    .A2(_032_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _546_ (.I(_287_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _547_ (.A1(_034_),
    .A2(_293_),
    .B(_288_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _548_ (.I(_288_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _549_ (.A1(_287_),
    .A2(_036_),
    .B(_464_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _550_ (.A1(_032_),
    .A2(_035_),
    .B1(_037_),
    .B2(_461_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _551_ (.I(_292_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _552_ (.I(_256_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _553_ (.I(_298_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _554_ (.A1(_297_),
    .A2(_040_),
    .B(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _555_ (.I(_250_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _556_ (.I(_301_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _557_ (.A1(_282_),
    .A2(_043_),
    .B(_044_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _558_ (.I(_030_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _559_ (.A1(_293_),
    .A2(_461_),
    .A3(_288_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _560_ (.A1(_039_),
    .A2(_042_),
    .B1(_045_),
    .B2(_046_),
    .C(_047_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _561_ (.A1(_031_),
    .A2(_033_),
    .B(_038_),
    .C(_048_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _562_ (.I(_049_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _563_ (.I(_366_),
    .ZN(_367_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _564_ (.I(_300_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _565_ (.A1(_028_),
    .A2(_327_),
    .B(_050_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _566_ (.A1(_255_),
    .A2(_051_),
    .B(_254_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _567_ (.I(_296_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _568_ (.A1(_026_),
    .A2(_052_),
    .B(_053_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _569_ (.A1(_292_),
    .A2(_054_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _570_ (.A1(net13),
    .A2(_286_),
    .A3(_291_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _571_ (.A1(net13),
    .A2(_287_),
    .A3(_286_),
    .B1(_055_),
    .B2(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _572_ (.A1(_461_),
    .A2(_057_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _573_ (.A1(_255_),
    .A2(_248_),
    .B(_254_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _574_ (.A1(_026_),
    .A2(_058_),
    .B(_053_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _575_ (.A1(_292_),
    .A2(_059_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _576_ (.A1(_291_),
    .A2(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _577_ (.A1(_287_),
    .A2(_061_),
    .B(_286_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _578_ (.A1(_464_),
    .A2(_062_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _579_ (.A1(_291_),
    .A2(_055_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _580_ (.A1(_287_),
    .A2(_063_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _581_ (.A1(_039_),
    .A2(_059_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _582_ (.A1(_297_),
    .A2(_052_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _583_ (.A1(_255_),
    .A2(_248_),
    .Z(_279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _584_ (.I(_255_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _585_ (.A1(_064_),
    .A2(_251_),
    .B(_256_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _586_ (.A1(_297_),
    .A2(_065_),
    .B(_041_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _587_ (.A1(_039_),
    .A2(_066_),
    .B(_293_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _588_ (.A1(_287_),
    .A2(_067_),
    .B(_036_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _589_ (.A1(_464_),
    .A2(_068_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _590_ (.A1(_293_),
    .A2(_031_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _591_ (.A1(_287_),
    .A2(_069_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _592_ (.A1(_292_),
    .A2(_066_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _593_ (.A1(_064_),
    .A2(_045_),
    .B(_256_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _594_ (.A1(_026_),
    .A2(_070_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _595_ (.A1(_255_),
    .A2(_251_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _596_ (.I(net1),
    .ZN(_437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _597_ (.I(net8),
    .ZN(_456_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _598_ (.I(net12),
    .ZN(_467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _599_ (.I(net11),
    .ZN(_470_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _600_ (.I(net10),
    .ZN(_473_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _601_ (.I(net9),
    .ZN(_476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _602_ (.I(net7),
    .ZN(_326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _603_ (.A1(\counter[6] ),
    .A2(\counter[7] ),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _604_ (.A1(net15),
    .A2(_365_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _605_ (.A1(\counter[3] ),
    .A2(\counter[2] ),
    .A3(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _606_ (.A1(\counter[5] ),
    .A2(\counter[4] ),
    .A3(_073_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _607_ (.A1(_071_),
    .A2(_074_),
    .B(net16),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _608_ (.I(_075_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _609_ (.A1(net15),
    .A2(\counter[0] ),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _610_ (.A1(_076_),
    .A2(_077_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _611_ (.I0(\counter[1] ),
    .I1(_366_),
    .S(net15),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _612_ (.A1(_076_),
    .A2(_078_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _613_ (.A1(_278_),
    .A2(_072_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _614_ (.A1(net16),
    .A2(_079_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _615_ (.A1(net15),
    .A2(\counter[0] ),
    .A3(_413_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _616_ (.A1(_274_),
    .A2(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _617_ (.A1(_076_),
    .A2(_081_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _618_ (.A1(_270_),
    .A2(_073_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _619_ (.A1(net16),
    .A2(_082_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _620_ (.A1(\counter[3] ),
    .A2(_080_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _621_ (.A1(\counter[4] ),
    .A2(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _622_ (.A1(_266_),
    .A2(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _623_ (.A1(_076_),
    .A2(_085_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _624_ (.A1(\counter[6] ),
    .A2(_074_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _625_ (.A1(net16),
    .A2(_086_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _626_ (.A1(\counter[6] ),
    .A2(\counter[5] ),
    .A3(\counter[4] ),
    .A4(_083_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _627_ (.A1(_258_),
    .A2(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _628_ (.A1(_076_),
    .A2(_088_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _629_ (.A1(_261_),
    .A2(_265_),
    .A3(_269_),
    .A4(_273_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _630_ (.A1(_284_),
    .A2(_371_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _631_ (.A1(_277_),
    .A2(_281_),
    .A3(_089_),
    .A4(_090_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _632_ (.I(_280_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _633_ (.A1(_372_),
    .A2(_284_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _634_ (.A1(_417_),
    .A2(_093_),
    .B(_281_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _635_ (.I(_277_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _636_ (.A1(_092_),
    .A2(_094_),
    .B(_095_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _637_ (.A1(_276_),
    .A2(_096_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _638_ (.I(_264_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _639_ (.A1(_272_),
    .A2(_269_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _640_ (.A1(_268_),
    .A2(_099_),
    .B(_265_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _641_ (.A1(_098_),
    .A2(_100_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _642_ (.A1(_089_),
    .A2(_097_),
    .B1(_101_),
    .B2(_261_),
    .C(_260_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _643_ (.A1(_091_),
    .A2(_102_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _644_ (.I(_341_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _645_ (.A1(_438_),
    .A2(_344_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _646_ (.A1(_345_),
    .A2(_105_),
    .B(_342_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _647_ (.A1(_340_),
    .A2(_338_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _648_ (.A1(_104_),
    .A2(_106_),
    .B(_107_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _649_ (.A1(_338_),
    .A2(_339_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _650_ (.A1(_337_),
    .A2(_108_),
    .A3(_109_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _651_ (.A1(_336_),
    .A2(_110_),
    .B(_335_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _652_ (.I(_332_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _653_ (.A1(_305_),
    .A2(_308_),
    .A3(_311_),
    .A4(_314_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _654_ (.A1(_317_),
    .A2(_323_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _655_ (.A1(_112_),
    .A2(_320_),
    .A3(_113_),
    .A4(_114_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _656_ (.I(_317_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _657_ (.I(_323_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _658_ (.I(_322_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _659_ (.A1(_117_),
    .A2(_333_),
    .B(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _660_ (.A1(_320_),
    .A2(_119_),
    .B(_319_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _661_ (.I(_316_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _662_ (.A1(_116_),
    .A2(_120_),
    .B(_121_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _663_ (.I(_307_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _664_ (.A1(_313_),
    .A2(_311_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _665_ (.A1(_310_),
    .A2(_124_),
    .B(_308_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _666_ (.A1(_123_),
    .A2(_125_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _667_ (.A1(_113_),
    .A2(_122_),
    .B1(_126_),
    .B2(_305_),
    .C(_304_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _668_ (.A1(_071_),
    .A2(_111_),
    .B1(_115_),
    .B2(_127_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _669_ (.A1(net16),
    .A2(net15),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _670_ (.A1(_103_),
    .A2(_128_),
    .B(_129_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _671_ (.A1(_381_),
    .A2(_377_),
    .A3(_379_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _672_ (.A1(_385_),
    .A2(_383_),
    .A3(_130_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _673_ (.A1(_332_),
    .A2(_375_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _674_ (.A1(_377_),
    .A2(_379_),
    .A3(_380_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _675_ (.A1(_374_),
    .A2(_376_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _676_ (.A1(_378_),
    .A2(_377_),
    .B(_133_),
    .C(_134_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _677_ (.A1(_383_),
    .A2(_384_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _678_ (.A1(_382_),
    .A2(_136_),
    .B(_130_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _679_ (.A1(_331_),
    .A2(_131_),
    .B(_135_),
    .C(_137_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _680_ (.A1(_375_),
    .A2(_374_),
    .B1(_131_),
    .B2(_132_),
    .C(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _681_ (.A1(_049_),
    .A2(_139_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _682_ (.A1(_391_),
    .A2(_389_),
    .A3(_393_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _683_ (.A1(_387_),
    .A2(_395_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _684_ (.A1(_439_),
    .A2(_141_),
    .A3(_142_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _685_ (.I(_440_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _686_ (.A1(_144_),
    .A2(_395_),
    .B(_394_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _687_ (.A1(_388_),
    .A2(_386_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _688_ (.A1(_391_),
    .A2(_392_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _689_ (.A1(_390_),
    .A2(_147_),
    .B(_389_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _690_ (.A1(_141_),
    .A2(_145_),
    .B(_146_),
    .C(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _691_ (.A1(_387_),
    .A2(_386_),
    .B(_143_),
    .C(_149_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _692_ (.A1(_020_),
    .A2(_150_),
    .B(_347_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _693_ (.A1(_347_),
    .A2(_049_),
    .A3(_139_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _694_ (.A1(_349_),
    .A2(_352_),
    .A3(_355_),
    .A4(_358_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _695_ (.A1(_371_),
    .A2(_361_),
    .A3(_364_),
    .A4(_369_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _696_ (.I(_351_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _697_ (.A1(_357_),
    .A2(_355_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _698_ (.A1(_354_),
    .A2(_156_),
    .B(_352_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _699_ (.A1(_155_),
    .A2(_157_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _700_ (.A1(_361_),
    .A2(_364_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _701_ (.I(_370_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _702_ (.A1(_369_),
    .A2(_160_),
    .B(_368_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _703_ (.A1(_361_),
    .A2(_363_),
    .B(_360_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _704_ (.A1(_159_),
    .A2(_161_),
    .B(_162_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _705_ (.A1(_349_),
    .A2(_158_),
    .B1(_163_),
    .B2(_153_),
    .C(_348_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _706_ (.A1(_153_),
    .A2(_154_),
    .B(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _707_ (.A1(_140_),
    .A2(_151_),
    .B(_152_),
    .C(_165_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _708_ (.A1(_129_),
    .A2(_166_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _709_ (.A1(_398_),
    .A2(_401_),
    .A3(_404_),
    .A4(_407_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _710_ (.I(_410_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _711_ (.I(_416_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _712_ (.A1(_371_),
    .A2(_168_),
    .A3(_418_),
    .A4(_169_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _713_ (.A1(_167_),
    .A2(_170_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _714_ (.I(_400_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _715_ (.A1(_406_),
    .A2(_404_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _716_ (.A1(_403_),
    .A2(_173_),
    .B(_401_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _717_ (.A1(_172_),
    .A2(_174_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _718_ (.I(_415_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _719_ (.A1(_372_),
    .A2(_418_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _720_ (.A1(_283_),
    .A2(_177_),
    .B(_416_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _721_ (.A1(_176_),
    .A2(_178_),
    .B(_168_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _722_ (.A1(_409_),
    .A2(_179_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _723_ (.A1(_398_),
    .A2(_175_),
    .B1(_180_),
    .B2(_167_),
    .C(_397_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _724_ (.I(_427_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _725_ (.A1(_323_),
    .A2(_333_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _726_ (.A1(_324_),
    .A2(_183_),
    .B(_428_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _727_ (.A1(_426_),
    .A2(_422_),
    .A3(_424_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _728_ (.A1(_182_),
    .A2(_184_),
    .B(_185_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _729_ (.I(_422_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _730_ (.A1(_424_),
    .A2(_425_),
    .B(_423_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _731_ (.A1(_187_),
    .A2(_188_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _732_ (.A1(_419_),
    .A2(_421_),
    .A3(_189_),
    .Z(_190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _733_ (.A1(_420_),
    .A2(_428_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _734_ (.A1(_323_),
    .A2(_332_),
    .A3(_185_),
    .A4(_191_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _735_ (.A1(_420_),
    .A2(_419_),
    .B1(_186_),
    .B2(_190_),
    .C(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _736_ (.A1(_431_),
    .A2(_430_),
    .B(_429_),
    .C(_433_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _737_ (.A1(_436_),
    .A2(_343_),
    .Z(_195_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _738_ (.I(_442_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _739_ (.A1(_344_),
    .A2(_436_),
    .A3(_196_),
    .Z(_197_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _740_ (.A1(_435_),
    .A2(_195_),
    .A3(_197_),
    .B(_434_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _741_ (.A1(_434_),
    .A2(_344_),
    .A3(_436_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _742_ (.A1(_439_),
    .A2(_430_),
    .A3(_432_),
    .A4(_199_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _743_ (.A1(_431_),
    .A2(_432_),
    .Z(_201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _744_ (.A1(_430_),
    .A2(_201_),
    .B(_429_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _745_ (.A1(_194_),
    .A2(_198_),
    .B(_200_),
    .C(_202_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _746_ (.A1(_049_),
    .A2(_193_),
    .B1(_203_),
    .B2(_399_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _747_ (.A1(_396_),
    .A2(_049_),
    .A3(_193_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _748_ (.A1(_171_),
    .A2(_181_),
    .B1(_204_),
    .B2(_396_),
    .C(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _749_ (.A1(net16),
    .A2(net15),
    .A3(_206_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _750_ (.I(_477_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _751_ (.I(_495_),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _752_ (.A1(_458_),
    .A2(_208_),
    .Z(_209_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _753_ (.A1(_457_),
    .A2(_209_),
    .B(_478_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _754_ (.A1(_207_),
    .A2(_210_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _755_ (.A1(_475_),
    .A2(_211_),
    .B(_474_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _756_ (.A1(_469_),
    .A2(_472_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _757_ (.A1(_471_),
    .A2(_469_),
    .B(_468_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _758_ (.A1(_212_),
    .A2(_213_),
    .B(_214_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _759_ (.A1(_463_),
    .A2(_466_),
    .Z(_216_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _760_ (.A1(_462_),
    .A2(_129_),
    .Z(_217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _761_ (.A1(_463_),
    .A2(_465_),
    .B1(_215_),
    .B2(_216_),
    .C(_217_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _762_ (.A1(_480_),
    .A2(_484_),
    .A3(_486_),
    .A4(_482_),
    .Z(_218_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _763_ (.A1(_494_),
    .A2(_488_),
    .A3(_490_),
    .A4(_492_),
    .Z(_219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _764_ (.I(_489_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _765_ (.I(_493_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _766_ (.A1(_492_),
    .A2(_221_),
    .Z(_222_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _767_ (.A1(_491_),
    .A2(_222_),
    .B(_490_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _768_ (.A1(_220_),
    .A2(_223_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _769_ (.A1(_488_),
    .A2(_224_),
    .Z(_225_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _770_ (.A1(_487_),
    .A2(_225_),
    .B(_218_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _771_ (.I(_481_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _772_ (.A1(_484_),
    .A2(_485_),
    .Z(_228_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _773_ (.A1(_483_),
    .A2(_228_),
    .B(_482_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _774_ (.A1(_227_),
    .A2(_229_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _775_ (.A1(_480_),
    .A2(_230_),
    .B(_479_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _776_ (.A1(_218_),
    .A2(_219_),
    .B1(_226_),
    .B2(_231_),
    .C(_129_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _777_ (.I(_454_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _778_ (.A1(_458_),
    .A2(_497_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _779_ (.A1(_459_),
    .A2(_233_),
    .B(_455_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _780_ (.A1(_232_),
    .A2(_234_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _781_ (.A1(_453_),
    .A2(_235_),
    .Z(_236_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _782_ (.A1(_445_),
    .A2(_447_),
    .A3(_449_),
    .A4(_451_),
    .Z(_237_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _783_ (.A1(_452_),
    .A2(_236_),
    .B(_237_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _784_ (.I(_446_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _785_ (.A1(_450_),
    .A2(_449_),
    .Z(_240_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _786_ (.A1(_448_),
    .A2(_240_),
    .B(_447_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _787_ (.A1(_239_),
    .A2(_241_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _788_ (.A1(_445_),
    .A2(_242_),
    .B(_444_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _789_ (.A1(_458_),
    .A2(_494_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _790_ (.A1(_453_),
    .A2(_455_),
    .A3(_237_),
    .A4(_244_),
    .Z(_245_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _791_ (.A1(_238_),
    .A2(_243_),
    .B(_129_),
    .C(_245_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _792_ (.A(_246_),
    .B(net8),
    .CI(_247_),
    .CO(_248_),
    .S(_249_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _793_ (.A(net2),
    .B(net8),
    .CI(_250_),
    .CO(_251_),
    .S(_252_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _794_ (.A(_253_),
    .B(net9),
    .CO(_254_),
    .S(_255_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _795_ (.A(net3),
    .B(net9),
    .CO(_256_),
    .S(_257_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _796_ (.A(_258_),
    .B(_259_),
    .CO(_260_),
    .S(_261_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _797_ (.A(_262_),
    .B(_263_),
    .CO(_264_),
    .S(_265_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _798_ (.A(_266_),
    .B(_267_),
    .CO(_268_),
    .S(_269_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _799_ (.A(_270_),
    .B(_271_),
    .CO(_272_),
    .S(_273_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _800_ (.A(_274_),
    .B(_275_),
    .CO(_276_),
    .S(_277_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _801_ (.A(_278_),
    .B(_279_),
    .CO(_280_),
    .S(_281_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _802_ (.A(_249_),
    .B(\counter[1] ),
    .CO(_283_),
    .S(_284_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _803_ (.A(_285_),
    .B(net12),
    .CO(_286_),
    .S(_287_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _804_ (.A(net6),
    .B(net12),
    .CO(_288_),
    .S(_289_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _805_ (.A(_290_),
    .B(net11),
    .CO(_291_),
    .S(_292_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _806_ (.A(net5),
    .B(net11),
    .CO(_293_),
    .S(_294_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _807_ (.A(_295_),
    .B(net10),
    .CO(_296_),
    .S(_297_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _808_ (.A(net4),
    .B(net10),
    .CO(_298_),
    .S(_299_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _809_ (.A(_246_),
    .B(net8),
    .CO(_300_),
    .S(_282_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _810_ (.A(net2),
    .B(net8),
    .CO(_301_),
    .S(_302_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _811_ (.A(_258_),
    .B(_303_),
    .CO(_304_),
    .S(_305_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _812_ (.A(_262_),
    .B(_306_),
    .CO(_307_),
    .S(_308_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _813_ (.A(_266_),
    .B(_309_),
    .CO(_310_),
    .S(_311_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _814_ (.A(_270_),
    .B(_312_),
    .CO(_313_),
    .S(_314_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _815_ (.A(_274_),
    .B(_315_),
    .CO(_316_),
    .S(_317_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _816_ (.A(_278_),
    .B(_318_),
    .CO(_319_),
    .S(_320_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _817_ (.A(_321_),
    .B(_252_),
    .CO(_322_),
    .S(_323_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _818_ (.A(\counter[1] ),
    .B(_252_),
    .CO(_324_),
    .S(_325_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _819_ (.A(net1),
    .B(_326_),
    .CO(_327_),
    .S(_328_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _820_ (.A(net1),
    .B(net7),
    .CO(_250_),
    .S(_329_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _821_ (.A(_330_),
    .B(_328_),
    .CO(_331_),
    .S(_332_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _822_ (.A(\counter[0] ),
    .B(_328_),
    .CO(_333_),
    .S(_334_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _823_ (.A(\counter[5] ),
    .B(net6),
    .CO(_335_),
    .S(_336_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _824_ (.A(\counter[4] ),
    .B(net5),
    .CO(_337_),
    .S(_338_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _825_ (.A(\counter[3] ),
    .B(net4),
    .CO(_339_),
    .S(_340_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _826_ (.A(\counter[2] ),
    .B(net3),
    .CO(_341_),
    .S(_342_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _827_ (.A(\counter[1] ),
    .B(_246_),
    .CO(_343_),
    .S(_344_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _828_ (.A(\counter[1] ),
    .B(net2),
    .CO(_345_),
    .S(_346_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _829_ (.A(_259_),
    .B(_347_),
    .CO(_348_),
    .S(_349_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _830_ (.A(_263_),
    .B(_350_),
    .CO(_351_),
    .S(_352_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _831_ (.A(_267_),
    .B(_353_),
    .CO(_354_),
    .S(_355_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _832_ (.A(_271_),
    .B(_356_),
    .CO(_357_),
    .S(_358_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _833_ (.A(_275_),
    .B(_359_),
    .CO(_360_),
    .S(_361_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _834_ (.A(_279_),
    .B(_362_),
    .CO(_363_),
    .S(_364_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _835_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_365_),
    .S(_366_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _836_ (.A(_249_),
    .B(_367_),
    .CO(_368_),
    .S(_369_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _837_ (.A(_330_),
    .B(_328_),
    .CO(_370_),
    .S(_371_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _838_ (.A(\counter[0] ),
    .B(_328_),
    .CO(_372_),
    .S(_373_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _839_ (.A(_306_),
    .B(_350_),
    .CO(_374_),
    .S(_375_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _840_ (.A(_309_),
    .B(_353_),
    .CO(_376_),
    .S(_377_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _841_ (.A(_312_),
    .B(_356_),
    .CO(_378_),
    .S(_379_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _842_ (.A(_315_),
    .B(_359_),
    .CO(_380_),
    .S(_381_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _843_ (.A(_318_),
    .B(_362_),
    .CO(_382_),
    .S(_383_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _844_ (.A(_252_),
    .B(_367_),
    .CO(_384_),
    .S(_385_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _845_ (.A(_285_),
    .B(_353_),
    .CO(_386_),
    .S(_387_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _846_ (.A(_290_),
    .B(_356_),
    .CO(_388_),
    .S(_389_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _847_ (.A(_295_),
    .B(_359_),
    .CO(_390_),
    .S(_391_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _848_ (.A(_253_),
    .B(_362_),
    .CO(_392_),
    .S(_393_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _849_ (.A(_246_),
    .B(_367_),
    .CO(_394_),
    .S(_395_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _850_ (.A(_396_),
    .B(_259_),
    .CO(_397_),
    .S(_398_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _851_ (.A(_399_),
    .B(_263_),
    .CO(_400_),
    .S(_401_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _852_ (.A(_402_),
    .B(_267_),
    .CO(_403_),
    .S(_404_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _853_ (.A(_405_),
    .B(_271_),
    .CO(_406_),
    .S(_407_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _854_ (.A(_408_),
    .B(_275_),
    .CO(_409_),
    .S(_410_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _855_ (.A(\counter[1] ),
    .B(_278_),
    .CO(_411_),
    .S(_412_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _856_ (.A(\counter[1] ),
    .B(\counter[2] ),
    .CO(_413_),
    .S(_414_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _857_ (.A(_412_),
    .B(_279_),
    .CO(_415_),
    .S(_416_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _858_ (.A(_321_),
    .B(_249_),
    .CO(_417_),
    .S(_418_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _859_ (.A(_399_),
    .B(_306_),
    .CO(_419_),
    .S(_420_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _860_ (.A(_402_),
    .B(_309_),
    .CO(_421_),
    .S(_422_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _861_ (.A(_405_),
    .B(_312_),
    .CO(_423_),
    .S(_424_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _862_ (.A(_408_),
    .B(_315_),
    .CO(_425_),
    .S(_426_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _863_ (.A(_412_),
    .B(_318_),
    .CO(_427_),
    .S(_428_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _864_ (.A(_285_),
    .B(_402_),
    .CO(_429_),
    .S(_430_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _865_ (.A(_290_),
    .B(_405_),
    .CO(_431_),
    .S(_432_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _866_ (.A(_295_),
    .B(_408_),
    .CO(_433_),
    .S(_434_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _867_ (.A(_253_),
    .B(_412_),
    .CO(_435_),
    .S(_436_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _868_ (.A(_330_),
    .B(_437_),
    .CO(_438_),
    .S(_439_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _869_ (.A(_330_),
    .B(net1),
    .CO(_440_),
    .S(_441_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _870_ (.A(\counter[0] ),
    .B(net1),
    .CO(_442_),
    .S(_443_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _871_ (.A(_396_),
    .B(net14),
    .CO(_444_),
    .S(_445_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _872_ (.A(_399_),
    .B(net13),
    .CO(_446_),
    .S(_447_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _873_ (.A(net12),
    .B(_402_),
    .CO(_448_),
    .S(_449_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _874_ (.A(net11),
    .B(_405_),
    .CO(_450_),
    .S(_451_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _875_ (.A(net10),
    .B(_408_),
    .CO(_452_),
    .S(_453_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _876_ (.A(net9),
    .B(_412_),
    .CO(_454_),
    .S(_455_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _877_ (.A(\counter[1] ),
    .B(_456_),
    .CO(_457_),
    .S(_458_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _878_ (.A(\counter[1] ),
    .B(net8),
    .CO(_459_),
    .S(_460_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _879_ (.A(\counter[7] ),
    .B(_461_),
    .CO(_462_),
    .S(_463_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _880_ (.A(\counter[6] ),
    .B(_464_),
    .CO(_465_),
    .S(_466_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _881_ (.A(\counter[5] ),
    .B(_467_),
    .CO(_468_),
    .S(_469_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _882_ (.A(\counter[4] ),
    .B(_470_),
    .CO(_471_),
    .S(_472_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _883_ (.A(\counter[3] ),
    .B(_473_),
    .CO(_474_),
    .S(_475_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _884_ (.A(\counter[2] ),
    .B(_476_),
    .CO(_477_),
    .S(_478_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _885_ (.A(net14),
    .B(_347_),
    .CO(_479_),
    .S(_480_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _886_ (.A(net13),
    .B(_350_),
    .CO(_481_),
    .S(_482_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _887_ (.A(net12),
    .B(_353_),
    .CO(_483_),
    .S(_484_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _888_ (.A(net11),
    .B(_356_),
    .CO(_485_),
    .S(_486_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _889_ (.A(net10),
    .B(_359_),
    .CO(_487_),
    .S(_488_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _890_ (.A(net9),
    .B(_362_),
    .CO(_489_),
    .S(_490_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _891_ (.A(net8),
    .B(_367_),
    .CO(_491_),
    .S(_492_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _892_ (.A(_330_),
    .B(_326_),
    .CO(_493_),
    .S(_494_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _893_ (.A(_330_),
    .B(net7),
    .CO(_495_),
    .S(_496_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _894_ (.A(\counter[0] ),
    .B(_326_),
    .CO(_497_),
    .S(_498_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[0]$_SDFFE_PN0P_  (.D(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[1]$_SDFFE_PN0P_  (.D(_001_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[2]$_SDFFE_PN0P_  (.D(_002_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[3]$_SDFFE_PN0P_  (.D(_003_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[4]$_SDFFE_PN0P_  (.D(_004_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[5]$_SDFFE_PN0P_  (.D(_005_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \counter[6]$_SDFFE_PN0P_  (.D(_006_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[7]$_SDFFE_PN0P_  (.D(_007_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_n_reg[0]$_SDFF_PN0_  (.D(_008_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_n_reg[1]$_SDFF_PN0_  (.D(_009_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_n_reg[2]$_SDFF_PN0_  (.D(_010_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_p_reg[0]$_SDFF_PN0_  (.D(_011_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_p_reg[1]$_SDFF_PN0_  (.D(_012_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_p_reg[2]$_SDFF_PN0_  (.D(_013_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_148 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(deadtime[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(deadtime[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(deadtime[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(deadtime[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(deadtime[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(deadtime[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(duty[0]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input8 (.I(duty[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input9 (.I(duty[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input10 (.I(duty[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input11 (.I(duty[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input12 (.I(duty[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input13 (.I(duty[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input14 (.I(duty[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input15 (.I(enable),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input16 (.I(rst_n),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net17),
    .Z(pwm_n_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net18),
    .Z(pwm_n_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net19),
    .Z(pwm_n_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net20),
    .Z(pwm_p_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net21),
    .Z(pwm_p_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net22),
    .Z(pwm_p_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_446 ();
endmodule
