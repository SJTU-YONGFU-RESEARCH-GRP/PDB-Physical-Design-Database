module clock_domain_crossing (dst_clk,
    dst_ready,
    dst_rst_n,
    dst_valid,
    src_clk,
    src_ready,
    src_rst_n,
    src_valid,
    dst_data,
    src_data);
 input dst_clk;
 input dst_ready;
 input dst_rst_n;
 output dst_valid;
 input src_clk;
 output src_ready;
 input src_rst_n;
 input src_valid;
 output [31:0] dst_data;
 input [31:0] src_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire dst_ack;
 wire dst_req_prev;
 wire \dst_req_sync[0] ;
 wire \dst_req_sync[1] ;
 wire src_ack;
 wire \src_ack_sync[0] ;
 wire \src_data_reg[0] ;
 wire \src_data_reg[10] ;
 wire \src_data_reg[11] ;
 wire \src_data_reg[12] ;
 wire \src_data_reg[13] ;
 wire \src_data_reg[14] ;
 wire \src_data_reg[15] ;
 wire \src_data_reg[16] ;
 wire \src_data_reg[17] ;
 wire \src_data_reg[18] ;
 wire \src_data_reg[19] ;
 wire \src_data_reg[1] ;
 wire \src_data_reg[20] ;
 wire \src_data_reg[21] ;
 wire \src_data_reg[22] ;
 wire \src_data_reg[23] ;
 wire \src_data_reg[24] ;
 wire \src_data_reg[25] ;
 wire \src_data_reg[26] ;
 wire \src_data_reg[27] ;
 wire \src_data_reg[28] ;
 wire \src_data_reg[29] ;
 wire \src_data_reg[2] ;
 wire \src_data_reg[30] ;
 wire \src_data_reg[31] ;
 wire \src_data_reg[3] ;
 wire \src_data_reg[4] ;
 wire \src_data_reg[5] ;
 wire \src_data_reg[6] ;
 wire \src_data_reg[7] ;
 wire \src_data_reg[8] ;
 wire \src_data_reg[9] ;
 wire src_req;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire clknet_0_src_clk;
 wire clknet_2_0__leaf_src_clk;
 wire clknet_2_1__leaf_src_clk;
 wire clknet_2_2__leaf_src_clk;
 wire clknet_2_3__leaf_src_clk;
 wire net72;
 wire net73;

 XNOR2_X2 _156_ (.A(src_req),
    .B(src_ack),
    .ZN(net71));
 INV_X1 _157_ (.A(net3),
    .ZN(_068_));
 OAI21_X1 _158_ (.A(dst_ack),
    .B1(_068_),
    .B2(\dst_req_sync[1] ),
    .ZN(_069_));
 AOI21_X1 _159_ (.A(dst_ack),
    .B1(net3),
    .B2(\dst_req_sync[1] ),
    .ZN(_070_));
 OAI21_X1 _160_ (.A(_069_),
    .B1(_070_),
    .B2(dst_req_prev),
    .ZN(_001_));
 XOR2_X2 _161_ (.A(dst_req_prev),
    .B(\dst_req_sync[1] ),
    .Z(_071_));
 BUF_X4 _162_ (.A(_071_),
    .Z(_072_));
 MUX2_X1 _163_ (.A(net38),
    .B(\src_data_reg[0] ),
    .S(_072_),
    .Z(_002_));
 MUX2_X1 _164_ (.A(net39),
    .B(\src_data_reg[10] ),
    .S(_072_),
    .Z(_003_));
 MUX2_X1 _165_ (.A(net40),
    .B(\src_data_reg[11] ),
    .S(_072_),
    .Z(_004_));
 MUX2_X1 _166_ (.A(net41),
    .B(\src_data_reg[12] ),
    .S(_072_),
    .Z(_005_));
 MUX2_X1 _167_ (.A(net42),
    .B(\src_data_reg[13] ),
    .S(_072_),
    .Z(_006_));
 MUX2_X1 _168_ (.A(net43),
    .B(\src_data_reg[14] ),
    .S(_072_),
    .Z(_007_));
 MUX2_X1 _169_ (.A(net44),
    .B(\src_data_reg[15] ),
    .S(_072_),
    .Z(_008_));
 MUX2_X1 _170_ (.A(net45),
    .B(\src_data_reg[16] ),
    .S(_072_),
    .Z(_009_));
 MUX2_X1 _171_ (.A(net46),
    .B(\src_data_reg[17] ),
    .S(_072_),
    .Z(_010_));
 BUF_X4 _172_ (.A(_071_),
    .Z(_073_));
 MUX2_X1 _173_ (.A(net47),
    .B(\src_data_reg[18] ),
    .S(_073_),
    .Z(_011_));
 MUX2_X1 _174_ (.A(net48),
    .B(\src_data_reg[19] ),
    .S(_073_),
    .Z(_012_));
 MUX2_X1 _175_ (.A(net49),
    .B(\src_data_reg[1] ),
    .S(_073_),
    .Z(_013_));
 MUX2_X1 _176_ (.A(net50),
    .B(\src_data_reg[20] ),
    .S(_073_),
    .Z(_014_));
 MUX2_X1 _177_ (.A(net51),
    .B(\src_data_reg[21] ),
    .S(_073_),
    .Z(_015_));
 MUX2_X1 _178_ (.A(net52),
    .B(\src_data_reg[22] ),
    .S(_073_),
    .Z(_016_));
 MUX2_X1 _179_ (.A(net53),
    .B(\src_data_reg[23] ),
    .S(_073_),
    .Z(_017_));
 MUX2_X1 _180_ (.A(net54),
    .B(\src_data_reg[24] ),
    .S(_073_),
    .Z(_018_));
 MUX2_X1 _181_ (.A(net55),
    .B(\src_data_reg[25] ),
    .S(_073_),
    .Z(_019_));
 MUX2_X1 _182_ (.A(net56),
    .B(\src_data_reg[26] ),
    .S(_073_),
    .Z(_020_));
 BUF_X4 _183_ (.A(_071_),
    .Z(_074_));
 MUX2_X1 _184_ (.A(net57),
    .B(\src_data_reg[27] ),
    .S(_074_),
    .Z(_021_));
 MUX2_X1 _185_ (.A(net58),
    .B(\src_data_reg[28] ),
    .S(_074_),
    .Z(_022_));
 MUX2_X1 _186_ (.A(net59),
    .B(\src_data_reg[29] ),
    .S(_074_),
    .Z(_023_));
 MUX2_X1 _187_ (.A(net60),
    .B(\src_data_reg[2] ),
    .S(_074_),
    .Z(_024_));
 MUX2_X1 _188_ (.A(net61),
    .B(\src_data_reg[30] ),
    .S(_074_),
    .Z(_025_));
 MUX2_X1 _189_ (.A(net62),
    .B(\src_data_reg[31] ),
    .S(_074_),
    .Z(_026_));
 MUX2_X1 _190_ (.A(net63),
    .B(\src_data_reg[3] ),
    .S(_074_),
    .Z(_027_));
 MUX2_X1 _191_ (.A(net64),
    .B(\src_data_reg[4] ),
    .S(_074_),
    .Z(_028_));
 MUX2_X1 _192_ (.A(net65),
    .B(\src_data_reg[5] ),
    .S(_074_),
    .Z(_029_));
 MUX2_X1 _193_ (.A(net66),
    .B(\src_data_reg[6] ),
    .S(_074_),
    .Z(_030_));
 MUX2_X1 _194_ (.A(net67),
    .B(\src_data_reg[7] ),
    .S(_071_),
    .Z(_031_));
 MUX2_X1 _195_ (.A(net68),
    .B(\src_data_reg[8] ),
    .S(_071_),
    .Z(_032_));
 MUX2_X1 _196_ (.A(net69),
    .B(\src_data_reg[9] ),
    .S(_071_),
    .Z(_033_));
 INV_X1 _197_ (.A(_072_),
    .ZN(_075_));
 INV_X1 _198_ (.A(net70),
    .ZN(_076_));
 OAI21_X1 _199_ (.A(_075_),
    .B1(_076_),
    .B2(net2),
    .ZN(_034_));
 NAND2_X4 _200_ (.A1(net37),
    .A2(net71),
    .ZN(_077_));
 BUF_X4 _201_ (.A(_077_),
    .Z(_078_));
 MUX2_X1 _202_ (.A(net4),
    .B(\src_data_reg[0] ),
    .S(_078_),
    .Z(_035_));
 MUX2_X1 _203_ (.A(net5),
    .B(\src_data_reg[10] ),
    .S(_078_),
    .Z(_036_));
 MUX2_X1 _204_ (.A(net6),
    .B(\src_data_reg[11] ),
    .S(_078_),
    .Z(_037_));
 MUX2_X1 _205_ (.A(net7),
    .B(\src_data_reg[12] ),
    .S(_078_),
    .Z(_038_));
 MUX2_X1 _206_ (.A(net8),
    .B(\src_data_reg[13] ),
    .S(_078_),
    .Z(_039_));
 MUX2_X1 _207_ (.A(net9),
    .B(\src_data_reg[14] ),
    .S(_078_),
    .Z(_040_));
 MUX2_X1 _208_ (.A(net10),
    .B(\src_data_reg[15] ),
    .S(_078_),
    .Z(_041_));
 MUX2_X1 _209_ (.A(net11),
    .B(\src_data_reg[16] ),
    .S(_078_),
    .Z(_042_));
 MUX2_X1 _210_ (.A(net12),
    .B(\src_data_reg[17] ),
    .S(_078_),
    .Z(_043_));
 MUX2_X1 _211_ (.A(net13),
    .B(\src_data_reg[18] ),
    .S(_078_),
    .Z(_044_));
 BUF_X8 _212_ (.A(_077_),
    .Z(_079_));
 MUX2_X1 _213_ (.A(net14),
    .B(\src_data_reg[19] ),
    .S(_079_),
    .Z(_045_));
 MUX2_X1 _214_ (.A(net15),
    .B(\src_data_reg[1] ),
    .S(_079_),
    .Z(_046_));
 MUX2_X1 _215_ (.A(net16),
    .B(\src_data_reg[20] ),
    .S(_079_),
    .Z(_047_));
 MUX2_X1 _216_ (.A(net17),
    .B(\src_data_reg[21] ),
    .S(_079_),
    .Z(_048_));
 MUX2_X1 _217_ (.A(net18),
    .B(\src_data_reg[22] ),
    .S(_079_),
    .Z(_049_));
 MUX2_X1 _218_ (.A(net19),
    .B(\src_data_reg[23] ),
    .S(_079_),
    .Z(_050_));
 MUX2_X1 _219_ (.A(net20),
    .B(\src_data_reg[24] ),
    .S(_079_),
    .Z(_051_));
 MUX2_X1 _220_ (.A(net21),
    .B(\src_data_reg[25] ),
    .S(_079_),
    .Z(_052_));
 MUX2_X1 _221_ (.A(net22),
    .B(\src_data_reg[26] ),
    .S(_079_),
    .Z(_053_));
 MUX2_X1 _222_ (.A(net23),
    .B(\src_data_reg[27] ),
    .S(_079_),
    .Z(_054_));
 BUF_X8 _223_ (.A(_077_),
    .Z(_080_));
 MUX2_X1 _224_ (.A(net24),
    .B(\src_data_reg[28] ),
    .S(_080_),
    .Z(_055_));
 MUX2_X1 _225_ (.A(net25),
    .B(\src_data_reg[29] ),
    .S(_080_),
    .Z(_056_));
 MUX2_X1 _226_ (.A(net26),
    .B(\src_data_reg[2] ),
    .S(_080_),
    .Z(_057_));
 MUX2_X1 _227_ (.A(net27),
    .B(\src_data_reg[30] ),
    .S(_080_),
    .Z(_058_));
 MUX2_X1 _228_ (.A(net28),
    .B(\src_data_reg[31] ),
    .S(_080_),
    .Z(_059_));
 MUX2_X1 _229_ (.A(net29),
    .B(\src_data_reg[3] ),
    .S(_080_),
    .Z(_060_));
 MUX2_X1 _230_ (.A(net30),
    .B(\src_data_reg[4] ),
    .S(_080_),
    .Z(_061_));
 MUX2_X1 _231_ (.A(net31),
    .B(\src_data_reg[5] ),
    .S(_080_),
    .Z(_062_));
 MUX2_X1 _232_ (.A(net32),
    .B(\src_data_reg[6] ),
    .S(_080_),
    .Z(_063_));
 MUX2_X1 _233_ (.A(net33),
    .B(\src_data_reg[7] ),
    .S(_080_),
    .Z(_064_));
 MUX2_X1 _234_ (.A(net34),
    .B(\src_data_reg[8] ),
    .S(_077_),
    .Z(_065_));
 MUX2_X1 _235_ (.A(net35),
    .B(\src_data_reg[9] ),
    .S(_077_),
    .Z(_066_));
 INV_X1 _236_ (.A(src_ack),
    .ZN(_081_));
 AOI21_X1 _237_ (.A(src_req),
    .B1(_081_),
    .B2(net37),
    .ZN(_082_));
 NAND2_X1 _238_ (.A1(net37),
    .A2(src_ack),
    .ZN(_083_));
 AOI21_X1 _239_ (.A(_000_),
    .B1(_083_),
    .B2(src_req),
    .ZN(_084_));
 NOR2_X1 _240_ (.A1(_082_),
    .A2(_084_),
    .ZN(_067_));
 DFF_X1 \dst_ack$_DFFE_PP_  (.D(_001_),
    .CK(net1),
    .Q(dst_ack),
    .QN(_150_));
 DFFR_X1 \dst_data[0]$_DFFE_PN0P_  (.D(_002_),
    .RN(net3),
    .CK(net1),
    .Q(net38),
    .QN(_149_));
 DFFR_X1 \dst_data[10]$_DFFE_PN0P_  (.D(_003_),
    .RN(net3),
    .CK(net1),
    .Q(net39),
    .QN(_148_));
 DFFR_X1 \dst_data[11]$_DFFE_PN0P_  (.D(_004_),
    .RN(net3),
    .CK(net1),
    .Q(net40),
    .QN(_147_));
 DFFR_X1 \dst_data[12]$_DFFE_PN0P_  (.D(_005_),
    .RN(net3),
    .CK(net1),
    .Q(net41),
    .QN(_146_));
 DFFR_X1 \dst_data[13]$_DFFE_PN0P_  (.D(_006_),
    .RN(net3),
    .CK(net1),
    .Q(net42),
    .QN(_145_));
 DFFR_X1 \dst_data[14]$_DFFE_PN0P_  (.D(_007_),
    .RN(net3),
    .CK(net1),
    .Q(net43),
    .QN(_144_));
 DFFR_X1 \dst_data[15]$_DFFE_PN0P_  (.D(_008_),
    .RN(net3),
    .CK(net1),
    .Q(net44),
    .QN(_143_));
 DFFR_X1 \dst_data[16]$_DFFE_PN0P_  (.D(_009_),
    .RN(net3),
    .CK(net1),
    .Q(net45),
    .QN(_142_));
 DFFR_X1 \dst_data[17]$_DFFE_PN0P_  (.D(_010_),
    .RN(net3),
    .CK(net1),
    .Q(net46),
    .QN(_141_));
 DFFR_X1 \dst_data[18]$_DFFE_PN0P_  (.D(_011_),
    .RN(net3),
    .CK(net1),
    .Q(net47),
    .QN(_140_));
 DFFR_X1 \dst_data[19]$_DFFE_PN0P_  (.D(_012_),
    .RN(net3),
    .CK(net1),
    .Q(net48),
    .QN(_139_));
 DFFR_X1 \dst_data[1]$_DFFE_PN0P_  (.D(_013_),
    .RN(net3),
    .CK(net1),
    .Q(net49),
    .QN(_138_));
 DFFR_X1 \dst_data[20]$_DFFE_PN0P_  (.D(_014_),
    .RN(net3),
    .CK(net1),
    .Q(net50),
    .QN(_137_));
 DFFR_X1 \dst_data[21]$_DFFE_PN0P_  (.D(_015_),
    .RN(net3),
    .CK(net1),
    .Q(net51),
    .QN(_136_));
 DFFR_X1 \dst_data[22]$_DFFE_PN0P_  (.D(_016_),
    .RN(net3),
    .CK(net1),
    .Q(net52),
    .QN(_135_));
 DFFR_X1 \dst_data[23]$_DFFE_PN0P_  (.D(_017_),
    .RN(net3),
    .CK(net1),
    .Q(net53),
    .QN(_134_));
 DFFR_X1 \dst_data[24]$_DFFE_PN0P_  (.D(_018_),
    .RN(net3),
    .CK(net1),
    .Q(net54),
    .QN(_133_));
 DFFR_X1 \dst_data[25]$_DFFE_PN0P_  (.D(_019_),
    .RN(net3),
    .CK(net1),
    .Q(net55),
    .QN(_132_));
 DFFR_X1 \dst_data[26]$_DFFE_PN0P_  (.D(_020_),
    .RN(net3),
    .CK(net1),
    .Q(net56),
    .QN(_131_));
 DFFR_X1 \dst_data[27]$_DFFE_PN0P_  (.D(_021_),
    .RN(net3),
    .CK(net1),
    .Q(net57),
    .QN(_130_));
 DFFR_X1 \dst_data[28]$_DFFE_PN0P_  (.D(_022_),
    .RN(net3),
    .CK(net1),
    .Q(net58),
    .QN(_129_));
 DFFR_X1 \dst_data[29]$_DFFE_PN0P_  (.D(_023_),
    .RN(net3),
    .CK(net1),
    .Q(net59),
    .QN(_128_));
 DFFR_X1 \dst_data[2]$_DFFE_PN0P_  (.D(_024_),
    .RN(net3),
    .CK(net1),
    .Q(net60),
    .QN(_127_));
 DFFR_X1 \dst_data[30]$_DFFE_PN0P_  (.D(_025_),
    .RN(net3),
    .CK(net1),
    .Q(net61),
    .QN(_126_));
 DFFR_X1 \dst_data[31]$_DFFE_PN0P_  (.D(_026_),
    .RN(net3),
    .CK(net1),
    .Q(net62),
    .QN(_125_));
 DFFR_X1 \dst_data[3]$_DFFE_PN0P_  (.D(_027_),
    .RN(net3),
    .CK(net1),
    .Q(net63),
    .QN(_124_));
 DFFR_X1 \dst_data[4]$_DFFE_PN0P_  (.D(_028_),
    .RN(net3),
    .CK(net1),
    .Q(net64),
    .QN(_123_));
 DFFR_X1 \dst_data[5]$_DFFE_PN0P_  (.D(_029_),
    .RN(net3),
    .CK(net1),
    .Q(net65),
    .QN(_122_));
 DFFR_X1 \dst_data[6]$_DFFE_PN0P_  (.D(_030_),
    .RN(net3),
    .CK(net1),
    .Q(net66),
    .QN(_121_));
 DFFR_X1 \dst_data[7]$_DFFE_PN0P_  (.D(_031_),
    .RN(net3),
    .CK(net1),
    .Q(net67),
    .QN(_120_));
 DFFR_X1 \dst_data[8]$_DFFE_PN0P_  (.D(_032_),
    .RN(net3),
    .CK(net1),
    .Q(net68),
    .QN(_119_));
 DFFR_X1 \dst_data[9]$_DFFE_PN0P_  (.D(_033_),
    .RN(net3),
    .CK(net1),
    .Q(net69),
    .QN(_151_));
 DFFR_X1 \dst_req_prev$_DFF_PN0_  (.D(\dst_req_sync[1] ),
    .RN(net3),
    .CK(net1),
    .Q(dst_req_prev),
    .QN(_152_));
 DFFR_X1 \dst_req_sync[0]$_DFF_PN0_  (.D(src_req),
    .RN(net3),
    .CK(net1),
    .Q(\dst_req_sync[0] ),
    .QN(_153_));
 DFFR_X2 \dst_req_sync[1]$_DFF_PN0_  (.D(\dst_req_sync[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\dst_req_sync[1] ),
    .QN(_118_));
 DFFR_X1 \dst_valid$_DFFE_PN0P_  (.D(_034_),
    .RN(net3),
    .CK(net1),
    .Q(net70),
    .QN(_154_));
 DFFR_X1 \src_ack_sync[0]$_DFF_PN0_  (.D(dst_ack),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\src_ack_sync[0] ),
    .QN(_155_));
 DFFR_X1 \src_ack_sync[1]$_DFF_PN0_  (.D(\src_ack_sync[0] ),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(src_ack),
    .QN(_117_));
 DFFR_X1 \src_data_reg[0]$_DFFE_PN0P_  (.D(_035_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[0] ),
    .QN(_116_));
 DFFR_X1 \src_data_reg[10]$_DFFE_PN0P_  (.D(_036_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[10] ),
    .QN(_115_));
 DFFR_X1 \src_data_reg[11]$_DFFE_PN0P_  (.D(_037_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[11] ),
    .QN(_114_));
 DFFR_X1 \src_data_reg[12]$_DFFE_PN0P_  (.D(_038_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[12] ),
    .QN(_113_));
 DFFR_X1 \src_data_reg[13]$_DFFE_PN0P_  (.D(_039_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[13] ),
    .QN(_112_));
 DFFR_X1 \src_data_reg[14]$_DFFE_PN0P_  (.D(_040_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[14] ),
    .QN(_111_));
 DFFR_X1 \src_data_reg[15]$_DFFE_PN0P_  (.D(_041_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[15] ),
    .QN(_110_));
 DFFR_X1 \src_data_reg[16]$_DFFE_PN0P_  (.D(_042_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[16] ),
    .QN(_109_));
 DFFR_X1 \src_data_reg[17]$_DFFE_PN0P_  (.D(_043_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[17] ),
    .QN(_108_));
 DFFR_X1 \src_data_reg[18]$_DFFE_PN0P_  (.D(_044_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[18] ),
    .QN(_107_));
 DFFR_X1 \src_data_reg[19]$_DFFE_PN0P_  (.D(_045_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[19] ),
    .QN(_106_));
 DFFR_X1 \src_data_reg[1]$_DFFE_PN0P_  (.D(_046_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[1] ),
    .QN(_105_));
 DFFR_X1 \src_data_reg[20]$_DFFE_PN0P_  (.D(_047_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[20] ),
    .QN(_104_));
 DFFR_X1 \src_data_reg[21]$_DFFE_PN0P_  (.D(_048_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[21] ),
    .QN(_103_));
 DFFR_X1 \src_data_reg[22]$_DFFE_PN0P_  (.D(_049_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[22] ),
    .QN(_102_));
 DFFR_X1 \src_data_reg[23]$_DFFE_PN0P_  (.D(_050_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[23] ),
    .QN(_101_));
 DFFR_X1 \src_data_reg[24]$_DFFE_PN0P_  (.D(_051_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[24] ),
    .QN(_100_));
 DFFR_X1 \src_data_reg[25]$_DFFE_PN0P_  (.D(_052_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[25] ),
    .QN(_099_));
 DFFR_X1 \src_data_reg[26]$_DFFE_PN0P_  (.D(_053_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[26] ),
    .QN(_098_));
 DFFR_X1 \src_data_reg[27]$_DFFE_PN0P_  (.D(_054_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[27] ),
    .QN(_097_));
 DFFR_X1 \src_data_reg[28]$_DFFE_PN0P_  (.D(_055_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[28] ),
    .QN(_096_));
 DFFR_X1 \src_data_reg[29]$_DFFE_PN0P_  (.D(_056_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[29] ),
    .QN(_095_));
 DFFR_X1 \src_data_reg[2]$_DFFE_PN0P_  (.D(_057_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[2] ),
    .QN(_094_));
 DFFR_X1 \src_data_reg[30]$_DFFE_PN0P_  (.D(_058_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[30] ),
    .QN(_093_));
 DFFR_X1 \src_data_reg[31]$_DFFE_PN0P_  (.D(_059_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[31] ),
    .QN(_092_));
 DFFR_X1 \src_data_reg[3]$_DFFE_PN0P_  (.D(_060_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[3] ),
    .QN(_091_));
 DFFR_X1 \src_data_reg[4]$_DFFE_PN0P_  (.D(_061_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[4] ),
    .QN(_090_));
 DFFR_X1 \src_data_reg[5]$_DFFE_PN0P_  (.D(_062_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[5] ),
    .QN(_089_));
 DFFR_X1 \src_data_reg[6]$_DFFE_PN0P_  (.D(_063_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[6] ),
    .QN(_088_));
 DFFR_X1 \src_data_reg[7]$_DFFE_PN0P_  (.D(_064_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[7] ),
    .QN(_087_));
 DFFR_X1 \src_data_reg[8]$_DFFE_PN0P_  (.D(_065_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[8] ),
    .QN(_086_));
 DFFR_X1 \src_data_reg[9]$_DFFE_PN0P_  (.D(_066_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[9] ),
    .QN(_085_));
 DFFR_X1 \src_req$_DFFE_PN0P_  (.D(_067_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(src_req),
    .QN(_000_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_45 ();
 BUF_X8 input1 (.A(dst_clk),
    .Z(net1));
 BUF_X1 input2 (.A(dst_ready),
    .Z(net2));
 BUF_X8 input3 (.A(dst_rst_n),
    .Z(net3));
 BUF_X1 input4 (.A(src_data[0]),
    .Z(net4));
 BUF_X1 input5 (.A(src_data[10]),
    .Z(net5));
 BUF_X1 input6 (.A(src_data[11]),
    .Z(net6));
 BUF_X1 input7 (.A(src_data[12]),
    .Z(net7));
 BUF_X1 input8 (.A(src_data[13]),
    .Z(net8));
 BUF_X1 input9 (.A(src_data[14]),
    .Z(net9));
 BUF_X1 input10 (.A(src_data[15]),
    .Z(net10));
 BUF_X1 input11 (.A(src_data[16]),
    .Z(net11));
 BUF_X1 input12 (.A(src_data[17]),
    .Z(net12));
 BUF_X1 input13 (.A(src_data[18]),
    .Z(net13));
 BUF_X1 input14 (.A(src_data[19]),
    .Z(net14));
 BUF_X1 input15 (.A(src_data[1]),
    .Z(net15));
 BUF_X1 input16 (.A(src_data[20]),
    .Z(net16));
 BUF_X1 input17 (.A(src_data[21]),
    .Z(net17));
 BUF_X1 input18 (.A(src_data[22]),
    .Z(net18));
 BUF_X1 input19 (.A(src_data[23]),
    .Z(net19));
 BUF_X1 input20 (.A(src_data[24]),
    .Z(net20));
 BUF_X1 input21 (.A(src_data[25]),
    .Z(net21));
 BUF_X1 input22 (.A(src_data[26]),
    .Z(net22));
 BUF_X1 input23 (.A(src_data[27]),
    .Z(net23));
 BUF_X1 input24 (.A(src_data[28]),
    .Z(net24));
 BUF_X1 input25 (.A(src_data[29]),
    .Z(net25));
 BUF_X1 input26 (.A(src_data[2]),
    .Z(net26));
 BUF_X1 input27 (.A(src_data[30]),
    .Z(net27));
 BUF_X1 input28 (.A(src_data[31]),
    .Z(net28));
 BUF_X1 input29 (.A(src_data[3]),
    .Z(net29));
 BUF_X1 input30 (.A(src_data[4]),
    .Z(net30));
 BUF_X1 input31 (.A(src_data[5]),
    .Z(net31));
 BUF_X1 input32 (.A(src_data[6]),
    .Z(net32));
 BUF_X1 input33 (.A(src_data[7]),
    .Z(net33));
 BUF_X1 input34 (.A(src_data[8]),
    .Z(net34));
 BUF_X1 input35 (.A(src_data[9]),
    .Z(net35));
 BUF_X8 input36 (.A(net72),
    .Z(net36));
 BUF_X1 input37 (.A(src_valid),
    .Z(net37));
 BUF_X1 output38 (.A(net38),
    .Z(dst_data[0]));
 BUF_X1 output39 (.A(net39),
    .Z(dst_data[10]));
 BUF_X1 output40 (.A(net40),
    .Z(dst_data[11]));
 BUF_X1 output41 (.A(net41),
    .Z(dst_data[12]));
 BUF_X1 output42 (.A(net42),
    .Z(dst_data[13]));
 BUF_X1 output43 (.A(net43),
    .Z(dst_data[14]));
 BUF_X1 output44 (.A(net44),
    .Z(dst_data[15]));
 BUF_X1 output45 (.A(net45),
    .Z(dst_data[16]));
 BUF_X1 output46 (.A(net46),
    .Z(dst_data[17]));
 BUF_X1 output47 (.A(net47),
    .Z(dst_data[18]));
 BUF_X1 output48 (.A(net48),
    .Z(dst_data[19]));
 BUF_X1 output49 (.A(net49),
    .Z(dst_data[1]));
 BUF_X1 output50 (.A(net50),
    .Z(dst_data[20]));
 BUF_X1 output51 (.A(net51),
    .Z(dst_data[21]));
 BUF_X1 output52 (.A(net52),
    .Z(dst_data[22]));
 BUF_X1 output53 (.A(net53),
    .Z(dst_data[23]));
 BUF_X1 output54 (.A(net54),
    .Z(dst_data[24]));
 BUF_X1 output55 (.A(net55),
    .Z(dst_data[25]));
 BUF_X1 output56 (.A(net56),
    .Z(dst_data[26]));
 BUF_X1 output57 (.A(net57),
    .Z(dst_data[27]));
 BUF_X1 output58 (.A(net58),
    .Z(dst_data[28]));
 BUF_X1 output59 (.A(net59),
    .Z(dst_data[29]));
 BUF_X1 output60 (.A(net60),
    .Z(dst_data[2]));
 BUF_X1 output61 (.A(net61),
    .Z(dst_data[30]));
 BUF_X1 output62 (.A(net62),
    .Z(dst_data[31]));
 BUF_X1 output63 (.A(net63),
    .Z(dst_data[3]));
 BUF_X1 output64 (.A(net64),
    .Z(dst_data[4]));
 BUF_X1 output65 (.A(net65),
    .Z(dst_data[5]));
 BUF_X1 output66 (.A(net66),
    .Z(dst_data[6]));
 BUF_X1 output67 (.A(net67),
    .Z(dst_data[7]));
 BUF_X1 output68 (.A(net68),
    .Z(dst_data[8]));
 BUF_X1 output69 (.A(net69),
    .Z(dst_data[9]));
 BUF_X1 output70 (.A(net70),
    .Z(dst_valid));
 BUF_X1 output71 (.A(net71),
    .Z(src_ready));
 CLKBUF_X3 clkbuf_0_src_clk (.A(src_clk),
    .Z(clknet_0_src_clk));
 CLKBUF_X3 clkbuf_2_0__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_0__leaf_src_clk));
 CLKBUF_X3 clkbuf_2_1__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_1__leaf_src_clk));
 CLKBUF_X3 clkbuf_2_2__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_2__leaf_src_clk));
 CLKBUF_X3 clkbuf_2_3__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_3__leaf_src_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_src_clk));
 INV_X1 clkload1 (.A(clknet_2_2__leaf_src_clk));
 CLKBUF_X1 hold1 (.A(src_rst_n),
    .Z(net72));
 BUF_X8 hold2 (.A(net36),
    .Z(net73));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_17 ();
 FILLCELL_X2 FILLER_0_25 ();
 FILLCELL_X2 FILLER_0_30 ();
 FILLCELL_X1 FILLER_0_32 ();
 FILLCELL_X8 FILLER_0_36 ();
 FILLCELL_X1 FILLER_0_44 ();
 FILLCELL_X2 FILLER_0_48 ();
 FILLCELL_X4 FILLER_0_53 ();
 FILLCELL_X2 FILLER_0_57 ();
 FILLCELL_X1 FILLER_0_59 ();
 FILLCELL_X2 FILLER_0_69 ();
 FILLCELL_X1 FILLER_0_71 ();
 FILLCELL_X4 FILLER_0_75 ();
 FILLCELL_X2 FILLER_0_79 ();
 FILLCELL_X4 FILLER_0_84 ();
 FILLCELL_X1 FILLER_0_88 ();
 FILLCELL_X2 FILLER_0_108 ();
 FILLCELL_X1 FILLER_0_110 ();
 FILLCELL_X8 FILLER_0_124 ();
 FILLCELL_X1 FILLER_0_135 ();
 FILLCELL_X4 FILLER_0_139 ();
 FILLCELL_X2 FILLER_0_143 ();
 FILLCELL_X4 FILLER_0_165 ();
 FILLCELL_X8 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_9 ();
 FILLCELL_X1 FILLER_1_11 ();
 FILLCELL_X2 FILLER_1_39 ();
 FILLCELL_X16 FILLER_1_68 ();
 FILLCELL_X4 FILLER_1_84 ();
 FILLCELL_X1 FILLER_1_88 ();
 FILLCELL_X1 FILLER_1_109 ();
 FILLCELL_X4 FILLER_1_130 ();
 FILLCELL_X2 FILLER_1_134 ();
 FILLCELL_X1 FILLER_1_136 ();
 FILLCELL_X2 FILLER_1_144 ();
 FILLCELL_X1 FILLER_1_146 ();
 FILLCELL_X2 FILLER_1_167 ();
 FILLCELL_X8 FILLER_2_1 ();
 FILLCELL_X2 FILLER_2_9 ();
 FILLCELL_X4 FILLER_2_38 ();
 FILLCELL_X2 FILLER_2_42 ();
 FILLCELL_X1 FILLER_2_78 ();
 FILLCELL_X2 FILLER_2_140 ();
 FILLCELL_X2 FILLER_2_149 ();
 FILLCELL_X8 FILLER_2_158 ();
 FILLCELL_X4 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_45 ();
 FILLCELL_X4 FILLER_3_53 ();
 FILLCELL_X2 FILLER_3_77 ();
 FILLCELL_X1 FILLER_3_93 ();
 FILLCELL_X1 FILLER_3_114 ();
 FILLCELL_X1 FILLER_3_122 ();
 FILLCELL_X2 FILLER_3_143 ();
 FILLCELL_X1 FILLER_3_165 ();
 FILLCELL_X2 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_17 ();
 FILLCELL_X8 FILLER_4_33 ();
 FILLCELL_X2 FILLER_4_41 ();
 FILLCELL_X32 FILLER_4_103 ();
 FILLCELL_X32 FILLER_4_135 ();
 FILLCELL_X2 FILLER_4_167 ();
 FILLCELL_X2 FILLER_5_1 ();
 FILLCELL_X2 FILLER_5_6 ();
 FILLCELL_X1 FILLER_5_8 ();
 FILLCELL_X1 FILLER_5_12 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_49 ();
 FILLCELL_X4 FILLER_5_57 ();
 FILLCELL_X2 FILLER_5_61 ();
 FILLCELL_X1 FILLER_5_63 ();
 FILLCELL_X32 FILLER_5_71 ();
 FILLCELL_X1 FILLER_5_103 ();
 FILLCELL_X16 FILLER_5_109 ();
 FILLCELL_X8 FILLER_5_125 ();
 FILLCELL_X4 FILLER_5_133 ();
 FILLCELL_X1 FILLER_5_137 ();
 FILLCELL_X4 FILLER_5_165 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_9 ();
 FILLCELL_X1 FILLER_6_13 ();
 FILLCELL_X4 FILLER_6_34 ();
 FILLCELL_X2 FILLER_6_38 ();
 FILLCELL_X32 FILLER_6_48 ();
 FILLCELL_X8 FILLER_6_80 ();
 FILLCELL_X4 FILLER_6_88 ();
 FILLCELL_X2 FILLER_6_92 ();
 FILLCELL_X1 FILLER_6_94 ();
 FILLCELL_X8 FILLER_6_102 ();
 FILLCELL_X4 FILLER_6_110 ();
 FILLCELL_X2 FILLER_6_114 ();
 FILLCELL_X1 FILLER_6_116 ();
 FILLCELL_X2 FILLER_6_144 ();
 FILLCELL_X8 FILLER_6_156 ();
 FILLCELL_X2 FILLER_6_164 ();
 FILLCELL_X2 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_3 ();
 FILLCELL_X4 FILLER_7_7 ();
 FILLCELL_X1 FILLER_7_18 ();
 FILLCELL_X32 FILLER_7_39 ();
 FILLCELL_X16 FILLER_7_71 ();
 FILLCELL_X4 FILLER_7_87 ();
 FILLCELL_X1 FILLER_7_91 ();
 FILLCELL_X8 FILLER_7_112 ();
 FILLCELL_X4 FILLER_7_120 ();
 FILLCELL_X2 FILLER_7_124 ();
 FILLCELL_X1 FILLER_7_126 ();
 FILLCELL_X2 FILLER_7_167 ();
 FILLCELL_X2 FILLER_8_14 ();
 FILLCELL_X4 FILLER_8_23 ();
 FILLCELL_X32 FILLER_8_47 ();
 FILLCELL_X8 FILLER_8_79 ();
 FILLCELL_X4 FILLER_8_87 ();
 FILLCELL_X2 FILLER_8_91 ();
 FILLCELL_X1 FILLER_8_93 ();
 FILLCELL_X8 FILLER_8_121 ();
 FILLCELL_X2 FILLER_8_129 ();
 FILLCELL_X4 FILLER_8_155 ();
 FILLCELL_X1 FILLER_8_159 ();
 FILLCELL_X32 FILLER_9_38 ();
 FILLCELL_X32 FILLER_9_70 ();
 FILLCELL_X16 FILLER_9_102 ();
 FILLCELL_X8 FILLER_9_118 ();
 FILLCELL_X2 FILLER_9_126 ();
 FILLCELL_X1 FILLER_9_168 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_3 ();
 FILLCELL_X32 FILLER_10_50 ();
 FILLCELL_X32 FILLER_10_82 ();
 FILLCELL_X16 FILLER_10_114 ();
 FILLCELL_X8 FILLER_10_130 ();
 FILLCELL_X4 FILLER_10_138 ();
 FILLCELL_X1 FILLER_10_142 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_5 ();
 FILLCELL_X8 FILLER_11_10 ();
 FILLCELL_X4 FILLER_11_18 ();
 FILLCELL_X1 FILLER_11_22 ();
 FILLCELL_X16 FILLER_11_30 ();
 FILLCELL_X8 FILLER_11_46 ();
 FILLCELL_X4 FILLER_11_54 ();
 FILLCELL_X1 FILLER_11_58 ();
 FILLCELL_X8 FILLER_11_66 ();
 FILLCELL_X1 FILLER_11_74 ();
 FILLCELL_X32 FILLER_11_87 ();
 FILLCELL_X8 FILLER_11_119 ();
 FILLCELL_X4 FILLER_11_127 ();
 FILLCELL_X2 FILLER_11_131 ();
 FILLCELL_X1 FILLER_11_140 ();
 FILLCELL_X4 FILLER_11_148 ();
 FILLCELL_X1 FILLER_11_152 ();
 FILLCELL_X8 FILLER_11_156 ();
 FILLCELL_X4 FILLER_11_164 ();
 FILLCELL_X1 FILLER_11_168 ();
 FILLCELL_X1 FILLER_12_4 ();
 FILLCELL_X2 FILLER_12_19 ();
 FILLCELL_X1 FILLER_12_21 ();
 FILLCELL_X2 FILLER_12_42 ();
 FILLCELL_X1 FILLER_12_44 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X4 FILLER_12_121 ();
 FILLCELL_X1 FILLER_12_125 ();
 FILLCELL_X4 FILLER_12_153 ();
 FILLCELL_X2 FILLER_12_157 ();
 FILLCELL_X1 FILLER_12_159 ();
 FILLCELL_X4 FILLER_12_163 ();
 FILLCELL_X2 FILLER_12_167 ();
 FILLCELL_X4 FILLER_13_7 ();
 FILLCELL_X1 FILLER_13_11 ();
 FILLCELL_X2 FILLER_13_39 ();
 FILLCELL_X1 FILLER_13_41 ();
 FILLCELL_X2 FILLER_13_49 ();
 FILLCELL_X1 FILLER_13_51 ();
 FILLCELL_X8 FILLER_13_59 ();
 FILLCELL_X4 FILLER_13_67 ();
 FILLCELL_X2 FILLER_13_71 ();
 FILLCELL_X16 FILLER_13_106 ();
 FILLCELL_X4 FILLER_13_122 ();
 FILLCELL_X2 FILLER_13_126 ();
 FILLCELL_X8 FILLER_13_158 ();
 FILLCELL_X2 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_3 ();
 FILLCELL_X4 FILLER_14_34 ();
 FILLCELL_X1 FILLER_14_74 ();
 FILLCELL_X8 FILLER_14_82 ();
 FILLCELL_X2 FILLER_14_90 ();
 FILLCELL_X8 FILLER_14_112 ();
 FILLCELL_X4 FILLER_14_120 ();
 FILLCELL_X2 FILLER_14_124 ();
 FILLCELL_X1 FILLER_14_126 ();
 FILLCELL_X2 FILLER_14_167 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_5 ();
 FILLCELL_X1 FILLER_15_7 ();
 FILLCELL_X16 FILLER_15_28 ();
 FILLCELL_X2 FILLER_15_44 ();
 FILLCELL_X1 FILLER_15_46 ();
 FILLCELL_X16 FILLER_15_64 ();
 FILLCELL_X2 FILLER_15_80 ();
 FILLCELL_X1 FILLER_15_82 ();
 FILLCELL_X16 FILLER_15_117 ();
 FILLCELL_X2 FILLER_15_133 ();
 FILLCELL_X2 FILLER_15_142 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X1 FILLER_15_165 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X8 FILLER_16_33 ();
 FILLCELL_X2 FILLER_16_41 ();
 FILLCELL_X1 FILLER_16_43 ();
 FILLCELL_X8 FILLER_16_70 ();
 FILLCELL_X2 FILLER_16_78 ();
 FILLCELL_X1 FILLER_16_101 ();
 FILLCELL_X8 FILLER_16_122 ();
 FILLCELL_X4 FILLER_16_130 ();
 FILLCELL_X1 FILLER_16_168 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X16 FILLER_17_8 ();
 FILLCELL_X1 FILLER_17_24 ();
 FILLCELL_X2 FILLER_17_45 ();
 FILLCELL_X1 FILLER_17_61 ();
 FILLCELL_X32 FILLER_17_70 ();
 FILLCELL_X8 FILLER_17_102 ();
 FILLCELL_X1 FILLER_17_110 ();
 FILLCELL_X16 FILLER_17_116 ();
 FILLCELL_X4 FILLER_17_132 ();
 FILLCELL_X2 FILLER_17_136 ();
 FILLCELL_X1 FILLER_17_165 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_3 ();
 FILLCELL_X4 FILLER_18_16 ();
 FILLCELL_X1 FILLER_18_20 ();
 FILLCELL_X8 FILLER_18_48 ();
 FILLCELL_X4 FILLER_18_58 ();
 FILLCELL_X1 FILLER_18_62 ();
 FILLCELL_X32 FILLER_18_70 ();
 FILLCELL_X32 FILLER_18_102 ();
 FILLCELL_X32 FILLER_18_134 ();
 FILLCELL_X1 FILLER_19_34 ();
 FILLCELL_X1 FILLER_19_55 ();
 FILLCELL_X1 FILLER_19_76 ();
 FILLCELL_X1 FILLER_19_83 ();
 FILLCELL_X1 FILLER_19_106 ();
 FILLCELL_X8 FILLER_19_154 ();
 FILLCELL_X4 FILLER_19_162 ();
 FILLCELL_X2 FILLER_19_166 ();
 FILLCELL_X1 FILLER_19_168 ();
 FILLCELL_X1 FILLER_20_4 ();
 FILLCELL_X4 FILLER_20_33 ();
 FILLCELL_X4 FILLER_20_164 ();
 FILLCELL_X1 FILLER_20_168 ();
 FILLCELL_X8 FILLER_21_34 ();
 FILLCELL_X4 FILLER_21_42 ();
 FILLCELL_X1 FILLER_21_49 ();
 FILLCELL_X2 FILLER_21_57 ();
 FILLCELL_X1 FILLER_21_59 ();
 FILLCELL_X4 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_74 ();
 FILLCELL_X2 FILLER_21_78 ();
 FILLCELL_X1 FILLER_21_80 ();
 FILLCELL_X1 FILLER_21_98 ();
 FILLCELL_X1 FILLER_21_109 ();
 FILLCELL_X2 FILLER_21_117 ();
 FILLCELL_X1 FILLER_21_126 ();
 FILLCELL_X2 FILLER_21_134 ();
 FILLCELL_X2 FILLER_21_143 ();
 FILLCELL_X4 FILLER_21_165 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_9 ();
 FILLCELL_X4 FILLER_22_39 ();
 FILLCELL_X2 FILLER_22_66 ();
 FILLCELL_X8 FILLER_22_71 ();
 FILLCELL_X4 FILLER_22_79 ();
 FILLCELL_X2 FILLER_22_86 ();
 FILLCELL_X1 FILLER_22_88 ();
 FILLCELL_X2 FILLER_22_92 ();
 FILLCELL_X1 FILLER_22_94 ();
 FILLCELL_X2 FILLER_22_104 ();
 FILLCELL_X1 FILLER_22_106 ();
 FILLCELL_X2 FILLER_22_110 ();
 FILLCELL_X2 FILLER_22_115 ();
 FILLCELL_X1 FILLER_22_117 ();
 FILLCELL_X4 FILLER_22_121 ();
 FILLCELL_X2 FILLER_22_125 ();
 FILLCELL_X2 FILLER_22_130 ();
 FILLCELL_X1 FILLER_22_132 ();
 FILLCELL_X8 FILLER_22_136 ();
 FILLCELL_X4 FILLER_22_144 ();
 FILLCELL_X2 FILLER_22_151 ();
 FILLCELL_X1 FILLER_22_153 ();
 FILLCELL_X2 FILLER_22_167 ();
endmodule
