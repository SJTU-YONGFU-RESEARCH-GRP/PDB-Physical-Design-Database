module configurable_lfsr (clk,
    enable,
    load_seed,
    rst_n,
    serial_out,
    parallel_out,
    seed,
    tap_pattern);
 input clk;
 input enable;
 input load_seed;
 input rst_n;
 output serial_out;
 output [7:0] parallel_out;
 input [7:0] seed;
 input [7:0] tap_pattern;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net28;

 sky130_fd_sc_hd__buf_2 _42_ (.A(net2),
    .X(_08_));
 sky130_fd_sc_hd__clkbuf_4 _43_ (.A(enable),
    .X(_09_));
 sky130_fd_sc_hd__mux2i_1 _44_ (.A0(net27),
    .A1(net20),
    .S(_09_),
    .Y(_10_));
 sky130_fd_sc_hd__nand2_1 _45_ (.A(_08_),
    .B(net3),
    .Y(_11_));
 sky130_fd_sc_hd__o21ai_0 _46_ (.A1(_08_),
    .A2(_10_),
    .B1(_11_),
    .Y(_00_));
 sky130_fd_sc_hd__mux2i_1 _47_ (.A0(net20),
    .A1(net21),
    .S(_09_),
    .Y(_12_));
 sky130_fd_sc_hd__nand2_1 _48_ (.A(_08_),
    .B(net4),
    .Y(_13_));
 sky130_fd_sc_hd__o21ai_0 _49_ (.A1(_08_),
    .A2(_12_),
    .B1(_13_),
    .Y(_01_));
 sky130_fd_sc_hd__mux2i_1 _50_ (.A0(net21),
    .A1(net22),
    .S(_09_),
    .Y(_14_));
 sky130_fd_sc_hd__nand2_1 _51_ (.A(_08_),
    .B(net5),
    .Y(_15_));
 sky130_fd_sc_hd__o21ai_0 _52_ (.A1(_08_),
    .A2(_14_),
    .B1(_15_),
    .Y(_02_));
 sky130_fd_sc_hd__mux2i_1 _53_ (.A0(net22),
    .A1(net23),
    .S(_09_),
    .Y(_16_));
 sky130_fd_sc_hd__nand2_1 _54_ (.A(_08_),
    .B(net6),
    .Y(_17_));
 sky130_fd_sc_hd__o21ai_0 _55_ (.A1(net2),
    .A2(_16_),
    .B1(_17_),
    .Y(_03_));
 sky130_fd_sc_hd__mux2i_1 _56_ (.A0(net23),
    .A1(net24),
    .S(_09_),
    .Y(_18_));
 sky130_fd_sc_hd__nand2_1 _57_ (.A(_08_),
    .B(net7),
    .Y(_19_));
 sky130_fd_sc_hd__o21ai_0 _58_ (.A1(net2),
    .A2(_18_),
    .B1(_19_),
    .Y(_04_));
 sky130_fd_sc_hd__mux2i_1 _59_ (.A0(net24),
    .A1(net25),
    .S(_09_),
    .Y(_20_));
 sky130_fd_sc_hd__nand2_1 _60_ (.A(_08_),
    .B(net8),
    .Y(_21_));
 sky130_fd_sc_hd__o21ai_0 _61_ (.A1(net2),
    .A2(_20_),
    .B1(_21_),
    .Y(_05_));
 sky130_fd_sc_hd__mux2i_1 _62_ (.A0(net25),
    .A1(net26),
    .S(_09_),
    .Y(_22_));
 sky130_fd_sc_hd__nand2_1 _63_ (.A(_08_),
    .B(net9),
    .Y(_23_));
 sky130_fd_sc_hd__o21ai_0 _64_ (.A1(net2),
    .A2(_22_),
    .B1(_23_),
    .Y(_06_));
 sky130_fd_sc_hd__nand2_1 _65_ (.A(net24),
    .B(net16),
    .Y(_24_));
 sky130_fd_sc_hd__nand2_1 _66_ (.A(net22),
    .B(net14),
    .Y(_25_));
 sky130_fd_sc_hd__xor2_1 _67_ (.A(_24_),
    .B(_25_),
    .X(_26_));
 sky130_fd_sc_hd__nand2_1 _68_ (.A(net25),
    .B(net17),
    .Y(_27_));
 sky130_fd_sc_hd__nand2_1 _69_ (.A(net23),
    .B(net15),
    .Y(_28_));
 sky130_fd_sc_hd__xnor2_1 _70_ (.A(_27_),
    .B(_28_),
    .Y(_29_));
 sky130_fd_sc_hd__xnor2_1 _71_ (.A(_26_),
    .B(_29_),
    .Y(_30_));
 sky130_fd_sc_hd__nand2_1 _72_ (.A(net20),
    .B(net12),
    .Y(_31_));
 sky130_fd_sc_hd__nand2_1 _73_ (.A(net11),
    .B(net27),
    .Y(_32_));
 sky130_fd_sc_hd__xor2_1 _74_ (.A(_31_),
    .B(_32_),
    .X(_33_));
 sky130_fd_sc_hd__nand2_1 _75_ (.A(net26),
    .B(net18),
    .Y(_34_));
 sky130_fd_sc_hd__nand2_1 _76_ (.A(net21),
    .B(net13),
    .Y(_35_));
 sky130_fd_sc_hd__xnor2_1 _77_ (.A(_34_),
    .B(_35_),
    .Y(_36_));
 sky130_fd_sc_hd__xnor2_1 _78_ (.A(_33_),
    .B(_36_),
    .Y(_37_));
 sky130_fd_sc_hd__xnor2_1 _79_ (.A(_30_),
    .B(_37_),
    .Y(_38_));
 sky130_fd_sc_hd__nand2b_1 _80_ (.A_N(net2),
    .B(_09_),
    .Y(_39_));
 sky130_fd_sc_hd__nor2_1 _81_ (.A(net2),
    .B(_09_),
    .Y(_40_));
 sky130_fd_sc_hd__a22oi_1 _82_ (.A1(net2),
    .A2(net10),
    .B1(_40_),
    .B2(net26),
    .Y(_41_));
 sky130_fd_sc_hd__o21ai_0 _83_ (.A1(_38_),
    .A2(_39_),
    .B1(_41_),
    .Y(_07_));
 sky130_fd_sc_hd__clkbuf_1 _84_ (.A(net27),
    .X(net19));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[4]$_DFFE_PN0P_  (.D(_04_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[5]$_DFFE_PN0P_  (.D(_05_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[6]$_DFFE_PN0P_  (.D(_06_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg[7]$_DFFE_PN0P_  (.D(_07_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 hold1 (.A(net28),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_30 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(load_seed),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(seed[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(seed[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(seed[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(seed[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(seed[4]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(seed[5]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(seed[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(seed[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(tap_pattern[0]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(tap_pattern[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(tap_pattern[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(tap_pattern[3]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(tap_pattern[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(tap_pattern[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(tap_pattern[6]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(tap_pattern[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(parallel_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(parallel_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(parallel_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(parallel_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(parallel_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(parallel_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(parallel_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(parallel_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(serial_out));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net28));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_115 ();
endmodule
