module dual_clock_fifo (almost_empty,
    almost_full,
    empty,
    full,
    rd_clk,
    rd_en,
    rd_rst_n,
    wr_clk,
    wr_en,
    wr_rst_n,
    fifo_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 output empty;
 output full;
 input rd_clk;
 input rd_en;
 input rd_rst_n;
 input wr_clk;
 input wr_en;
 input wr_rst_n;
 output [4:0] fifo_count;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_bin_wr_sync[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_wr_sync1[0] ;
 wire \rd_ptr_gray_wr_sync1[1] ;
 wire \rd_ptr_gray_wr_sync1[2] ;
 wire \rd_ptr_gray_wr_sync1[3] ;
 wire \rd_ptr_gray_wr_sync1[4] ;
 wire \rd_ptr_gray_wr_sync2[0] ;
 wire \rd_ptr_gray_wr_sync2[1] ;
 wire \rd_ptr_gray_wr_sync2[2] ;
 wire \rd_ptr_gray_wr_sync2[3] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_bin_rd_sync[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_rd_sync1[0] ;
 wire \wr_ptr_gray_rd_sync1[1] ;
 wire \wr_ptr_gray_rd_sync1[2] ;
 wire \wr_ptr_gray_rd_sync1[3] ;
 wire \wr_ptr_gray_rd_sync1[4] ;
 wire \wr_ptr_gray_rd_sync2[0] ;
 wire \wr_ptr_gray_rd_sync2[1] ;
 wire \wr_ptr_gray_rd_sync2[2] ;
 wire \wr_ptr_gray_rd_sync2[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;

 XOR2_X2 _0654_ (.A(\wr_ptr_gray[1] ),
    .B(\rd_ptr_gray_wr_sync2[1] ),
    .Z(_0160_));
 XOR2_X2 _0655_ (.A(\wr_ptr_gray[2] ),
    .B(\rd_ptr_gray_wr_sync2[2] ),
    .Z(_0161_));
 XOR2_X2 _0656_ (.A(\wr_ptr_gray[3] ),
    .B(\rd_ptr_gray_wr_sync2[3] ),
    .Z(_0162_));
 NOR3_X4 _0657_ (.A1(_0160_),
    .A2(_0161_),
    .A3(_0162_),
    .ZN(_0163_));
 XNOR2_X2 _0658_ (.A(\wr_ptr_bin[4] ),
    .B(\rd_ptr_bin_wr_sync[4] ),
    .ZN(_0164_));
 XOR2_X2 _0659_ (.A(\wr_ptr_gray[0] ),
    .B(\rd_ptr_gray_wr_sync2[0] ),
    .Z(_0165_));
 NOR2_X2 _0660_ (.A1(_0164_),
    .A2(_0165_),
    .ZN(_0166_));
 NAND2_X2 _0661_ (.A1(_0163_),
    .A2(_0166_),
    .ZN(_0167_));
 INV_X4 _0662_ (.A(_0167_),
    .ZN(net15));
 XOR2_X2 _0663_ (.A(\wr_ptr_bin_rd_sync[4] ),
    .B(\rd_ptr_bin[4] ),
    .Z(_0168_));
 XNOR2_X1 _0664_ (.A(\wr_ptr_gray_rd_sync2[3] ),
    .B(\rd_ptr_gray[3] ),
    .ZN(_0169_));
 XNOR2_X2 _0665_ (.A(\wr_ptr_gray_rd_sync2[0] ),
    .B(\rd_ptr_gray[0] ),
    .ZN(_0170_));
 XNOR2_X1 _0666_ (.A(\wr_ptr_gray_rd_sync2[1] ),
    .B(\rd_ptr_gray[1] ),
    .ZN(_0171_));
 XNOR2_X2 _0667_ (.A(\wr_ptr_gray_rd_sync2[2] ),
    .B(\rd_ptr_gray[2] ),
    .ZN(_0172_));
 NAND4_X2 _0668_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0171_),
    .A4(_0172_),
    .ZN(_0173_));
 NOR2_X1 _0669_ (.A1(_0168_),
    .A2(_0173_),
    .ZN(net9));
 XOR2_X2 _0670_ (.A(\wr_ptr_gray_rd_sync2[3] ),
    .B(\wr_ptr_bin_rd_sync[4] ),
    .Z(_0621_));
 XOR2_X2 _0671_ (.A(\wr_ptr_gray_rd_sync2[2] ),
    .B(_0621_),
    .Z(_0625_));
 XNOR2_X2 _0672_ (.A(\wr_ptr_gray_rd_sync2[1] ),
    .B(_0625_),
    .ZN(_0618_));
 INV_X1 _0673_ (.A(_0626_),
    .ZN(_0174_));
 INV_X1 _0674_ (.A(_0617_),
    .ZN(_0175_));
 AOI21_X1 _0675_ (.A(_0630_),
    .B1(_0175_),
    .B2(_0631_),
    .ZN(_0176_));
 INV_X1 _0676_ (.A(_0627_),
    .ZN(_0177_));
 OAI21_X1 _0677_ (.A(_0174_),
    .B1(_0176_),
    .B2(_0177_),
    .ZN(_0178_));
 XOR2_X1 _0678_ (.A(_0623_),
    .B(_0178_),
    .Z(net13));
 INV_X1 _0679_ (.A(_0653_),
    .ZN(net10));
 OAI21_X1 _0680_ (.A(_0174_),
    .B1(_0177_),
    .B2(_0619_),
    .ZN(_0179_));
 AOI21_X1 _0681_ (.A(_0622_),
    .B1(_0179_),
    .B2(_0623_),
    .ZN(_0180_));
 XOR2_X1 _0682_ (.A(_0168_),
    .B(_0180_),
    .Z(net14));
 XNOR2_X2 _0683_ (.A(\rd_ptr_bin_wr_sync[4] ),
    .B(\rd_ptr_gray_wr_sync2[3] ),
    .ZN(_0632_));
 XOR2_X2 _0684_ (.A(\rd_ptr_gray_wr_sync2[2] ),
    .B(_0632_),
    .Z(_0635_));
 XOR2_X2 _0685_ (.A(\rd_ptr_gray_wr_sync2[1] ),
    .B(_0635_),
    .Z(_0614_));
 INV_X1 _0686_ (.A(_0641_),
    .ZN(_0613_));
 INV_X1 _0687_ (.A(_0618_),
    .ZN(_0629_));
 XNOR2_X1 _0688_ (.A(\rd_ptr_gray_wr_sync2[0] ),
    .B(_0614_),
    .ZN(_0640_));
 XOR2_X2 _0689_ (.A(\wr_ptr_gray_rd_sync2[0] ),
    .B(_0618_),
    .Z(_0652_));
 BUF_X1 _0690_ (.A(wr_data[0]),
    .Z(_0181_));
 BUF_X2 _0691_ (.A(_0181_),
    .Z(_0182_));
 BUF_X4 _0692_ (.A(\wr_ptr_bin[3] ),
    .Z(_0183_));
 INV_X1 _0693_ (.A(_0645_),
    .ZN(_0184_));
 INV_X1 _0694_ (.A(\wr_ptr_bin[2] ),
    .ZN(_0185_));
 NAND2_X4 _0695_ (.A1(net5),
    .A2(_0185_),
    .ZN(_0186_));
 NOR4_X4 _0696_ (.A1(_0183_),
    .A2(_0184_),
    .A3(net15),
    .A4(_0186_),
    .ZN(_0187_));
 MUX2_X1 _0697_ (.A(\mem[0][0] ),
    .B(_0182_),
    .S(_0187_),
    .Z(_0006_));
 CLKBUF_X2 _0698_ (.A(wr_data[1]),
    .Z(_0188_));
 BUF_X2 _0699_ (.A(_0188_),
    .Z(_0189_));
 MUX2_X1 _0700_ (.A(\mem[0][1] ),
    .B(_0189_),
    .S(_0187_),
    .Z(_0007_));
 CLKBUF_X2 _0701_ (.A(wr_data[2]),
    .Z(_0190_));
 BUF_X2 _0702_ (.A(_0190_),
    .Z(_0191_));
 MUX2_X1 _0703_ (.A(\mem[0][2] ),
    .B(_0191_),
    .S(_0187_),
    .Z(_0008_));
 BUF_X1 _0704_ (.A(wr_data[3]),
    .Z(_0192_));
 BUF_X2 _0705_ (.A(_0192_),
    .Z(_0193_));
 MUX2_X1 _0706_ (.A(\mem[0][3] ),
    .B(_0193_),
    .S(_0187_),
    .Z(_0009_));
 BUF_X1 _0707_ (.A(wr_data[4]),
    .Z(_0194_));
 BUF_X2 _0708_ (.A(_0194_),
    .Z(_0195_));
 MUX2_X1 _0709_ (.A(\mem[0][4] ),
    .B(_0195_),
    .S(_0187_),
    .Z(_0010_));
 BUF_X1 _0710_ (.A(wr_data[5]),
    .Z(_0196_));
 BUF_X2 _0711_ (.A(_0196_),
    .Z(_0197_));
 MUX2_X1 _0712_ (.A(\mem[0][5] ),
    .B(_0197_),
    .S(_0187_),
    .Z(_0011_));
 BUF_X1 _0713_ (.A(wr_data[6]),
    .Z(_0198_));
 BUF_X2 _0714_ (.A(_0198_),
    .Z(_0199_));
 MUX2_X1 _0715_ (.A(\mem[0][6] ),
    .B(_0199_),
    .S(_0187_),
    .Z(_0012_));
 BUF_X1 _0716_ (.A(wr_data[7]),
    .Z(_0200_));
 BUF_X2 _0717_ (.A(_0200_),
    .Z(_0201_));
 MUX2_X1 _0718_ (.A(\mem[0][7] ),
    .B(_0201_),
    .S(_0187_),
    .Z(_0013_));
 INV_X1 _0719_ (.A(net5),
    .ZN(_0202_));
 NOR2_X1 _0720_ (.A1(_0202_),
    .A2(\wr_ptr_bin[2] ),
    .ZN(_0203_));
 AND4_X1 _0721_ (.A1(_0183_),
    .A2(_0646_),
    .A3(_0167_),
    .A4(_0203_),
    .ZN(_0204_));
 CLKBUF_X3 _0722_ (.A(_0204_),
    .Z(_0205_));
 MUX2_X1 _0723_ (.A(\mem[10][0] ),
    .B(_0182_),
    .S(_0205_),
    .Z(_0014_));
 MUX2_X1 _0724_ (.A(\mem[10][1] ),
    .B(_0189_),
    .S(_0205_),
    .Z(_0015_));
 MUX2_X1 _0725_ (.A(\mem[10][2] ),
    .B(_0191_),
    .S(_0205_),
    .Z(_0016_));
 MUX2_X1 _0726_ (.A(\mem[10][3] ),
    .B(_0193_),
    .S(_0205_),
    .Z(_0017_));
 MUX2_X1 _0727_ (.A(\mem[10][4] ),
    .B(_0195_),
    .S(_0205_),
    .Z(_0018_));
 MUX2_X1 _0728_ (.A(\mem[10][5] ),
    .B(_0197_),
    .S(_0205_),
    .Z(_0019_));
 MUX2_X1 _0729_ (.A(\mem[10][6] ),
    .B(_0199_),
    .S(_0205_),
    .Z(_0020_));
 MUX2_X1 _0730_ (.A(\mem[10][7] ),
    .B(_0201_),
    .S(_0205_),
    .Z(_0021_));
 BUF_X2 _0731_ (.A(_0650_),
    .Z(_0206_));
 AND4_X1 _0732_ (.A1(_0183_),
    .A2(_0206_),
    .A3(_0167_),
    .A4(_0203_),
    .ZN(_0207_));
 CLKBUF_X3 _0733_ (.A(_0207_),
    .Z(_0208_));
 MUX2_X1 _0734_ (.A(\mem[11][0] ),
    .B(_0182_),
    .S(_0208_),
    .Z(_0022_));
 MUX2_X1 _0735_ (.A(\mem[11][1] ),
    .B(_0189_),
    .S(_0208_),
    .Z(_0023_));
 MUX2_X1 _0736_ (.A(\mem[11][2] ),
    .B(_0191_),
    .S(_0208_),
    .Z(_0024_));
 MUX2_X1 _0737_ (.A(\mem[11][3] ),
    .B(_0193_),
    .S(_0208_),
    .Z(_0025_));
 MUX2_X1 _0738_ (.A(\mem[11][4] ),
    .B(_0195_),
    .S(_0208_),
    .Z(_0026_));
 MUX2_X1 _0739_ (.A(\mem[11][5] ),
    .B(_0197_),
    .S(_0208_),
    .Z(_0027_));
 MUX2_X1 _0740_ (.A(\mem[11][6] ),
    .B(_0199_),
    .S(_0208_),
    .Z(_0028_));
 MUX2_X1 _0741_ (.A(\mem[11][7] ),
    .B(_0201_),
    .S(_0208_),
    .Z(_0029_));
 AOI21_X4 _0742_ (.A(_0202_),
    .B1(_0163_),
    .B2(_0166_),
    .ZN(_0209_));
 BUF_X4 _0743_ (.A(_0209_),
    .Z(_0210_));
 AND2_X1 _0744_ (.A1(\wr_ptr_bin[2] ),
    .A2(\wr_ptr_bin[3] ),
    .ZN(_0211_));
 BUF_X4 _0745_ (.A(_0211_),
    .Z(_0212_));
 NAND3_X4 _0746_ (.A1(_0645_),
    .A2(_0210_),
    .A3(_0212_),
    .ZN(_0213_));
 MUX2_X1 _0747_ (.A(_0181_),
    .B(\mem[12][0] ),
    .S(_0213_),
    .Z(_0030_));
 MUX2_X1 _0748_ (.A(_0188_),
    .B(\mem[12][1] ),
    .S(_0213_),
    .Z(_0031_));
 MUX2_X1 _0749_ (.A(_0190_),
    .B(\mem[12][2] ),
    .S(_0213_),
    .Z(_0032_));
 MUX2_X1 _0750_ (.A(_0192_),
    .B(\mem[12][3] ),
    .S(_0213_),
    .Z(_0033_));
 MUX2_X1 _0751_ (.A(_0194_),
    .B(\mem[12][4] ),
    .S(_0213_),
    .Z(_0034_));
 MUX2_X1 _0752_ (.A(_0196_),
    .B(\mem[12][5] ),
    .S(_0213_),
    .Z(_0035_));
 MUX2_X1 _0753_ (.A(_0198_),
    .B(\mem[12][6] ),
    .S(_0213_),
    .Z(_0036_));
 MUX2_X1 _0754_ (.A(_0200_),
    .B(\mem[12][7] ),
    .S(_0213_),
    .Z(_0037_));
 NAND3_X4 _0755_ (.A1(_0648_),
    .A2(_0210_),
    .A3(_0212_),
    .ZN(_0214_));
 MUX2_X1 _0756_ (.A(_0181_),
    .B(\mem[13][0] ),
    .S(_0214_),
    .Z(_0038_));
 MUX2_X1 _0757_ (.A(_0188_),
    .B(\mem[13][1] ),
    .S(_0214_),
    .Z(_0039_));
 MUX2_X1 _0758_ (.A(_0190_),
    .B(\mem[13][2] ),
    .S(_0214_),
    .Z(_0040_));
 MUX2_X1 _0759_ (.A(_0192_),
    .B(\mem[13][3] ),
    .S(_0214_),
    .Z(_0041_));
 MUX2_X1 _0760_ (.A(_0194_),
    .B(\mem[13][4] ),
    .S(_0214_),
    .Z(_0042_));
 MUX2_X1 _0761_ (.A(_0196_),
    .B(\mem[13][5] ),
    .S(_0214_),
    .Z(_0043_));
 MUX2_X1 _0762_ (.A(_0198_),
    .B(\mem[13][6] ),
    .S(_0214_),
    .Z(_0044_));
 MUX2_X1 _0763_ (.A(_0200_),
    .B(\mem[13][7] ),
    .S(_0214_),
    .Z(_0045_));
 NAND3_X4 _0764_ (.A1(_0646_),
    .A2(_0209_),
    .A3(_0212_),
    .ZN(_0215_));
 MUX2_X1 _0765_ (.A(_0181_),
    .B(\mem[14][0] ),
    .S(_0215_),
    .Z(_0046_));
 MUX2_X1 _0766_ (.A(_0188_),
    .B(\mem[14][1] ),
    .S(_0215_),
    .Z(_0047_));
 MUX2_X1 _0767_ (.A(_0190_),
    .B(\mem[14][2] ),
    .S(_0215_),
    .Z(_0048_));
 MUX2_X1 _0768_ (.A(_0192_),
    .B(\mem[14][3] ),
    .S(_0215_),
    .Z(_0049_));
 MUX2_X1 _0769_ (.A(_0194_),
    .B(\mem[14][4] ),
    .S(_0215_),
    .Z(_0050_));
 MUX2_X1 _0770_ (.A(_0196_),
    .B(\mem[14][5] ),
    .S(_0215_),
    .Z(_0051_));
 MUX2_X1 _0771_ (.A(_0198_),
    .B(\mem[14][6] ),
    .S(_0215_),
    .Z(_0052_));
 MUX2_X1 _0772_ (.A(_0200_),
    .B(\mem[14][7] ),
    .S(_0215_),
    .Z(_0053_));
 NAND3_X4 _0773_ (.A1(_0206_),
    .A2(_0209_),
    .A3(_0212_),
    .ZN(_0216_));
 MUX2_X1 _0774_ (.A(_0181_),
    .B(\mem[15][0] ),
    .S(_0216_),
    .Z(_0054_));
 MUX2_X1 _0775_ (.A(_0188_),
    .B(\mem[15][1] ),
    .S(_0216_),
    .Z(_0055_));
 MUX2_X1 _0776_ (.A(_0190_),
    .B(\mem[15][2] ),
    .S(_0216_),
    .Z(_0056_));
 MUX2_X1 _0777_ (.A(_0192_),
    .B(\mem[15][3] ),
    .S(_0216_),
    .Z(_0057_));
 MUX2_X1 _0778_ (.A(_0194_),
    .B(\mem[15][4] ),
    .S(_0216_),
    .Z(_0058_));
 MUX2_X1 _0779_ (.A(_0196_),
    .B(\mem[15][5] ),
    .S(_0216_),
    .Z(_0059_));
 MUX2_X1 _0780_ (.A(_0198_),
    .B(\mem[15][6] ),
    .S(_0216_),
    .Z(_0060_));
 MUX2_X1 _0781_ (.A(_0200_),
    .B(\mem[15][7] ),
    .S(_0216_),
    .Z(_0061_));
 INV_X1 _0782_ (.A(_0648_),
    .ZN(_0217_));
 NOR4_X4 _0783_ (.A1(_0183_),
    .A2(_0217_),
    .A3(net15),
    .A4(_0186_),
    .ZN(_0218_));
 MUX2_X1 _0784_ (.A(\mem[1][0] ),
    .B(_0182_),
    .S(_0218_),
    .Z(_0062_));
 MUX2_X1 _0785_ (.A(\mem[1][1] ),
    .B(_0189_),
    .S(_0218_),
    .Z(_0063_));
 MUX2_X1 _0786_ (.A(\mem[1][2] ),
    .B(_0191_),
    .S(_0218_),
    .Z(_0064_));
 MUX2_X1 _0787_ (.A(\mem[1][3] ),
    .B(_0193_),
    .S(_0218_),
    .Z(_0065_));
 MUX2_X1 _0788_ (.A(\mem[1][4] ),
    .B(_0195_),
    .S(_0218_),
    .Z(_0066_));
 MUX2_X1 _0789_ (.A(\mem[1][5] ),
    .B(_0197_),
    .S(_0218_),
    .Z(_0067_));
 MUX2_X1 _0790_ (.A(\mem[1][6] ),
    .B(_0199_),
    .S(_0218_),
    .Z(_0068_));
 MUX2_X1 _0791_ (.A(\mem[1][7] ),
    .B(_0201_),
    .S(_0218_),
    .Z(_0069_));
 INV_X1 _0792_ (.A(_0646_),
    .ZN(_0219_));
 NOR4_X4 _0793_ (.A1(_0183_),
    .A2(_0219_),
    .A3(net15),
    .A4(_0186_),
    .ZN(_0220_));
 MUX2_X1 _0794_ (.A(\mem[2][0] ),
    .B(_0182_),
    .S(_0220_),
    .Z(_0070_));
 MUX2_X1 _0795_ (.A(\mem[2][1] ),
    .B(_0189_),
    .S(_0220_),
    .Z(_0071_));
 MUX2_X1 _0796_ (.A(\mem[2][2] ),
    .B(_0191_),
    .S(_0220_),
    .Z(_0072_));
 MUX2_X1 _0797_ (.A(\mem[2][3] ),
    .B(_0193_),
    .S(_0220_),
    .Z(_0073_));
 MUX2_X1 _0798_ (.A(\mem[2][4] ),
    .B(_0195_),
    .S(_0220_),
    .Z(_0074_));
 MUX2_X1 _0799_ (.A(\mem[2][5] ),
    .B(_0197_),
    .S(_0220_),
    .Z(_0075_));
 MUX2_X1 _0800_ (.A(\mem[2][6] ),
    .B(_0199_),
    .S(_0220_),
    .Z(_0076_));
 MUX2_X1 _0801_ (.A(\mem[2][7] ),
    .B(_0201_),
    .S(_0220_),
    .Z(_0077_));
 INV_X1 _0802_ (.A(_0206_),
    .ZN(_0221_));
 NOR4_X4 _0803_ (.A1(_0183_),
    .A2(_0221_),
    .A3(net15),
    .A4(_0186_),
    .ZN(_0222_));
 MUX2_X1 _0804_ (.A(\mem[3][0] ),
    .B(_0182_),
    .S(_0222_),
    .Z(_0078_));
 MUX2_X1 _0805_ (.A(\mem[3][1] ),
    .B(_0189_),
    .S(_0222_),
    .Z(_0079_));
 MUX2_X1 _0806_ (.A(\mem[3][2] ),
    .B(_0191_),
    .S(_0222_),
    .Z(_0080_));
 MUX2_X1 _0807_ (.A(\mem[3][3] ),
    .B(_0193_),
    .S(_0222_),
    .Z(_0081_));
 MUX2_X1 _0808_ (.A(\mem[3][4] ),
    .B(_0195_),
    .S(_0222_),
    .Z(_0082_));
 MUX2_X1 _0809_ (.A(\mem[3][5] ),
    .B(_0197_),
    .S(_0222_),
    .Z(_0083_));
 MUX2_X1 _0810_ (.A(\mem[3][6] ),
    .B(_0199_),
    .S(_0222_),
    .Z(_0084_));
 MUX2_X1 _0811_ (.A(\mem[3][7] ),
    .B(_0201_),
    .S(_0222_),
    .Z(_0085_));
 NOR2_X1 _0812_ (.A1(_0185_),
    .A2(_0183_),
    .ZN(_0223_));
 AND3_X1 _0813_ (.A1(_0645_),
    .A2(_0209_),
    .A3(_0223_),
    .ZN(_0224_));
 BUF_X4 _0814_ (.A(_0224_),
    .Z(_0225_));
 MUX2_X1 _0815_ (.A(\mem[4][0] ),
    .B(_0182_),
    .S(_0225_),
    .Z(_0086_));
 MUX2_X1 _0816_ (.A(\mem[4][1] ),
    .B(_0189_),
    .S(_0225_),
    .Z(_0087_));
 MUX2_X1 _0817_ (.A(\mem[4][2] ),
    .B(_0191_),
    .S(_0225_),
    .Z(_0088_));
 MUX2_X1 _0818_ (.A(\mem[4][3] ),
    .B(_0193_),
    .S(_0225_),
    .Z(_0089_));
 MUX2_X1 _0819_ (.A(\mem[4][4] ),
    .B(_0195_),
    .S(_0225_),
    .Z(_0090_));
 MUX2_X1 _0820_ (.A(\mem[4][5] ),
    .B(_0197_),
    .S(_0225_),
    .Z(_0091_));
 MUX2_X1 _0821_ (.A(\mem[4][6] ),
    .B(_0199_),
    .S(_0225_),
    .Z(_0092_));
 MUX2_X1 _0822_ (.A(\mem[4][7] ),
    .B(_0201_),
    .S(_0225_),
    .Z(_0093_));
 AND3_X1 _0823_ (.A1(_0648_),
    .A2(_0209_),
    .A3(_0223_),
    .ZN(_0226_));
 BUF_X4 _0824_ (.A(_0226_),
    .Z(_0227_));
 MUX2_X1 _0825_ (.A(\mem[5][0] ),
    .B(_0182_),
    .S(_0227_),
    .Z(_0094_));
 MUX2_X1 _0826_ (.A(\mem[5][1] ),
    .B(_0189_),
    .S(_0227_),
    .Z(_0095_));
 MUX2_X1 _0827_ (.A(\mem[5][2] ),
    .B(_0191_),
    .S(_0227_),
    .Z(_0096_));
 MUX2_X1 _0828_ (.A(\mem[5][3] ),
    .B(_0193_),
    .S(_0227_),
    .Z(_0097_));
 MUX2_X1 _0829_ (.A(\mem[5][4] ),
    .B(_0195_),
    .S(_0227_),
    .Z(_0098_));
 MUX2_X1 _0830_ (.A(\mem[5][5] ),
    .B(_0197_),
    .S(_0227_),
    .Z(_0099_));
 MUX2_X1 _0831_ (.A(\mem[5][6] ),
    .B(_0199_),
    .S(_0227_),
    .Z(_0100_));
 MUX2_X1 _0832_ (.A(\mem[5][7] ),
    .B(_0201_),
    .S(_0227_),
    .Z(_0101_));
 AND3_X1 _0833_ (.A1(_0646_),
    .A2(_0209_),
    .A3(_0223_),
    .ZN(_0228_));
 BUF_X4 _0834_ (.A(_0228_),
    .Z(_0229_));
 MUX2_X1 _0835_ (.A(\mem[6][0] ),
    .B(_0182_),
    .S(_0229_),
    .Z(_0102_));
 MUX2_X1 _0836_ (.A(\mem[6][1] ),
    .B(_0189_),
    .S(_0229_),
    .Z(_0103_));
 MUX2_X1 _0837_ (.A(\mem[6][2] ),
    .B(_0191_),
    .S(_0229_),
    .Z(_0104_));
 MUX2_X1 _0838_ (.A(\mem[6][3] ),
    .B(_0193_),
    .S(_0229_),
    .Z(_0105_));
 MUX2_X1 _0839_ (.A(\mem[6][4] ),
    .B(_0195_),
    .S(_0229_),
    .Z(_0106_));
 MUX2_X1 _0840_ (.A(\mem[6][5] ),
    .B(_0197_),
    .S(_0229_),
    .Z(_0107_));
 MUX2_X1 _0841_ (.A(\mem[6][6] ),
    .B(_0199_),
    .S(_0229_),
    .Z(_0108_));
 MUX2_X1 _0842_ (.A(\mem[6][7] ),
    .B(_0201_),
    .S(_0229_),
    .Z(_0109_));
 AND3_X1 _0843_ (.A1(_0206_),
    .A2(_0209_),
    .A3(_0223_),
    .ZN(_0230_));
 BUF_X4 _0844_ (.A(_0230_),
    .Z(_0231_));
 MUX2_X1 _0845_ (.A(\mem[7][0] ),
    .B(_0182_),
    .S(_0231_),
    .Z(_0110_));
 MUX2_X1 _0846_ (.A(\mem[7][1] ),
    .B(_0189_),
    .S(_0231_),
    .Z(_0111_));
 MUX2_X1 _0847_ (.A(\mem[7][2] ),
    .B(_0191_),
    .S(_0231_),
    .Z(_0112_));
 MUX2_X1 _0848_ (.A(\mem[7][3] ),
    .B(_0193_),
    .S(_0231_),
    .Z(_0113_));
 MUX2_X1 _0849_ (.A(\mem[7][4] ),
    .B(_0195_),
    .S(_0231_),
    .Z(_0114_));
 MUX2_X1 _0850_ (.A(\mem[7][5] ),
    .B(_0197_),
    .S(_0231_),
    .Z(_0115_));
 MUX2_X1 _0851_ (.A(\mem[7][6] ),
    .B(_0199_),
    .S(_0231_),
    .Z(_0116_));
 MUX2_X1 _0852_ (.A(\mem[7][7] ),
    .B(_0201_),
    .S(_0231_),
    .Z(_0117_));
 AND4_X1 _0853_ (.A1(_0183_),
    .A2(_0645_),
    .A3(_0167_),
    .A4(_0203_),
    .ZN(_0232_));
 CLKBUF_X3 _0854_ (.A(_0232_),
    .Z(_0233_));
 MUX2_X1 _0855_ (.A(\mem[8][0] ),
    .B(_0181_),
    .S(_0233_),
    .Z(_0118_));
 MUX2_X1 _0856_ (.A(\mem[8][1] ),
    .B(_0188_),
    .S(_0233_),
    .Z(_0119_));
 MUX2_X1 _0857_ (.A(\mem[8][2] ),
    .B(_0190_),
    .S(_0233_),
    .Z(_0120_));
 MUX2_X1 _0858_ (.A(\mem[8][3] ),
    .B(_0192_),
    .S(_0233_),
    .Z(_0121_));
 MUX2_X1 _0859_ (.A(\mem[8][4] ),
    .B(_0194_),
    .S(_0233_),
    .Z(_0122_));
 MUX2_X1 _0860_ (.A(\mem[8][5] ),
    .B(_0196_),
    .S(_0233_),
    .Z(_0123_));
 MUX2_X1 _0861_ (.A(\mem[8][6] ),
    .B(_0198_),
    .S(_0233_),
    .Z(_0124_));
 MUX2_X1 _0862_ (.A(\mem[8][7] ),
    .B(_0200_),
    .S(_0233_),
    .Z(_0125_));
 AND4_X1 _0863_ (.A1(_0183_),
    .A2(_0648_),
    .A3(_0167_),
    .A4(_0203_),
    .ZN(_0234_));
 CLKBUF_X3 _0864_ (.A(_0234_),
    .Z(_0235_));
 MUX2_X1 _0865_ (.A(\mem[9][0] ),
    .B(_0181_),
    .S(_0235_),
    .Z(_0126_));
 MUX2_X1 _0866_ (.A(\mem[9][1] ),
    .B(_0188_),
    .S(_0235_),
    .Z(_0127_));
 MUX2_X1 _0867_ (.A(\mem[9][2] ),
    .B(_0190_),
    .S(_0235_),
    .Z(_0128_));
 MUX2_X1 _0868_ (.A(\mem[9][3] ),
    .B(_0192_),
    .S(_0235_),
    .Z(_0129_));
 MUX2_X1 _0869_ (.A(\mem[9][4] ),
    .B(_0194_),
    .S(_0235_),
    .Z(_0130_));
 MUX2_X1 _0870_ (.A(\mem[9][5] ),
    .B(_0196_),
    .S(_0235_),
    .Z(_0131_));
 MUX2_X1 _0871_ (.A(\mem[9][6] ),
    .B(_0198_),
    .S(_0235_),
    .Z(_0132_));
 MUX2_X1 _0872_ (.A(\mem[9][7] ),
    .B(_0200_),
    .S(_0235_),
    .Z(_0133_));
 OAI21_X4 _0873_ (.A(net2),
    .B1(_0168_),
    .B2(_0173_),
    .ZN(_0236_));
 BUF_X4 _0874_ (.A(_0236_),
    .Z(_0237_));
 BUF_X4 _0875_ (.A(\rd_ptr_bin[2] ),
    .Z(_0238_));
 BUF_X8 _0876_ (.A(_0238_),
    .Z(_0239_));
 BUF_X4 _0877_ (.A(_0239_),
    .Z(_0240_));
 MUX2_X1 _0878_ (.A(\mem[3][0] ),
    .B(\mem[7][0] ),
    .S(_0240_),
    .Z(_0241_));
 BUF_X2 _0879_ (.A(\rd_ptr_bin[0] ),
    .Z(_0242_));
 BUF_X2 _0880_ (.A(\rd_ptr_bin[1] ),
    .Z(_0243_));
 BUF_X4 _0881_ (.A(_0243_),
    .Z(_0244_));
 NAND2_X4 _0882_ (.A1(_0242_),
    .A2(_0244_),
    .ZN(_0245_));
 NOR2_X1 _0883_ (.A1(_0241_),
    .A2(_0245_),
    .ZN(_0246_));
 INV_X4 _0884_ (.A(_0242_),
    .ZN(_0247_));
 NOR2_X4 _0885_ (.A1(_0247_),
    .A2(_0244_),
    .ZN(_0248_));
 MUX2_X1 _0886_ (.A(\mem[1][0] ),
    .B(\mem[5][0] ),
    .S(_0240_),
    .Z(_0249_));
 INV_X1 _0887_ (.A(_0249_),
    .ZN(_0250_));
 AOI21_X1 _0888_ (.A(_0246_),
    .B1(_0248_),
    .B2(_0250_),
    .ZN(_0251_));
 CLKBUF_X3 _0889_ (.A(\rd_ptr_bin[3] ),
    .Z(_0252_));
 BUF_X4 _0890_ (.A(_0252_),
    .Z(_0253_));
 MUX2_X1 _0891_ (.A(\mem[0][0] ),
    .B(\mem[4][0] ),
    .S(_0240_),
    .Z(_0254_));
 OR2_X1 _0892_ (.A1(_0242_),
    .A2(_0243_),
    .ZN(_0255_));
 BUF_X2 _0893_ (.A(_0255_),
    .Z(_0256_));
 NOR2_X1 _0894_ (.A1(_0254_),
    .A2(_0256_),
    .ZN(_0257_));
 CLKBUF_X3 _0895_ (.A(_0242_),
    .Z(_0258_));
 INV_X2 _0896_ (.A(_0243_),
    .ZN(_0259_));
 BUF_X8 _0897_ (.A(_0239_),
    .Z(_0260_));
 MUX2_X1 _0898_ (.A(\mem[2][0] ),
    .B(\mem[6][0] ),
    .S(_0260_),
    .Z(_0261_));
 NOR3_X1 _0899_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0261_),
    .ZN(_0262_));
 NOR3_X1 _0900_ (.A1(_0253_),
    .A2(_0257_),
    .A3(_0262_),
    .ZN(_0263_));
 MUX2_X1 _0901_ (.A(\mem[9][0] ),
    .B(\mem[13][0] ),
    .S(_0239_),
    .Z(_0264_));
 BUF_X4 _0902_ (.A(_0238_),
    .Z(_0265_));
 MUX2_X1 _0903_ (.A(\mem[11][0] ),
    .B(\mem[15][0] ),
    .S(_0265_),
    .Z(_0266_));
 BUF_X4 _0904_ (.A(_0243_),
    .Z(_0267_));
 MUX2_X1 _0905_ (.A(_0264_),
    .B(_0266_),
    .S(_0267_),
    .Z(_0268_));
 BUF_X4 _0906_ (.A(_0238_),
    .Z(_0269_));
 MUX2_X1 _0907_ (.A(\mem[8][0] ),
    .B(\mem[12][0] ),
    .S(_0269_),
    .Z(_0270_));
 BUF_X4 _0908_ (.A(_0238_),
    .Z(_0271_));
 MUX2_X1 _0909_ (.A(\mem[10][0] ),
    .B(\mem[14][0] ),
    .S(_0271_),
    .Z(_0272_));
 MUX2_X1 _0910_ (.A(_0270_),
    .B(_0272_),
    .S(_0244_),
    .Z(_0273_));
 MUX2_X1 _0911_ (.A(_0268_),
    .B(_0273_),
    .S(_0247_),
    .Z(_0274_));
 AOI221_X2 _0912_ (.A(_0237_),
    .B1(_0251_),
    .B2(_0263_),
    .C1(_0274_),
    .C2(_0253_),
    .ZN(_0275_));
 BUF_X4 _0913_ (.A(_0237_),
    .Z(_0276_));
 INV_X1 _0914_ (.A(net16),
    .ZN(_0277_));
 AOI21_X1 _0915_ (.A(_0275_),
    .B1(_0276_),
    .B2(_0277_),
    .ZN(_0134_));
 MUX2_X1 _0916_ (.A(\mem[3][1] ),
    .B(\mem[7][1] ),
    .S(_0240_),
    .Z(_0278_));
 NOR2_X1 _0917_ (.A1(_0245_),
    .A2(_0278_),
    .ZN(_0279_));
 BUF_X8 _0918_ (.A(_0260_),
    .Z(_0280_));
 MUX2_X1 _0919_ (.A(\mem[1][1] ),
    .B(\mem[5][1] ),
    .S(_0280_),
    .Z(_0281_));
 INV_X1 _0920_ (.A(_0281_),
    .ZN(_0282_));
 AOI21_X1 _0921_ (.A(_0279_),
    .B1(_0282_),
    .B2(_0248_),
    .ZN(_0283_));
 MUX2_X1 _0922_ (.A(\mem[0][1] ),
    .B(\mem[4][1] ),
    .S(_0260_),
    .Z(_0284_));
 NOR2_X1 _0923_ (.A1(_0256_),
    .A2(_0284_),
    .ZN(_0285_));
 MUX2_X1 _0924_ (.A(\mem[2][1] ),
    .B(\mem[6][1] ),
    .S(_0260_),
    .Z(_0286_));
 NOR3_X1 _0925_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0286_),
    .ZN(_0287_));
 NOR3_X1 _0926_ (.A1(_0252_),
    .A2(_0285_),
    .A3(_0287_),
    .ZN(_0288_));
 MUX2_X1 _0927_ (.A(\mem[9][1] ),
    .B(\mem[13][1] ),
    .S(_0239_),
    .Z(_0289_));
 MUX2_X1 _0928_ (.A(\mem[11][1] ),
    .B(\mem[15][1] ),
    .S(_0265_),
    .Z(_0290_));
 MUX2_X1 _0929_ (.A(_0289_),
    .B(_0290_),
    .S(_0267_),
    .Z(_0291_));
 MUX2_X1 _0930_ (.A(\mem[8][1] ),
    .B(\mem[12][1] ),
    .S(_0269_),
    .Z(_0292_));
 MUX2_X1 _0931_ (.A(\mem[10][1] ),
    .B(\mem[14][1] ),
    .S(_0271_),
    .Z(_0293_));
 MUX2_X1 _0932_ (.A(_0292_),
    .B(_0293_),
    .S(_0244_),
    .Z(_0294_));
 MUX2_X1 _0933_ (.A(_0291_),
    .B(_0294_),
    .S(_0247_),
    .Z(_0295_));
 AOI221_X2 _0934_ (.A(_0237_),
    .B1(_0283_),
    .B2(_0288_),
    .C1(_0295_),
    .C2(_0253_),
    .ZN(_0296_));
 INV_X1 _0935_ (.A(net17),
    .ZN(_0297_));
 AOI21_X1 _0936_ (.A(_0296_),
    .B1(_0276_),
    .B2(_0297_),
    .ZN(_0135_));
 MUX2_X1 _0937_ (.A(\mem[3][2] ),
    .B(\mem[7][2] ),
    .S(_0240_),
    .Z(_0298_));
 NOR2_X1 _0938_ (.A1(_0245_),
    .A2(_0298_),
    .ZN(_0299_));
 MUX2_X1 _0939_ (.A(\mem[1][2] ),
    .B(\mem[5][2] ),
    .S(_0280_),
    .Z(_0300_));
 INV_X1 _0940_ (.A(_0300_),
    .ZN(_0301_));
 AOI21_X1 _0941_ (.A(_0299_),
    .B1(_0301_),
    .B2(_0248_),
    .ZN(_0302_));
 MUX2_X1 _0942_ (.A(\mem[0][2] ),
    .B(\mem[4][2] ),
    .S(_0260_),
    .Z(_0303_));
 NOR2_X1 _0943_ (.A1(_0256_),
    .A2(_0303_),
    .ZN(_0304_));
 MUX2_X1 _0944_ (.A(\mem[2][2] ),
    .B(\mem[6][2] ),
    .S(_0271_),
    .Z(_0305_));
 NOR3_X1 _0945_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0305_),
    .ZN(_0306_));
 NOR3_X1 _0946_ (.A1(_0252_),
    .A2(_0304_),
    .A3(_0306_),
    .ZN(_0307_));
 MUX2_X1 _0947_ (.A(\mem[9][2] ),
    .B(\mem[13][2] ),
    .S(_0239_),
    .Z(_0308_));
 MUX2_X1 _0948_ (.A(\mem[11][2] ),
    .B(\mem[15][2] ),
    .S(_0265_),
    .Z(_0309_));
 MUX2_X1 _0949_ (.A(_0308_),
    .B(_0309_),
    .S(_0267_),
    .Z(_0310_));
 MUX2_X1 _0950_ (.A(\mem[8][2] ),
    .B(\mem[12][2] ),
    .S(_0269_),
    .Z(_0311_));
 MUX2_X1 _0951_ (.A(\mem[10][2] ),
    .B(\mem[14][2] ),
    .S(_0271_),
    .Z(_0312_));
 MUX2_X1 _0952_ (.A(_0311_),
    .B(_0312_),
    .S(_0244_),
    .Z(_0313_));
 MUX2_X1 _0953_ (.A(_0310_),
    .B(_0313_),
    .S(_0247_),
    .Z(_0314_));
 AOI221_X2 _0954_ (.A(_0236_),
    .B1(_0302_),
    .B2(_0307_),
    .C1(_0314_),
    .C2(_0253_),
    .ZN(_0315_));
 INV_X1 _0955_ (.A(net18),
    .ZN(_0316_));
 AOI21_X1 _0956_ (.A(_0315_),
    .B1(_0276_),
    .B2(_0316_),
    .ZN(_0136_));
 MUX2_X1 _0957_ (.A(\mem[3][3] ),
    .B(\mem[7][3] ),
    .S(_0240_),
    .Z(_0317_));
 NOR2_X1 _0958_ (.A1(_0245_),
    .A2(_0317_),
    .ZN(_0318_));
 MUX2_X1 _0959_ (.A(\mem[1][3] ),
    .B(\mem[5][3] ),
    .S(_0280_),
    .Z(_0319_));
 INV_X1 _0960_ (.A(_0319_),
    .ZN(_0320_));
 AOI21_X1 _0961_ (.A(_0318_),
    .B1(_0320_),
    .B2(_0248_),
    .ZN(_0321_));
 MUX2_X1 _0962_ (.A(\mem[0][3] ),
    .B(\mem[4][3] ),
    .S(_0260_),
    .Z(_0322_));
 NOR2_X1 _0963_ (.A1(_0256_),
    .A2(_0322_),
    .ZN(_0323_));
 MUX2_X1 _0964_ (.A(\mem[2][3] ),
    .B(\mem[6][3] ),
    .S(_0271_),
    .Z(_0324_));
 NOR3_X1 _0965_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0324_),
    .ZN(_0325_));
 NOR3_X1 _0966_ (.A1(_0252_),
    .A2(_0323_),
    .A3(_0325_),
    .ZN(_0326_));
 MUX2_X1 _0967_ (.A(\mem[9][3] ),
    .B(\mem[13][3] ),
    .S(_0239_),
    .Z(_0327_));
 MUX2_X1 _0968_ (.A(\mem[11][3] ),
    .B(\mem[15][3] ),
    .S(_0265_),
    .Z(_0328_));
 MUX2_X1 _0969_ (.A(_0327_),
    .B(_0328_),
    .S(_0267_),
    .Z(_0329_));
 MUX2_X1 _0970_ (.A(\mem[8][3] ),
    .B(\mem[12][3] ),
    .S(_0269_),
    .Z(_0330_));
 MUX2_X1 _0971_ (.A(\mem[10][3] ),
    .B(\mem[14][3] ),
    .S(_0271_),
    .Z(_0331_));
 MUX2_X1 _0972_ (.A(_0330_),
    .B(_0331_),
    .S(_0244_),
    .Z(_0332_));
 MUX2_X1 _0973_ (.A(_0329_),
    .B(_0332_),
    .S(_0247_),
    .Z(_0333_));
 AOI221_X2 _0974_ (.A(_0236_),
    .B1(_0321_),
    .B2(_0326_),
    .C1(_0333_),
    .C2(_0253_),
    .ZN(_0334_));
 INV_X1 _0975_ (.A(net19),
    .ZN(_0335_));
 AOI21_X1 _0976_ (.A(_0334_),
    .B1(_0276_),
    .B2(_0335_),
    .ZN(_0137_));
 MUX2_X1 _0977_ (.A(\mem[3][4] ),
    .B(\mem[7][4] ),
    .S(_0240_),
    .Z(_0336_));
 NOR2_X1 _0978_ (.A1(_0245_),
    .A2(_0336_),
    .ZN(_0337_));
 MUX2_X1 _0979_ (.A(\mem[1][4] ),
    .B(\mem[5][4] ),
    .S(_0280_),
    .Z(_0338_));
 INV_X1 _0980_ (.A(_0338_),
    .ZN(_0339_));
 AOI21_X1 _0981_ (.A(_0337_),
    .B1(_0339_),
    .B2(_0248_),
    .ZN(_0340_));
 MUX2_X1 _0982_ (.A(\mem[0][4] ),
    .B(\mem[4][4] ),
    .S(_0260_),
    .Z(_0341_));
 NOR2_X1 _0983_ (.A1(_0256_),
    .A2(_0341_),
    .ZN(_0342_));
 MUX2_X1 _0984_ (.A(\mem[2][4] ),
    .B(\mem[6][4] ),
    .S(_0271_),
    .Z(_0343_));
 NOR3_X1 _0985_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0343_),
    .ZN(_0344_));
 NOR3_X1 _0986_ (.A1(_0252_),
    .A2(_0342_),
    .A3(_0344_),
    .ZN(_0345_));
 MUX2_X1 _0987_ (.A(\mem[9][4] ),
    .B(\mem[13][4] ),
    .S(_0239_),
    .Z(_0346_));
 MUX2_X1 _0988_ (.A(\mem[11][4] ),
    .B(\mem[15][4] ),
    .S(_0265_),
    .Z(_0347_));
 MUX2_X1 _0989_ (.A(_0346_),
    .B(_0347_),
    .S(_0267_),
    .Z(_0348_));
 MUX2_X1 _0990_ (.A(\mem[8][4] ),
    .B(\mem[12][4] ),
    .S(_0269_),
    .Z(_0349_));
 MUX2_X1 _0991_ (.A(\mem[10][4] ),
    .B(\mem[14][4] ),
    .S(_0269_),
    .Z(_0350_));
 MUX2_X1 _0992_ (.A(_0349_),
    .B(_0350_),
    .S(_0244_),
    .Z(_0351_));
 MUX2_X1 _0993_ (.A(_0348_),
    .B(_0351_),
    .S(_0247_),
    .Z(_0352_));
 AOI221_X2 _0994_ (.A(_0236_),
    .B1(_0340_),
    .B2(_0345_),
    .C1(_0352_),
    .C2(_0253_),
    .ZN(_0353_));
 INV_X1 _0995_ (.A(net20),
    .ZN(_0354_));
 AOI21_X1 _0996_ (.A(_0353_),
    .B1(_0276_),
    .B2(_0354_),
    .ZN(_0138_));
 MUX2_X1 _0997_ (.A(\mem[3][5] ),
    .B(\mem[7][5] ),
    .S(_0240_),
    .Z(_0355_));
 NOR2_X1 _0998_ (.A1(_0245_),
    .A2(_0355_),
    .ZN(_0356_));
 MUX2_X1 _0999_ (.A(\mem[1][5] ),
    .B(\mem[5][5] ),
    .S(_0280_),
    .Z(_0357_));
 INV_X1 _1000_ (.A(_0357_),
    .ZN(_0358_));
 AOI21_X1 _1001_ (.A(_0356_),
    .B1(_0358_),
    .B2(_0248_),
    .ZN(_0359_));
 MUX2_X1 _1002_ (.A(\mem[0][5] ),
    .B(\mem[4][5] ),
    .S(_0260_),
    .Z(_0360_));
 NOR2_X1 _1003_ (.A1(_0256_),
    .A2(_0360_),
    .ZN(_0361_));
 MUX2_X1 _1004_ (.A(\mem[2][5] ),
    .B(\mem[6][5] ),
    .S(_0271_),
    .Z(_0362_));
 NOR3_X1 _1005_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0362_),
    .ZN(_0363_));
 NOR3_X1 _1006_ (.A1(_0252_),
    .A2(_0361_),
    .A3(_0363_),
    .ZN(_0364_));
 MUX2_X1 _1007_ (.A(\mem[9][5] ),
    .B(\mem[13][5] ),
    .S(_0239_),
    .Z(_0365_));
 MUX2_X1 _1008_ (.A(\mem[11][5] ),
    .B(\mem[15][5] ),
    .S(_0265_),
    .Z(_0366_));
 MUX2_X1 _1009_ (.A(_0365_),
    .B(_0366_),
    .S(_0267_),
    .Z(_0367_));
 MUX2_X1 _1010_ (.A(\mem[8][5] ),
    .B(\mem[12][5] ),
    .S(_0269_),
    .Z(_0368_));
 MUX2_X1 _1011_ (.A(\mem[10][5] ),
    .B(\mem[14][5] ),
    .S(_0269_),
    .Z(_0369_));
 MUX2_X1 _1012_ (.A(_0368_),
    .B(_0369_),
    .S(_0244_),
    .Z(_0370_));
 MUX2_X1 _1013_ (.A(_0367_),
    .B(_0370_),
    .S(_0247_),
    .Z(_0371_));
 AOI221_X2 _1014_ (.A(_0236_),
    .B1(_0359_),
    .B2(_0364_),
    .C1(_0371_),
    .C2(_0253_),
    .ZN(_0372_));
 INV_X1 _1015_ (.A(net21),
    .ZN(_0373_));
 AOI21_X1 _1016_ (.A(_0372_),
    .B1(_0276_),
    .B2(_0373_),
    .ZN(_0139_));
 MUX2_X1 _1017_ (.A(\mem[3][6] ),
    .B(\mem[7][6] ),
    .S(_0240_),
    .Z(_0374_));
 NOR2_X1 _1018_ (.A1(_0245_),
    .A2(_0374_),
    .ZN(_0375_));
 MUX2_X1 _1019_ (.A(\mem[1][6] ),
    .B(\mem[5][6] ),
    .S(_0280_),
    .Z(_0376_));
 INV_X1 _1020_ (.A(_0376_),
    .ZN(_0377_));
 AOI21_X1 _1021_ (.A(_0375_),
    .B1(_0377_),
    .B2(_0248_),
    .ZN(_0378_));
 MUX2_X1 _1022_ (.A(\mem[0][6] ),
    .B(\mem[4][6] ),
    .S(_0260_),
    .Z(_0379_));
 NOR2_X1 _1023_ (.A1(_0256_),
    .A2(_0379_),
    .ZN(_0380_));
 MUX2_X1 _1024_ (.A(\mem[2][6] ),
    .B(\mem[6][6] ),
    .S(_0271_),
    .Z(_0381_));
 NOR3_X1 _1025_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0381_),
    .ZN(_0382_));
 NOR3_X1 _1026_ (.A1(_0252_),
    .A2(_0380_),
    .A3(_0382_),
    .ZN(_0383_));
 MUX2_X1 _1027_ (.A(\mem[9][6] ),
    .B(\mem[13][6] ),
    .S(_0239_),
    .Z(_0384_));
 MUX2_X1 _1028_ (.A(\mem[11][6] ),
    .B(\mem[15][6] ),
    .S(_0265_),
    .Z(_0385_));
 MUX2_X1 _1029_ (.A(_0384_),
    .B(_0385_),
    .S(_0267_),
    .Z(_0386_));
 MUX2_X1 _1030_ (.A(\mem[8][6] ),
    .B(\mem[12][6] ),
    .S(_0265_),
    .Z(_0387_));
 MUX2_X1 _1031_ (.A(\mem[10][6] ),
    .B(\mem[14][6] ),
    .S(_0269_),
    .Z(_0388_));
 MUX2_X1 _1032_ (.A(_0387_),
    .B(_0388_),
    .S(_0267_),
    .Z(_0389_));
 MUX2_X1 _1033_ (.A(_0386_),
    .B(_0389_),
    .S(_0247_),
    .Z(_0390_));
 AOI221_X2 _1034_ (.A(_0236_),
    .B1(_0378_),
    .B2(_0383_),
    .C1(_0390_),
    .C2(_0253_),
    .ZN(_0391_));
 INV_X1 _1035_ (.A(net22),
    .ZN(_0392_));
 AOI21_X1 _1036_ (.A(_0391_),
    .B1(_0276_),
    .B2(_0392_),
    .ZN(_0140_));
 MUX2_X1 _1037_ (.A(\mem[3][7] ),
    .B(\mem[7][7] ),
    .S(_0240_),
    .Z(_0393_));
 NOR2_X1 _1038_ (.A1(_0245_),
    .A2(_0393_),
    .ZN(_0394_));
 MUX2_X1 _1039_ (.A(\mem[1][7] ),
    .B(\mem[5][7] ),
    .S(_0280_),
    .Z(_0395_));
 INV_X1 _1040_ (.A(_0395_),
    .ZN(_0396_));
 AOI21_X1 _1041_ (.A(_0394_),
    .B1(_0396_),
    .B2(_0248_),
    .ZN(_0397_));
 MUX2_X1 _1042_ (.A(\mem[0][7] ),
    .B(\mem[4][7] ),
    .S(_0260_),
    .Z(_0398_));
 NOR2_X1 _1043_ (.A1(_0256_),
    .A2(_0398_),
    .ZN(_0399_));
 MUX2_X1 _1044_ (.A(\mem[2][7] ),
    .B(\mem[6][7] ),
    .S(_0271_),
    .Z(_0400_));
 NOR3_X1 _1045_ (.A1(_0258_),
    .A2(_0259_),
    .A3(_0400_),
    .ZN(_0401_));
 NOR3_X1 _1046_ (.A1(_0252_),
    .A2(_0399_),
    .A3(_0401_),
    .ZN(_0402_));
 MUX2_X1 _1047_ (.A(\mem[9][7] ),
    .B(\mem[13][7] ),
    .S(_0239_),
    .Z(_0403_));
 MUX2_X1 _1048_ (.A(\mem[11][7] ),
    .B(\mem[15][7] ),
    .S(_0265_),
    .Z(_0404_));
 MUX2_X1 _1049_ (.A(_0403_),
    .B(_0404_),
    .S(_0267_),
    .Z(_0405_));
 MUX2_X1 _1050_ (.A(\mem[8][7] ),
    .B(\mem[12][7] ),
    .S(_0265_),
    .Z(_0406_));
 MUX2_X1 _1051_ (.A(\mem[10][7] ),
    .B(\mem[14][7] ),
    .S(_0269_),
    .Z(_0407_));
 MUX2_X1 _1052_ (.A(_0406_),
    .B(_0407_),
    .S(_0267_),
    .Z(_0408_));
 MUX2_X1 _1053_ (.A(_0405_),
    .B(_0408_),
    .S(_0247_),
    .Z(_0409_));
 AOI221_X1 _1054_ (.A(_0236_),
    .B1(_0397_),
    .B2(_0402_),
    .C1(_0409_),
    .C2(_0253_),
    .ZN(_0410_));
 INV_X1 _1055_ (.A(net23),
    .ZN(_0411_));
 AOI21_X1 _1056_ (.A(_0410_),
    .B1(_0276_),
    .B2(_0411_),
    .ZN(_0141_));
 MUX2_X1 _1057_ (.A(_0004_),
    .B(_0258_),
    .S(_0276_),
    .Z(_0142_));
 MUX2_X1 _1058_ (.A(_0005_),
    .B(_0244_),
    .S(_0276_),
    .Z(_0143_));
 XNOR2_X2 _1059_ (.A(_0643_),
    .B(_0624_),
    .ZN(_0412_));
 MUX2_X1 _1060_ (.A(_0412_),
    .B(_0280_),
    .S(_0237_),
    .Z(_0144_));
 NAND3_X1 _1061_ (.A1(_0242_),
    .A2(_0244_),
    .A3(_0280_),
    .ZN(_0413_));
 XOR2_X2 _1062_ (.A(_0620_),
    .B(_0413_),
    .Z(_0414_));
 MUX2_X1 _1063_ (.A(_0414_),
    .B(_0253_),
    .S(_0237_),
    .Z(_0145_));
 XNOR2_X1 _1064_ (.A(_0258_),
    .B(_0005_),
    .ZN(_0415_));
 MUX2_X1 _1065_ (.A(_0415_),
    .B(\rd_ptr_gray[0] ),
    .S(_0237_),
    .Z(_0146_));
 XOR2_X1 _1066_ (.A(_0005_),
    .B(_0412_),
    .Z(_0416_));
 MUX2_X1 _1067_ (.A(_0416_),
    .B(\rd_ptr_gray[1] ),
    .S(_0237_),
    .Z(_0147_));
 XOR2_X1 _1068_ (.A(_0412_),
    .B(_0414_),
    .Z(_0417_));
 MUX2_X1 _1069_ (.A(_0417_),
    .B(\rd_ptr_gray[2] ),
    .S(_0237_),
    .Z(_0148_));
 NAND3_X1 _1070_ (.A1(_0280_),
    .A2(_0252_),
    .A3(_0643_),
    .ZN(_0418_));
 XOR2_X1 _1071_ (.A(\rd_ptr_bin[4] ),
    .B(_0418_),
    .Z(_0419_));
 XNOR2_X1 _1072_ (.A(_0414_),
    .B(_0419_),
    .ZN(_0420_));
 MUX2_X1 _1073_ (.A(_0420_),
    .B(\rd_ptr_gray[3] ),
    .S(_0237_),
    .Z(_0149_));
 NOR2_X1 _1074_ (.A1(_0237_),
    .A2(_0418_),
    .ZN(_0421_));
 XOR2_X1 _1075_ (.A(\rd_ptr_bin[4] ),
    .B(_0421_),
    .Z(_0150_));
 MUX2_X1 _1076_ (.A(\wr_ptr_bin[0] ),
    .B(_0002_),
    .S(_0210_),
    .Z(_0151_));
 MUX2_X1 _1077_ (.A(\wr_ptr_bin[1] ),
    .B(_0003_),
    .S(_0210_),
    .Z(_0152_));
 OR2_X1 _1078_ (.A1(_0185_),
    .A2(_0210_),
    .ZN(_0422_));
 XOR2_X2 _1079_ (.A(_0206_),
    .B(_0001_),
    .Z(_0423_));
 NAND2_X1 _1080_ (.A1(net5),
    .A2(_0167_),
    .ZN(_0424_));
 OAI21_X1 _1081_ (.A(_0422_),
    .B1(_0423_),
    .B2(_0424_),
    .ZN(_0153_));
 NAND3_X1 _1082_ (.A1(\wr_ptr_bin[2] ),
    .A2(\wr_ptr_bin[1] ),
    .A3(\wr_ptr_bin[0] ),
    .ZN(_0425_));
 XOR2_X2 _1083_ (.A(_0000_),
    .B(_0425_),
    .Z(_0426_));
 MUX2_X1 _1084_ (.A(_0183_),
    .B(_0426_),
    .S(_0210_),
    .Z(_0154_));
 XNOR2_X1 _1085_ (.A(\wr_ptr_bin[0] ),
    .B(_0003_),
    .ZN(_0427_));
 MUX2_X1 _1086_ (.A(\wr_ptr_gray[0] ),
    .B(_0427_),
    .S(_0210_),
    .Z(_0155_));
 XNOR2_X1 _1087_ (.A(_0003_),
    .B(_0423_),
    .ZN(_0428_));
 MUX2_X1 _1088_ (.A(\wr_ptr_gray[1] ),
    .B(_0428_),
    .S(_0210_),
    .Z(_0156_));
 XNOR2_X1 _1089_ (.A(_0423_),
    .B(_0426_),
    .ZN(_0429_));
 MUX2_X1 _1090_ (.A(\wr_ptr_gray[2] ),
    .B(_0429_),
    .S(_0210_),
    .Z(_0157_));
 NAND2_X1 _1091_ (.A1(_0206_),
    .A2(_0212_),
    .ZN(_0430_));
 XOR2_X1 _1092_ (.A(\wr_ptr_bin[4] ),
    .B(_0430_),
    .Z(_0431_));
 XNOR2_X1 _1093_ (.A(_0426_),
    .B(_0431_),
    .ZN(_0432_));
 MUX2_X1 _1094_ (.A(\wr_ptr_gray[3] ),
    .B(_0432_),
    .S(_0210_),
    .Z(_0158_));
 XNOR2_X1 _1095_ (.A(\wr_ptr_bin[4] ),
    .B(_0216_),
    .ZN(_0159_));
 NAND2_X1 _1096_ (.A1(_0169_),
    .A2(_0170_),
    .ZN(_0433_));
 NAND2_X1 _1097_ (.A1(_0171_),
    .A2(_0172_),
    .ZN(_0434_));
 XNOR2_X1 _1098_ (.A(_0619_),
    .B(_0627_),
    .ZN(net12));
 OR2_X1 _1099_ (.A1(net11),
    .A2(net10),
    .ZN(_0435_));
 AND2_X1 _1100_ (.A1(net12),
    .A2(_0435_),
    .ZN(_0436_));
 OAI33_X1 _1101_ (.A1(_0433_),
    .A2(_0168_),
    .A3(_0434_),
    .B1(net13),
    .B2(net14),
    .B3(_0436_),
    .ZN(net7));
 XNOR2_X1 _1102_ (.A(_0637_),
    .B(_0615_),
    .ZN(_0437_));
 INV_X1 _1103_ (.A(_0636_),
    .ZN(_0438_));
 AOI21_X1 _1104_ (.A(_0638_),
    .B1(_0639_),
    .B2(_0613_),
    .ZN(_0439_));
 INV_X1 _1105_ (.A(_0637_),
    .ZN(_0440_));
 OAI21_X1 _1106_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0440_),
    .ZN(_0441_));
 XNOR2_X1 _1107_ (.A(_0634_),
    .B(_0441_),
    .ZN(_0442_));
 AOI21_X1 _1108_ (.A(_0636_),
    .B1(_0615_),
    .B2(_0637_),
    .ZN(_0443_));
 INV_X1 _1109_ (.A(_0443_),
    .ZN(_0444_));
 AOI21_X1 _1110_ (.A(_0633_),
    .B1(_0444_),
    .B2(_0634_),
    .ZN(_0445_));
 XOR2_X1 _1111_ (.A(_0164_),
    .B(_0445_),
    .Z(_0446_));
 NAND4_X1 _1112_ (.A1(_0167_),
    .A2(_0437_),
    .A3(_0442_),
    .A4(_0446_),
    .ZN(net8));
 FA_X1 _1113_ (.A(\wr_ptr_bin[1] ),
    .B(_0613_),
    .CI(_0614_),
    .CO(_0615_),
    .S(_0616_));
 FA_X1 _1114_ (.A(\rd_ptr_bin[1] ),
    .B(_0617_),
    .CI(_0618_),
    .CO(_0619_),
    .S(net11));
 HA_X1 _1115_ (.A(_0620_),
    .B(_0621_),
    .CO(_0622_),
    .S(_0623_));
 HA_X1 _1116_ (.A(_0624_),
    .B(_0625_),
    .CO(_0626_),
    .S(_0627_));
 HA_X1 _1117_ (.A(_0628_),
    .B(_0629_),
    .CO(_0630_),
    .S(_0631_));
 HA_X1 _1118_ (.A(\wr_ptr_bin[3] ),
    .B(_0632_),
    .CO(_0633_),
    .S(_0634_));
 HA_X1 _1119_ (.A(\wr_ptr_bin[2] ),
    .B(_0635_),
    .CO(_0636_),
    .S(_0637_));
 HA_X1 _1120_ (.A(\wr_ptr_bin[1] ),
    .B(_0614_),
    .CO(_0638_),
    .S(_0639_));
 HA_X1 _1121_ (.A(_0002_),
    .B(_0640_),
    .CO(_0641_),
    .S(_0642_));
 HA_X1 _1122_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .CO(_0643_),
    .S(_0005_));
 HA_X1 _1123_ (.A(_0002_),
    .B(_0644_),
    .CO(_0645_),
    .S(_0003_));
 HA_X1 _1124_ (.A(_0002_),
    .B(\wr_ptr_bin[1] ),
    .CO(_0646_),
    .S(_0647_));
 HA_X1 _1125_ (.A(\wr_ptr_bin[0] ),
    .B(_0644_),
    .CO(_0648_),
    .S(_0649_));
 HA_X1 _1126_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .CO(_0650_),
    .S(_0651_));
 HA_X1 _1127_ (.A(\rd_ptr_bin[0] ),
    .B(_0652_),
    .CO(_0617_),
    .S(_0653_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0006_),
    .CK(net4),
    .Q(\mem[0][0] ),
    .QN(_0592_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0007_),
    .CK(net4),
    .Q(\mem[0][1] ),
    .QN(_0591_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0008_),
    .CK(net4),
    .Q(\mem[0][2] ),
    .QN(_0590_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0009_),
    .CK(net4),
    .Q(\mem[0][3] ),
    .QN(_0589_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0010_),
    .CK(net4),
    .Q(\mem[0][4] ),
    .QN(_0588_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0011_),
    .CK(net4),
    .Q(\mem[0][5] ),
    .QN(_0587_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0012_),
    .CK(net4),
    .Q(\mem[0][6] ),
    .QN(_0586_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0013_),
    .CK(net4),
    .Q(\mem[0][7] ),
    .QN(_0585_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0014_),
    .CK(net4),
    .Q(\mem[10][0] ),
    .QN(_0584_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0015_),
    .CK(net4),
    .Q(\mem[10][1] ),
    .QN(_0583_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0016_),
    .CK(net4),
    .Q(\mem[10][2] ),
    .QN(_0582_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0017_),
    .CK(net4),
    .Q(\mem[10][3] ),
    .QN(_0581_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0018_),
    .CK(net4),
    .Q(\mem[10][4] ),
    .QN(_0580_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0019_),
    .CK(net4),
    .Q(\mem[10][5] ),
    .QN(_0579_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0020_),
    .CK(net4),
    .Q(\mem[10][6] ),
    .QN(_0578_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0021_),
    .CK(net4),
    .Q(\mem[10][7] ),
    .QN(_0577_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0022_),
    .CK(net4),
    .Q(\mem[11][0] ),
    .QN(_0576_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0023_),
    .CK(net4),
    .Q(\mem[11][1] ),
    .QN(_0575_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0024_),
    .CK(net4),
    .Q(\mem[11][2] ),
    .QN(_0574_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0025_),
    .CK(net4),
    .Q(\mem[11][3] ),
    .QN(_0573_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0026_),
    .CK(net4),
    .Q(\mem[11][4] ),
    .QN(_0572_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0027_),
    .CK(net4),
    .Q(\mem[11][5] ),
    .QN(_0571_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0028_),
    .CK(net4),
    .Q(\mem[11][6] ),
    .QN(_0570_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0029_),
    .CK(net4),
    .Q(\mem[11][7] ),
    .QN(_0569_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0030_),
    .CK(net4),
    .Q(\mem[12][0] ),
    .QN(_0568_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0031_),
    .CK(net4),
    .Q(\mem[12][1] ),
    .QN(_0567_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0032_),
    .CK(net4),
    .Q(\mem[12][2] ),
    .QN(_0566_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0033_),
    .CK(net4),
    .Q(\mem[12][3] ),
    .QN(_0565_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0034_),
    .CK(net4),
    .Q(\mem[12][4] ),
    .QN(_0564_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0035_),
    .CK(net4),
    .Q(\mem[12][5] ),
    .QN(_0563_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0036_),
    .CK(net4),
    .Q(\mem[12][6] ),
    .QN(_0562_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0037_),
    .CK(net4),
    .Q(\mem[12][7] ),
    .QN(_0561_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0038_),
    .CK(net4),
    .Q(\mem[13][0] ),
    .QN(_0560_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0039_),
    .CK(net4),
    .Q(\mem[13][1] ),
    .QN(_0559_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0040_),
    .CK(net4),
    .Q(\mem[13][2] ),
    .QN(_0558_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0041_),
    .CK(net4),
    .Q(\mem[13][3] ),
    .QN(_0557_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0042_),
    .CK(net4),
    .Q(\mem[13][4] ),
    .QN(_0556_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0043_),
    .CK(net4),
    .Q(\mem[13][5] ),
    .QN(_0555_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0044_),
    .CK(net4),
    .Q(\mem[13][6] ),
    .QN(_0554_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0045_),
    .CK(net4),
    .Q(\mem[13][7] ),
    .QN(_0553_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0046_),
    .CK(net4),
    .Q(\mem[14][0] ),
    .QN(_0552_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0047_),
    .CK(net4),
    .Q(\mem[14][1] ),
    .QN(_0551_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0048_),
    .CK(net4),
    .Q(\mem[14][2] ),
    .QN(_0550_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0049_),
    .CK(net4),
    .Q(\mem[14][3] ),
    .QN(_0549_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0050_),
    .CK(net4),
    .Q(\mem[14][4] ),
    .QN(_0548_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0051_),
    .CK(net4),
    .Q(\mem[14][5] ),
    .QN(_0547_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0052_),
    .CK(net4),
    .Q(\mem[14][6] ),
    .QN(_0546_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0053_),
    .CK(net4),
    .Q(\mem[14][7] ),
    .QN(_0545_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0054_),
    .CK(net4),
    .Q(\mem[15][0] ),
    .QN(_0544_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0055_),
    .CK(net4),
    .Q(\mem[15][1] ),
    .QN(_0543_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0056_),
    .CK(net4),
    .Q(\mem[15][2] ),
    .QN(_0542_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0057_),
    .CK(net4),
    .Q(\mem[15][3] ),
    .QN(_0541_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0058_),
    .CK(net4),
    .Q(\mem[15][4] ),
    .QN(_0540_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0059_),
    .CK(net4),
    .Q(\mem[15][5] ),
    .QN(_0539_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0060_),
    .CK(net4),
    .Q(\mem[15][6] ),
    .QN(_0538_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0061_),
    .CK(net4),
    .Q(\mem[15][7] ),
    .QN(_0537_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0062_),
    .CK(net4),
    .Q(\mem[1][0] ),
    .QN(_0536_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0063_),
    .CK(net4),
    .Q(\mem[1][1] ),
    .QN(_0535_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0064_),
    .CK(net4),
    .Q(\mem[1][2] ),
    .QN(_0534_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0065_),
    .CK(net4),
    .Q(\mem[1][3] ),
    .QN(_0533_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0066_),
    .CK(net4),
    .Q(\mem[1][4] ),
    .QN(_0532_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0067_),
    .CK(net4),
    .Q(\mem[1][5] ),
    .QN(_0531_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0068_),
    .CK(net4),
    .Q(\mem[1][6] ),
    .QN(_0530_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0069_),
    .CK(net4),
    .Q(\mem[1][7] ),
    .QN(_0529_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0070_),
    .CK(net4),
    .Q(\mem[2][0] ),
    .QN(_0528_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0071_),
    .CK(net4),
    .Q(\mem[2][1] ),
    .QN(_0527_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0072_),
    .CK(net4),
    .Q(\mem[2][2] ),
    .QN(_0526_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0073_),
    .CK(net4),
    .Q(\mem[2][3] ),
    .QN(_0525_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0074_),
    .CK(net4),
    .Q(\mem[2][4] ),
    .QN(_0524_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0075_),
    .CK(net4),
    .Q(\mem[2][5] ),
    .QN(_0523_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0076_),
    .CK(net4),
    .Q(\mem[2][6] ),
    .QN(_0522_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0077_),
    .CK(net4),
    .Q(\mem[2][7] ),
    .QN(_0521_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0078_),
    .CK(net4),
    .Q(\mem[3][0] ),
    .QN(_0520_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0079_),
    .CK(net4),
    .Q(\mem[3][1] ),
    .QN(_0519_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0080_),
    .CK(net4),
    .Q(\mem[3][2] ),
    .QN(_0518_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0081_),
    .CK(net4),
    .Q(\mem[3][3] ),
    .QN(_0517_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0082_),
    .CK(net4),
    .Q(\mem[3][4] ),
    .QN(_0516_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0083_),
    .CK(net4),
    .Q(\mem[3][5] ),
    .QN(_0515_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0084_),
    .CK(net4),
    .Q(\mem[3][6] ),
    .QN(_0514_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0085_),
    .CK(net4),
    .Q(\mem[3][7] ),
    .QN(_0513_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0086_),
    .CK(net4),
    .Q(\mem[4][0] ),
    .QN(_0512_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0087_),
    .CK(net4),
    .Q(\mem[4][1] ),
    .QN(_0511_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0088_),
    .CK(net4),
    .Q(\mem[4][2] ),
    .QN(_0510_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0089_),
    .CK(net4),
    .Q(\mem[4][3] ),
    .QN(_0509_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0090_),
    .CK(net4),
    .Q(\mem[4][4] ),
    .QN(_0508_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0091_),
    .CK(net4),
    .Q(\mem[4][5] ),
    .QN(_0507_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0092_),
    .CK(net4),
    .Q(\mem[4][6] ),
    .QN(_0506_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0093_),
    .CK(net4),
    .Q(\mem[4][7] ),
    .QN(_0505_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0094_),
    .CK(net4),
    .Q(\mem[5][0] ),
    .QN(_0504_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0095_),
    .CK(net4),
    .Q(\mem[5][1] ),
    .QN(_0503_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0096_),
    .CK(net4),
    .Q(\mem[5][2] ),
    .QN(_0502_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0097_),
    .CK(net4),
    .Q(\mem[5][3] ),
    .QN(_0501_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0098_),
    .CK(net4),
    .Q(\mem[5][4] ),
    .QN(_0500_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0099_),
    .CK(net4),
    .Q(\mem[5][5] ),
    .QN(_0499_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0100_),
    .CK(net4),
    .Q(\mem[5][6] ),
    .QN(_0498_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0101_),
    .CK(net4),
    .Q(\mem[5][7] ),
    .QN(_0497_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0102_),
    .CK(net4),
    .Q(\mem[6][0] ),
    .QN(_0496_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0103_),
    .CK(net4),
    .Q(\mem[6][1] ),
    .QN(_0495_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0104_),
    .CK(net4),
    .Q(\mem[6][2] ),
    .QN(_0494_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0105_),
    .CK(net4),
    .Q(\mem[6][3] ),
    .QN(_0493_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0106_),
    .CK(net4),
    .Q(\mem[6][4] ),
    .QN(_0492_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0107_),
    .CK(net4),
    .Q(\mem[6][5] ),
    .QN(_0491_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0108_),
    .CK(net4),
    .Q(\mem[6][6] ),
    .QN(_0490_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0109_),
    .CK(net4),
    .Q(\mem[6][7] ),
    .QN(_0489_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0110_),
    .CK(net4),
    .Q(\mem[7][0] ),
    .QN(_0488_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0111_),
    .CK(net4),
    .Q(\mem[7][1] ),
    .QN(_0487_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0112_),
    .CK(net4),
    .Q(\mem[7][2] ),
    .QN(_0486_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0113_),
    .CK(net4),
    .Q(\mem[7][3] ),
    .QN(_0485_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0114_),
    .CK(net4),
    .Q(\mem[7][4] ),
    .QN(_0484_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0115_),
    .CK(net4),
    .Q(\mem[7][5] ),
    .QN(_0483_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0116_),
    .CK(net4),
    .Q(\mem[7][6] ),
    .QN(_0482_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0117_),
    .CK(net4),
    .Q(\mem[7][7] ),
    .QN(_0481_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0118_),
    .CK(net4),
    .Q(\mem[8][0] ),
    .QN(_0480_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0119_),
    .CK(net4),
    .Q(\mem[8][1] ),
    .QN(_0479_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0120_),
    .CK(net4),
    .Q(\mem[8][2] ),
    .QN(_0478_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0121_),
    .CK(net4),
    .Q(\mem[8][3] ),
    .QN(_0477_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0122_),
    .CK(net4),
    .Q(\mem[8][4] ),
    .QN(_0476_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0123_),
    .CK(net4),
    .Q(\mem[8][5] ),
    .QN(_0475_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0124_),
    .CK(net4),
    .Q(\mem[8][6] ),
    .QN(_0474_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0125_),
    .CK(net4),
    .Q(\mem[8][7] ),
    .QN(_0473_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0126_),
    .CK(net4),
    .Q(\mem[9][0] ),
    .QN(_0472_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0127_),
    .CK(net4),
    .Q(\mem[9][1] ),
    .QN(_0471_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0128_),
    .CK(net4),
    .Q(\mem[9][2] ),
    .QN(_0470_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0129_),
    .CK(net4),
    .Q(\mem[9][3] ),
    .QN(_0469_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0130_),
    .CK(net4),
    .Q(\mem[9][4] ),
    .QN(_0468_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0131_),
    .CK(net4),
    .Q(\mem[9][5] ),
    .QN(_0467_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0132_),
    .CK(net4),
    .Q(\mem[9][6] ),
    .QN(_0466_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0133_),
    .CK(net4),
    .Q(\mem[9][7] ),
    .QN(_0465_));
 DFF_X1 \rd_data_reg[0]$_DFFE_PP_  (.D(_0134_),
    .CK(net1),
    .Q(net16),
    .QN(_0464_));
 DFF_X1 \rd_data_reg[1]$_DFFE_PP_  (.D(_0135_),
    .CK(net1),
    .Q(net17),
    .QN(_0463_));
 DFF_X1 \rd_data_reg[2]$_DFFE_PP_  (.D(_0136_),
    .CK(net1),
    .Q(net18),
    .QN(_0462_));
 DFF_X1 \rd_data_reg[3]$_DFFE_PP_  (.D(_0137_),
    .CK(net1),
    .Q(net19),
    .QN(_0461_));
 DFF_X1 \rd_data_reg[4]$_DFFE_PP_  (.D(_0138_),
    .CK(net1),
    .Q(net20),
    .QN(_0460_));
 DFF_X1 \rd_data_reg[5]$_DFFE_PP_  (.D(_0139_),
    .CK(net1),
    .Q(net21),
    .QN(_0459_));
 DFF_X1 \rd_data_reg[6]$_DFFE_PP_  (.D(_0140_),
    .CK(net1),
    .Q(net22),
    .QN(_0458_));
 DFF_X1 \rd_data_reg[7]$_DFFE_PP_  (.D(_0141_),
    .CK(net1),
    .Q(net23),
    .QN(_0457_));
 DFFR_X1 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_0142_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[0] ),
    .QN(_0004_));
 DFFR_X2 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_0143_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[1] ),
    .QN(_0628_));
 DFFR_X1 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_0144_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[2] ),
    .QN(_0624_));
 DFFR_X2 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_0145_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[3] ),
    .QN(_0620_));
 DFFR_X1 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_0146_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[0] ),
    .QN(_0456_));
 DFFR_X1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_0147_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[1] ),
    .QN(_0455_));
 DFFR_X2 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_0148_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[2] ),
    .QN(_0454_));
 DFFR_X1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_0149_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[3] ),
    .QN(_0453_));
 DFFR_X2 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_0150_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[4] ),
    .QN(_0593_));
 DFFR_X1 \rd_ptr_gray_wr_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync1[0] ),
    .QN(_0594_));
 DFFR_X1 \rd_ptr_gray_wr_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync1[1] ),
    .QN(_0595_));
 DFFR_X1 \rd_ptr_gray_wr_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync1[2] ),
    .QN(_0596_));
 DFFR_X1 \rd_ptr_gray_wr_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync1[3] ),
    .QN(_0597_));
 DFFR_X1 \rd_ptr_gray_wr_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync1[4] ),
    .QN(_0598_));
 DFFR_X1 \rd_ptr_gray_wr_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[0] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync2[0] ),
    .QN(_0599_));
 DFFR_X2 \rd_ptr_gray_wr_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[1] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync2[1] ),
    .QN(_0600_));
 DFFR_X2 \rd_ptr_gray_wr_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[2] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync2[2] ),
    .QN(_0601_));
 DFFR_X2 \rd_ptr_gray_wr_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[3] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_wr_sync2[3] ),
    .QN(_0602_));
 DFFR_X2 \rd_ptr_gray_wr_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[4] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_bin_wr_sync[4] ),
    .QN(_0452_));
 DFFR_X2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_0151_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[0] ),
    .QN(_0002_));
 DFFR_X2 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_0152_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[1] ),
    .QN(_0644_));
 DFFR_X2 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_0153_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[2] ),
    .QN(_0001_));
 DFFR_X1 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_0154_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[3] ),
    .QN(_0000_));
 DFFR_X2 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_0155_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[0] ),
    .QN(_0451_));
 DFFR_X1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_0156_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[1] ),
    .QN(_0450_));
 DFFR_X1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_0157_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[2] ),
    .QN(_0449_));
 DFFR_X1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_0158_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[3] ),
    .QN(_0448_));
 DFFR_X2 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_0159_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[4] ),
    .QN(_0603_));
 DFFR_X1 \wr_ptr_gray_rd_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync1[0] ),
    .QN(_0604_));
 DFFR_X1 \wr_ptr_gray_rd_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync1[1] ),
    .QN(_0605_));
 DFFR_X1 \wr_ptr_gray_rd_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync1[2] ),
    .QN(_0606_));
 DFFR_X1 \wr_ptr_gray_rd_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync1[3] ),
    .QN(_0607_));
 DFFR_X1 \wr_ptr_gray_rd_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync1[4] ),
    .QN(_0608_));
 DFFR_X1 \wr_ptr_gray_rd_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync2[0] ),
    .QN(_0609_));
 DFFR_X1 \wr_ptr_gray_rd_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync2[1] ),
    .QN(_0610_));
 DFFR_X2 \wr_ptr_gray_rd_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync2[2] ),
    .QN(_0611_));
 DFFR_X1 \wr_ptr_gray_rd_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_rd_sync2[3] ),
    .QN(_0612_));
 DFFR_X2 \wr_ptr_gray_rd_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_bin_rd_sync[4] ),
    .QN(_0447_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_77 ();
 BUF_X4 input1 (.A(rd_clk),
    .Z(net1));
 BUF_X1 input2 (.A(rd_en),
    .Z(net2));
 BUF_X4 input3 (.A(rd_rst_n),
    .Z(net3));
 BUF_X16 input4 (.A(wr_clk),
    .Z(net4));
 CLKBUF_X2 input5 (.A(wr_en),
    .Z(net5));
 BUF_X4 input6 (.A(wr_rst_n),
    .Z(net6));
 BUF_X1 output7 (.A(net7),
    .Z(almost_empty));
 BUF_X1 output8 (.A(net8),
    .Z(almost_full));
 BUF_X1 output9 (.A(net9),
    .Z(empty));
 BUF_X1 output10 (.A(net10),
    .Z(fifo_count[0]));
 BUF_X1 output11 (.A(net11),
    .Z(fifo_count[1]));
 BUF_X1 output12 (.A(net12),
    .Z(fifo_count[2]));
 BUF_X1 output13 (.A(net13),
    .Z(fifo_count[3]));
 BUF_X1 output14 (.A(net14),
    .Z(fifo_count[4]));
 BUF_X1 output15 (.A(net15),
    .Z(full));
 BUF_X1 output16 (.A(net16),
    .Z(rd_data[0]));
 BUF_X1 output17 (.A(net17),
    .Z(rd_data[1]));
 BUF_X1 output18 (.A(net18),
    .Z(rd_data[2]));
 BUF_X1 output19 (.A(net19),
    .Z(rd_data[3]));
 BUF_X1 output20 (.A(net20),
    .Z(rd_data[4]));
 BUF_X1 output21 (.A(net21),
    .Z(rd_data[5]));
 BUF_X1 output22 (.A(net22),
    .Z(rd_data[6]));
 BUF_X1 output23 (.A(net23),
    .Z(rd_data[7]));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_17 ();
 FILLCELL_X4 FILLER_0_25 ();
 FILLCELL_X2 FILLER_0_29 ();
 FILLCELL_X1 FILLER_0_31 ();
 FILLCELL_X16 FILLER_0_36 ();
 FILLCELL_X8 FILLER_0_52 ();
 FILLCELL_X2 FILLER_0_60 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_81 ();
 FILLCELL_X16 FILLER_0_92 ();
 FILLCELL_X8 FILLER_0_108 ();
 FILLCELL_X8 FILLER_0_147 ();
 FILLCELL_X2 FILLER_0_155 ();
 FILLCELL_X1 FILLER_0_157 ();
 FILLCELL_X8 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_186 ();
 FILLCELL_X4 FILLER_0_218 ();
 FILLCELL_X2 FILLER_0_222 ();
 FILLCELL_X32 FILLER_0_233 ();
 FILLCELL_X16 FILLER_0_265 ();
 FILLCELL_X8 FILLER_0_281 ();
 FILLCELL_X4 FILLER_0_289 ();
 FILLCELL_X1 FILLER_0_293 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X16 FILLER_1_33 ();
 FILLCELL_X8 FILLER_1_49 ();
 FILLCELL_X1 FILLER_1_57 ();
 FILLCELL_X1 FILLER_1_82 ();
 FILLCELL_X1 FILLER_1_117 ();
 FILLCELL_X16 FILLER_1_142 ();
 FILLCELL_X8 FILLER_1_158 ();
 FILLCELL_X16 FILLER_1_183 ();
 FILLCELL_X1 FILLER_1_232 ();
 FILLCELL_X32 FILLER_1_253 ();
 FILLCELL_X8 FILLER_1_285 ();
 FILLCELL_X1 FILLER_1_293 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X4 FILLER_2_33 ();
 FILLCELL_X1 FILLER_2_37 ();
 FILLCELL_X8 FILLER_2_79 ();
 FILLCELL_X4 FILLER_2_87 ();
 FILLCELL_X1 FILLER_2_91 ();
 FILLCELL_X4 FILLER_2_113 ();
 FILLCELL_X2 FILLER_2_117 ();
 FILLCELL_X1 FILLER_2_119 ();
 FILLCELL_X4 FILLER_2_127 ();
 FILLCELL_X2 FILLER_2_131 ();
 FILLCELL_X1 FILLER_2_133 ();
 FILLCELL_X4 FILLER_2_158 ();
 FILLCELL_X2 FILLER_2_162 ();
 FILLCELL_X8 FILLER_2_185 ();
 FILLCELL_X4 FILLER_2_193 ();
 FILLCELL_X2 FILLER_2_197 ();
 FILLCELL_X1 FILLER_2_199 ();
 FILLCELL_X2 FILLER_2_228 ();
 FILLCELL_X32 FILLER_2_237 ();
 FILLCELL_X16 FILLER_2_269 ();
 FILLCELL_X2 FILLER_2_292 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X4 FILLER_3_49 ();
 FILLCELL_X2 FILLER_3_53 ();
 FILLCELL_X8 FILLER_3_69 ();
 FILLCELL_X8 FILLER_3_84 ();
 FILLCELL_X2 FILLER_3_92 ();
 FILLCELL_X8 FILLER_3_111 ();
 FILLCELL_X4 FILLER_3_119 ();
 FILLCELL_X2 FILLER_3_123 ();
 FILLCELL_X4 FILLER_3_142 ();
 FILLCELL_X1 FILLER_3_146 ();
 FILLCELL_X32 FILLER_3_154 ();
 FILLCELL_X8 FILLER_3_186 ();
 FILLCELL_X4 FILLER_3_194 ();
 FILLCELL_X8 FILLER_3_215 ();
 FILLCELL_X2 FILLER_3_223 ();
 FILLCELL_X32 FILLER_3_254 ();
 FILLCELL_X8 FILLER_3_286 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_25 ();
 FILLCELL_X2 FILLER_4_29 ();
 FILLCELL_X8 FILLER_4_48 ();
 FILLCELL_X1 FILLER_4_56 ();
 FILLCELL_X16 FILLER_4_81 ();
 FILLCELL_X16 FILLER_4_114 ();
 FILLCELL_X8 FILLER_4_130 ();
 FILLCELL_X2 FILLER_4_138 ();
 FILLCELL_X16 FILLER_4_147 ();
 FILLCELL_X4 FILLER_4_197 ();
 FILLCELL_X16 FILLER_4_221 ();
 FILLCELL_X2 FILLER_4_237 ();
 FILLCELL_X1 FILLER_4_239 ();
 FILLCELL_X32 FILLER_4_252 ();
 FILLCELL_X8 FILLER_4_284 ();
 FILLCELL_X2 FILLER_4_292 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X2 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_59 ();
 FILLCELL_X4 FILLER_5_105 ();
 FILLCELL_X2 FILLER_5_109 ();
 FILLCELL_X1 FILLER_5_111 ();
 FILLCELL_X8 FILLER_5_119 ();
 FILLCELL_X4 FILLER_5_127 ();
 FILLCELL_X1 FILLER_5_131 ();
 FILLCELL_X16 FILLER_5_149 ();
 FILLCELL_X4 FILLER_5_165 ();
 FILLCELL_X1 FILLER_5_169 ();
 FILLCELL_X8 FILLER_5_191 ();
 FILLCELL_X4 FILLER_5_199 ();
 FILLCELL_X2 FILLER_5_203 ();
 FILLCELL_X1 FILLER_5_205 ();
 FILLCELL_X4 FILLER_5_216 ();
 FILLCELL_X8 FILLER_5_224 ();
 FILLCELL_X4 FILLER_5_232 ();
 FILLCELL_X2 FILLER_5_236 ();
 FILLCELL_X16 FILLER_5_270 ();
 FILLCELL_X8 FILLER_5_286 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_9 ();
 FILLCELL_X4 FILLER_6_34 ();
 FILLCELL_X1 FILLER_6_38 ();
 FILLCELL_X4 FILLER_6_53 ();
 FILLCELL_X1 FILLER_6_57 ();
 FILLCELL_X16 FILLER_6_82 ();
 FILLCELL_X4 FILLER_6_98 ();
 FILLCELL_X16 FILLER_6_109 ();
 FILLCELL_X8 FILLER_6_125 ();
 FILLCELL_X1 FILLER_6_133 ();
 FILLCELL_X2 FILLER_6_141 ();
 FILLCELL_X1 FILLER_6_143 ();
 FILLCELL_X4 FILLER_6_158 ();
 FILLCELL_X2 FILLER_6_162 ();
 FILLCELL_X1 FILLER_6_164 ();
 FILLCELL_X2 FILLER_6_172 ();
 FILLCELL_X16 FILLER_6_191 ();
 FILLCELL_X4 FILLER_6_211 ();
 FILLCELL_X1 FILLER_6_215 ();
 FILLCELL_X4 FILLER_6_229 ();
 FILLCELL_X2 FILLER_6_233 ();
 FILLCELL_X1 FILLER_6_235 ();
 FILLCELL_X2 FILLER_6_242 ();
 FILLCELL_X2 FILLER_6_248 ();
 FILLCELL_X1 FILLER_6_250 ();
 FILLCELL_X4 FILLER_6_253 ();
 FILLCELL_X2 FILLER_6_257 ();
 FILLCELL_X4 FILLER_6_263 ();
 FILLCELL_X1 FILLER_6_267 ();
 FILLCELL_X4 FILLER_6_288 ();
 FILLCELL_X2 FILLER_6_292 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_34 ();
 FILLCELL_X4 FILLER_7_42 ();
 FILLCELL_X1 FILLER_7_46 ();
 FILLCELL_X1 FILLER_7_54 ();
 FILLCELL_X4 FILLER_7_59 ();
 FILLCELL_X2 FILLER_7_63 ();
 FILLCELL_X1 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_90 ();
 FILLCELL_X1 FILLER_7_98 ();
 FILLCELL_X32 FILLER_7_116 ();
 FILLCELL_X2 FILLER_7_148 ();
 FILLCELL_X8 FILLER_7_167 ();
 FILLCELL_X1 FILLER_7_175 ();
 FILLCELL_X8 FILLER_7_194 ();
 FILLCELL_X1 FILLER_7_202 ();
 FILLCELL_X2 FILLER_7_228 ();
 FILLCELL_X4 FILLER_7_249 ();
 FILLCELL_X4 FILLER_7_266 ();
 FILLCELL_X2 FILLER_7_270 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_17 ();
 FILLCELL_X2 FILLER_8_26 ();
 FILLCELL_X4 FILLER_8_35 ();
 FILLCELL_X2 FILLER_8_39 ();
 FILLCELL_X8 FILLER_8_58 ();
 FILLCELL_X2 FILLER_8_66 ();
 FILLCELL_X1 FILLER_8_68 ();
 FILLCELL_X4 FILLER_8_76 ();
 FILLCELL_X1 FILLER_8_80 ();
 FILLCELL_X8 FILLER_8_88 ();
 FILLCELL_X2 FILLER_8_96 ();
 FILLCELL_X1 FILLER_8_98 ();
 FILLCELL_X4 FILLER_8_130 ();
 FILLCELL_X2 FILLER_8_134 ();
 FILLCELL_X1 FILLER_8_136 ();
 FILLCELL_X16 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_201 ();
 FILLCELL_X2 FILLER_8_205 ();
 FILLCELL_X4 FILLER_8_213 ();
 FILLCELL_X2 FILLER_8_217 ();
 FILLCELL_X1 FILLER_8_219 ();
 FILLCELL_X4 FILLER_8_229 ();
 FILLCELL_X1 FILLER_8_233 ();
 FILLCELL_X32 FILLER_8_260 ();
 FILLCELL_X2 FILLER_8_292 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_17 ();
 FILLCELL_X2 FILLER_9_21 ();
 FILLCELL_X8 FILLER_9_37 ();
 FILLCELL_X1 FILLER_9_45 ();
 FILLCELL_X8 FILLER_9_67 ();
 FILLCELL_X4 FILLER_9_75 ();
 FILLCELL_X2 FILLER_9_79 ();
 FILLCELL_X1 FILLER_9_81 ();
 FILLCELL_X2 FILLER_9_89 ();
 FILLCELL_X1 FILLER_9_91 ();
 FILLCELL_X4 FILLER_9_131 ();
 FILLCELL_X2 FILLER_9_149 ();
 FILLCELL_X4 FILLER_9_158 ();
 FILLCELL_X4 FILLER_9_179 ();
 FILLCELL_X2 FILLER_9_190 ();
 FILLCELL_X1 FILLER_9_192 ();
 FILLCELL_X8 FILLER_9_200 ();
 FILLCELL_X1 FILLER_9_208 ();
 FILLCELL_X8 FILLER_9_235 ();
 FILLCELL_X1 FILLER_9_243 ();
 FILLCELL_X8 FILLER_9_284 ();
 FILLCELL_X2 FILLER_9_292 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_41 ();
 FILLCELL_X2 FILLER_10_79 ();
 FILLCELL_X8 FILLER_10_88 ();
 FILLCELL_X4 FILLER_10_96 ();
 FILLCELL_X2 FILLER_10_100 ();
 FILLCELL_X8 FILLER_10_119 ();
 FILLCELL_X4 FILLER_10_127 ();
 FILLCELL_X2 FILLER_10_131 ();
 FILLCELL_X1 FILLER_10_133 ();
 FILLCELL_X16 FILLER_10_182 ();
 FILLCELL_X8 FILLER_10_198 ();
 FILLCELL_X1 FILLER_10_206 ();
 FILLCELL_X8 FILLER_10_225 ();
 FILLCELL_X2 FILLER_10_269 ();
 FILLCELL_X1 FILLER_10_271 ();
 FILLCELL_X2 FILLER_10_292 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_9 ();
 FILLCELL_X4 FILLER_11_35 ();
 FILLCELL_X8 FILLER_11_43 ();
 FILLCELL_X4 FILLER_11_51 ();
 FILLCELL_X1 FILLER_11_55 ();
 FILLCELL_X4 FILLER_11_80 ();
 FILLCELL_X1 FILLER_11_84 ();
 FILLCELL_X16 FILLER_11_116 ();
 FILLCELL_X8 FILLER_11_132 ();
 FILLCELL_X8 FILLER_11_165 ();
 FILLCELL_X1 FILLER_11_173 ();
 FILLCELL_X1 FILLER_11_186 ();
 FILLCELL_X8 FILLER_11_193 ();
 FILLCELL_X4 FILLER_11_201 ();
 FILLCELL_X2 FILLER_11_205 ();
 FILLCELL_X1 FILLER_11_207 ();
 FILLCELL_X8 FILLER_11_213 ();
 FILLCELL_X8 FILLER_11_227 ();
 FILLCELL_X1 FILLER_11_235 ();
 FILLCELL_X4 FILLER_11_245 ();
 FILLCELL_X1 FILLER_11_249 ();
 FILLCELL_X16 FILLER_11_264 ();
 FILLCELL_X8 FILLER_11_280 ();
 FILLCELL_X4 FILLER_11_288 ();
 FILLCELL_X2 FILLER_11_292 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_17 ();
 FILLCELL_X1 FILLER_12_21 ();
 FILLCELL_X32 FILLER_12_29 ();
 FILLCELL_X8 FILLER_12_61 ();
 FILLCELL_X32 FILLER_12_83 ();
 FILLCELL_X16 FILLER_12_115 ();
 FILLCELL_X4 FILLER_12_131 ();
 FILLCELL_X1 FILLER_12_135 ();
 FILLCELL_X1 FILLER_12_153 ();
 FILLCELL_X16 FILLER_12_168 ();
 FILLCELL_X4 FILLER_12_184 ();
 FILLCELL_X1 FILLER_12_194 ();
 FILLCELL_X1 FILLER_12_208 ();
 FILLCELL_X1 FILLER_12_216 ();
 FILLCELL_X1 FILLER_12_230 ();
 FILLCELL_X1 FILLER_12_236 ();
 FILLCELL_X4 FILLER_12_242 ();
 FILLCELL_X2 FILLER_12_246 ();
 FILLCELL_X1 FILLER_12_248 ();
 FILLCELL_X8 FILLER_12_279 ();
 FILLCELL_X4 FILLER_12_287 ();
 FILLCELL_X2 FILLER_12_291 ();
 FILLCELL_X1 FILLER_12_293 ();
 FILLCELL_X4 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_5 ();
 FILLCELL_X1 FILLER_13_7 ();
 FILLCELL_X4 FILLER_13_25 ();
 FILLCELL_X8 FILLER_13_36 ();
 FILLCELL_X4 FILLER_13_44 ();
 FILLCELL_X32 FILLER_13_72 ();
 FILLCELL_X8 FILLER_13_104 ();
 FILLCELL_X4 FILLER_13_112 ();
 FILLCELL_X2 FILLER_13_116 ();
 FILLCELL_X2 FILLER_13_149 ();
 FILLCELL_X4 FILLER_13_168 ();
 FILLCELL_X1 FILLER_13_172 ();
 FILLCELL_X1 FILLER_13_183 ();
 FILLCELL_X4 FILLER_13_213 ();
 FILLCELL_X1 FILLER_13_223 ();
 FILLCELL_X4 FILLER_13_231 ();
 FILLCELL_X2 FILLER_13_235 ();
 FILLCELL_X1 FILLER_13_237 ();
 FILLCELL_X4 FILLER_13_248 ();
 FILLCELL_X1 FILLER_13_252 ();
 FILLCELL_X2 FILLER_13_262 ();
 FILLCELL_X1 FILLER_13_264 ();
 FILLCELL_X1 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_19 ();
 FILLCELL_X2 FILLER_14_28 ();
 FILLCELL_X2 FILLER_14_47 ();
 FILLCELL_X4 FILLER_14_73 ();
 FILLCELL_X2 FILLER_14_84 ();
 FILLCELL_X1 FILLER_14_86 ();
 FILLCELL_X2 FILLER_14_111 ();
 FILLCELL_X1 FILLER_14_113 ();
 FILLCELL_X32 FILLER_14_138 ();
 FILLCELL_X2 FILLER_14_170 ();
 FILLCELL_X8 FILLER_14_177 ();
 FILLCELL_X4 FILLER_14_185 ();
 FILLCELL_X4 FILLER_14_195 ();
 FILLCELL_X8 FILLER_14_212 ();
 FILLCELL_X1 FILLER_14_220 ();
 FILLCELL_X2 FILLER_14_246 ();
 FILLCELL_X1 FILLER_14_271 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_29 ();
 FILLCELL_X16 FILLER_15_38 ();
 FILLCELL_X4 FILLER_15_54 ();
 FILLCELL_X2 FILLER_15_58 ();
 FILLCELL_X1 FILLER_15_60 ();
 FILLCELL_X4 FILLER_15_68 ();
 FILLCELL_X1 FILLER_15_72 ();
 FILLCELL_X32 FILLER_15_104 ();
 FILLCELL_X8 FILLER_15_136 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X16 FILLER_15_169 ();
 FILLCELL_X4 FILLER_15_185 ();
 FILLCELL_X2 FILLER_15_189 ();
 FILLCELL_X16 FILLER_15_222 ();
 FILLCELL_X2 FILLER_15_238 ();
 FILLCELL_X8 FILLER_15_260 ();
 FILLCELL_X4 FILLER_15_268 ();
 FILLCELL_X2 FILLER_15_292 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X2 FILLER_16_21 ();
 FILLCELL_X32 FILLER_16_30 ();
 FILLCELL_X8 FILLER_16_69 ();
 FILLCELL_X4 FILLER_16_84 ();
 FILLCELL_X1 FILLER_16_88 ();
 FILLCELL_X8 FILLER_16_113 ();
 FILLCELL_X4 FILLER_16_121 ();
 FILLCELL_X2 FILLER_16_125 ();
 FILLCELL_X2 FILLER_16_134 ();
 FILLCELL_X2 FILLER_16_143 ();
 FILLCELL_X1 FILLER_16_145 ();
 FILLCELL_X1 FILLER_16_150 ();
 FILLCELL_X2 FILLER_16_158 ();
 FILLCELL_X1 FILLER_16_160 ();
 FILLCELL_X2 FILLER_16_168 ();
 FILLCELL_X1 FILLER_16_170 ();
 FILLCELL_X16 FILLER_16_178 ();
 FILLCELL_X2 FILLER_16_194 ();
 FILLCELL_X1 FILLER_16_198 ();
 FILLCELL_X4 FILLER_16_209 ();
 FILLCELL_X1 FILLER_16_213 ();
 FILLCELL_X2 FILLER_16_236 ();
 FILLCELL_X1 FILLER_16_238 ();
 FILLCELL_X4 FILLER_16_259 ();
 FILLCELL_X2 FILLER_16_263 ();
 FILLCELL_X2 FILLER_16_292 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_9 ();
 FILLCELL_X1 FILLER_17_11 ();
 FILLCELL_X1 FILLER_17_29 ();
 FILLCELL_X8 FILLER_17_44 ();
 FILLCELL_X2 FILLER_17_56 ();
 FILLCELL_X4 FILLER_17_82 ();
 FILLCELL_X2 FILLER_17_86 ();
 FILLCELL_X8 FILLER_17_112 ();
 FILLCELL_X2 FILLER_17_120 ();
 FILLCELL_X1 FILLER_17_122 ();
 FILLCELL_X4 FILLER_17_147 ();
 FILLCELL_X8 FILLER_17_182 ();
 FILLCELL_X2 FILLER_17_190 ();
 FILLCELL_X16 FILLER_17_210 ();
 FILLCELL_X8 FILLER_17_226 ();
 FILLCELL_X16 FILLER_17_276 ();
 FILLCELL_X2 FILLER_17_292 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_5 ();
 FILLCELL_X1 FILLER_18_7 ();
 FILLCELL_X4 FILLER_18_42 ();
 FILLCELL_X1 FILLER_18_46 ();
 FILLCELL_X4 FILLER_18_51 ();
 FILLCELL_X1 FILLER_18_55 ();
 FILLCELL_X8 FILLER_18_87 ();
 FILLCELL_X2 FILLER_18_95 ();
 FILLCELL_X1 FILLER_18_97 ();
 FILLCELL_X16 FILLER_18_112 ();
 FILLCELL_X1 FILLER_18_128 ();
 FILLCELL_X16 FILLER_18_153 ();
 FILLCELL_X2 FILLER_18_169 ();
 FILLCELL_X1 FILLER_18_171 ();
 FILLCELL_X2 FILLER_18_179 ();
 FILLCELL_X1 FILLER_18_199 ();
 FILLCELL_X2 FILLER_18_205 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X1 FILLER_18_257 ();
 FILLCELL_X8 FILLER_18_286 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_9 ();
 FILLCELL_X1 FILLER_19_11 ();
 FILLCELL_X32 FILLER_19_36 ();
 FILLCELL_X16 FILLER_19_68 ();
 FILLCELL_X8 FILLER_19_84 ();
 FILLCELL_X32 FILLER_19_123 ();
 FILLCELL_X8 FILLER_19_155 ();
 FILLCELL_X4 FILLER_19_163 ();
 FILLCELL_X8 FILLER_19_174 ();
 FILLCELL_X4 FILLER_19_182 ();
 FILLCELL_X2 FILLER_19_186 ();
 FILLCELL_X2 FILLER_19_190 ();
 FILLCELL_X8 FILLER_19_214 ();
 FILLCELL_X2 FILLER_19_262 ();
 FILLCELL_X1 FILLER_19_264 ();
 FILLCELL_X8 FILLER_19_286 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_17 ();
 FILLCELL_X2 FILLER_20_21 ();
 FILLCELL_X16 FILLER_20_40 ();
 FILLCELL_X4 FILLER_20_56 ();
 FILLCELL_X4 FILLER_20_77 ();
 FILLCELL_X8 FILLER_20_105 ();
 FILLCELL_X4 FILLER_20_113 ();
 FILLCELL_X2 FILLER_20_117 ();
 FILLCELL_X32 FILLER_20_126 ();
 FILLCELL_X4 FILLER_20_158 ();
 FILLCELL_X2 FILLER_20_162 ();
 FILLCELL_X1 FILLER_20_164 ();
 FILLCELL_X4 FILLER_20_178 ();
 FILLCELL_X1 FILLER_20_182 ();
 FILLCELL_X4 FILLER_20_197 ();
 FILLCELL_X1 FILLER_20_201 ();
 FILLCELL_X4 FILLER_20_207 ();
 FILLCELL_X2 FILLER_20_211 ();
 FILLCELL_X1 FILLER_20_213 ();
 FILLCELL_X32 FILLER_20_234 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_9 ();
 FILLCELL_X1 FILLER_21_13 ();
 FILLCELL_X16 FILLER_21_38 ();
 FILLCELL_X4 FILLER_21_54 ();
 FILLCELL_X4 FILLER_21_89 ();
 FILLCELL_X2 FILLER_21_93 ();
 FILLCELL_X4 FILLER_21_112 ();
 FILLCELL_X8 FILLER_21_140 ();
 FILLCELL_X16 FILLER_21_155 ();
 FILLCELL_X4 FILLER_21_171 ();
 FILLCELL_X2 FILLER_21_175 ();
 FILLCELL_X1 FILLER_21_177 ();
 FILLCELL_X16 FILLER_21_185 ();
 FILLCELL_X2 FILLER_21_201 ();
 FILLCELL_X16 FILLER_21_210 ();
 FILLCELL_X8 FILLER_21_226 ();
 FILLCELL_X2 FILLER_21_234 ();
 FILLCELL_X1 FILLER_21_236 ();
 FILLCELL_X2 FILLER_21_282 ();
 FILLCELL_X1 FILLER_21_293 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X2 FILLER_22_5 ();
 FILLCELL_X8 FILLER_22_31 ();
 FILLCELL_X4 FILLER_22_39 ();
 FILLCELL_X1 FILLER_22_43 ();
 FILLCELL_X16 FILLER_22_68 ();
 FILLCELL_X8 FILLER_22_84 ();
 FILLCELL_X4 FILLER_22_92 ();
 FILLCELL_X1 FILLER_22_96 ();
 FILLCELL_X32 FILLER_22_111 ();
 FILLCELL_X32 FILLER_22_194 ();
 FILLCELL_X16 FILLER_22_226 ();
 FILLCELL_X4 FILLER_22_242 ();
 FILLCELL_X2 FILLER_22_292 ();
 FILLCELL_X8 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_9 ();
 FILLCELL_X8 FILLER_23_35 ();
 FILLCELL_X2 FILLER_23_43 ();
 FILLCELL_X1 FILLER_23_45 ();
 FILLCELL_X16 FILLER_23_94 ();
 FILLCELL_X8 FILLER_23_110 ();
 FILLCELL_X4 FILLER_23_118 ();
 FILLCELL_X2 FILLER_23_146 ();
 FILLCELL_X32 FILLER_23_220 ();
 FILLCELL_X4 FILLER_23_252 ();
 FILLCELL_X1 FILLER_23_256 ();
 FILLCELL_X4 FILLER_23_290 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X8 FILLER_24_17 ();
 FILLCELL_X1 FILLER_24_25 ();
 FILLCELL_X8 FILLER_24_33 ();
 FILLCELL_X4 FILLER_24_41 ();
 FILLCELL_X1 FILLER_24_45 ();
 FILLCELL_X4 FILLER_24_53 ();
 FILLCELL_X2 FILLER_24_57 ();
 FILLCELL_X1 FILLER_24_59 ();
 FILLCELL_X4 FILLER_24_80 ();
 FILLCELL_X2 FILLER_24_84 ();
 FILLCELL_X1 FILLER_24_86 ();
 FILLCELL_X16 FILLER_24_94 ();
 FILLCELL_X4 FILLER_24_110 ();
 FILLCELL_X8 FILLER_24_138 ();
 FILLCELL_X2 FILLER_24_146 ();
 FILLCELL_X2 FILLER_24_155 ();
 FILLCELL_X2 FILLER_24_164 ();
 FILLCELL_X1 FILLER_24_166 ();
 FILLCELL_X4 FILLER_24_181 ();
 FILLCELL_X1 FILLER_24_185 ();
 FILLCELL_X1 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_201 ();
 FILLCELL_X16 FILLER_24_233 ();
 FILLCELL_X8 FILLER_24_249 ();
 FILLCELL_X4 FILLER_24_257 ();
 FILLCELL_X1 FILLER_24_261 ();
 FILLCELL_X2 FILLER_24_291 ();
 FILLCELL_X1 FILLER_24_293 ();
 FILLCELL_X2 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_3 ();
 FILLCELL_X8 FILLER_25_45 ();
 FILLCELL_X1 FILLER_25_53 ();
 FILLCELL_X1 FILLER_25_71 ();
 FILLCELL_X1 FILLER_25_89 ();
 FILLCELL_X1 FILLER_25_104 ();
 FILLCELL_X2 FILLER_25_112 ();
 FILLCELL_X1 FILLER_25_114 ();
 FILLCELL_X2 FILLER_25_117 ();
 FILLCELL_X1 FILLER_25_119 ();
 FILLCELL_X16 FILLER_25_131 ();
 FILLCELL_X8 FILLER_25_147 ();
 FILLCELL_X4 FILLER_25_155 ();
 FILLCELL_X2 FILLER_25_159 ();
 FILLCELL_X1 FILLER_25_161 ();
 FILLCELL_X8 FILLER_25_166 ();
 FILLCELL_X4 FILLER_25_174 ();
 FILLCELL_X2 FILLER_25_182 ();
 FILLCELL_X4 FILLER_25_187 ();
 FILLCELL_X1 FILLER_25_191 ();
 FILLCELL_X1 FILLER_25_204 ();
 FILLCELL_X1 FILLER_25_222 ();
 FILLCELL_X1 FILLER_25_229 ();
 FILLCELL_X2 FILLER_25_254 ();
 FILLCELL_X1 FILLER_25_256 ();
 FILLCELL_X2 FILLER_25_292 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X8 FILLER_26_17 ();
 FILLCELL_X4 FILLER_26_25 ();
 FILLCELL_X2 FILLER_26_29 ();
 FILLCELL_X1 FILLER_26_48 ();
 FILLCELL_X4 FILLER_26_56 ();
 FILLCELL_X2 FILLER_26_60 ();
 FILLCELL_X4 FILLER_26_69 ();
 FILLCELL_X8 FILLER_26_80 ();
 FILLCELL_X2 FILLER_26_88 ();
 FILLCELL_X1 FILLER_26_90 ();
 FILLCELL_X1 FILLER_26_127 ();
 FILLCELL_X16 FILLER_26_132 ();
 FILLCELL_X8 FILLER_26_162 ();
 FILLCELL_X1 FILLER_26_170 ();
 FILLCELL_X1 FILLER_26_202 ();
 FILLCELL_X1 FILLER_26_225 ();
 FILLCELL_X2 FILLER_26_259 ();
 FILLCELL_X1 FILLER_26_261 ();
 FILLCELL_X2 FILLER_26_280 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_33 ();
 FILLCELL_X8 FILLER_27_52 ();
 FILLCELL_X2 FILLER_27_60 ();
 FILLCELL_X8 FILLER_27_79 ();
 FILLCELL_X4 FILLER_27_87 ();
 FILLCELL_X1 FILLER_27_91 ();
 FILLCELL_X4 FILLER_27_123 ();
 FILLCELL_X2 FILLER_27_127 ();
 FILLCELL_X1 FILLER_27_133 ();
 FILLCELL_X2 FILLER_27_151 ();
 FILLCELL_X1 FILLER_27_160 ();
 FILLCELL_X1 FILLER_27_164 ();
 FILLCELL_X1 FILLER_27_182 ();
 FILLCELL_X1 FILLER_27_186 ();
 FILLCELL_X2 FILLER_27_198 ();
 FILLCELL_X1 FILLER_27_200 ();
 FILLCELL_X1 FILLER_27_208 ();
 FILLCELL_X2 FILLER_27_216 ();
 FILLCELL_X4 FILLER_27_245 ();
 FILLCELL_X2 FILLER_27_249 ();
 FILLCELL_X8 FILLER_27_261 ();
 FILLCELL_X16 FILLER_27_275 ();
 FILLCELL_X2 FILLER_27_291 ();
 FILLCELL_X1 FILLER_27_293 ();
 FILLCELL_X8 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_9 ();
 FILLCELL_X1 FILLER_28_13 ();
 FILLCELL_X32 FILLER_28_52 ();
 FILLCELL_X1 FILLER_28_84 ();
 FILLCELL_X8 FILLER_28_113 ();
 FILLCELL_X4 FILLER_28_121 ();
 FILLCELL_X1 FILLER_28_125 ();
 FILLCELL_X4 FILLER_28_137 ();
 FILLCELL_X1 FILLER_28_141 ();
 FILLCELL_X2 FILLER_28_159 ();
 FILLCELL_X1 FILLER_28_165 ();
 FILLCELL_X2 FILLER_28_173 ();
 FILLCELL_X1 FILLER_28_182 ();
 FILLCELL_X1 FILLER_28_192 ();
 FILLCELL_X1 FILLER_28_205 ();
 FILLCELL_X2 FILLER_28_213 ();
 FILLCELL_X1 FILLER_28_215 ();
 FILLCELL_X4 FILLER_28_223 ();
 FILLCELL_X2 FILLER_28_227 ();
 FILLCELL_X1 FILLER_28_229 ();
 FILLCELL_X16 FILLER_28_237 ();
 FILLCELL_X2 FILLER_28_253 ();
 FILLCELL_X1 FILLER_28_255 ();
 FILLCELL_X2 FILLER_28_269 ();
 FILLCELL_X1 FILLER_28_271 ();
 FILLCELL_X2 FILLER_28_292 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X2 FILLER_29_9 ();
 FILLCELL_X1 FILLER_29_11 ();
 FILLCELL_X4 FILLER_29_36 ();
 FILLCELL_X2 FILLER_29_40 ();
 FILLCELL_X4 FILLER_29_49 ();
 FILLCELL_X2 FILLER_29_53 ();
 FILLCELL_X1 FILLER_29_55 ();
 FILLCELL_X2 FILLER_29_80 ();
 FILLCELL_X1 FILLER_29_82 ();
 FILLCELL_X4 FILLER_29_90 ();
 FILLCELL_X2 FILLER_29_94 ();
 FILLCELL_X1 FILLER_29_96 ();
 FILLCELL_X1 FILLER_29_100 ();
 FILLCELL_X8 FILLER_29_107 ();
 FILLCELL_X4 FILLER_29_115 ();
 FILLCELL_X2 FILLER_29_119 ();
 FILLCELL_X1 FILLER_29_121 ();
 FILLCELL_X16 FILLER_29_133 ();
 FILLCELL_X8 FILLER_29_149 ();
 FILLCELL_X4 FILLER_29_168 ();
 FILLCELL_X1 FILLER_29_172 ();
 FILLCELL_X4 FILLER_29_184 ();
 FILLCELL_X1 FILLER_29_188 ();
 FILLCELL_X16 FILLER_29_209 ();
 FILLCELL_X8 FILLER_29_225 ();
 FILLCELL_X2 FILLER_29_237 ();
 FILLCELL_X1 FILLER_29_239 ();
 FILLCELL_X4 FILLER_29_247 ();
 FILLCELL_X4 FILLER_29_265 ();
 FILLCELL_X4 FILLER_29_289 ();
 FILLCELL_X1 FILLER_29_293 ();
 FILLCELL_X16 FILLER_30_1 ();
 FILLCELL_X8 FILLER_30_17 ();
 FILLCELL_X2 FILLER_30_25 ();
 FILLCELL_X8 FILLER_30_51 ();
 FILLCELL_X4 FILLER_30_59 ();
 FILLCELL_X2 FILLER_30_63 ();
 FILLCELL_X4 FILLER_30_72 ();
 FILLCELL_X4 FILLER_30_83 ();
 FILLCELL_X1 FILLER_30_87 ();
 FILLCELL_X4 FILLER_30_95 ();
 FILLCELL_X1 FILLER_30_99 ();
 FILLCELL_X1 FILLER_30_107 ();
 FILLCELL_X8 FILLER_30_111 ();
 FILLCELL_X4 FILLER_30_119 ();
 FILLCELL_X2 FILLER_30_123 ();
 FILLCELL_X8 FILLER_30_129 ();
 FILLCELL_X4 FILLER_30_137 ();
 FILLCELL_X1 FILLER_30_141 ();
 FILLCELL_X8 FILLER_30_144 ();
 FILLCELL_X4 FILLER_30_152 ();
 FILLCELL_X2 FILLER_30_156 ();
 FILLCELL_X1 FILLER_30_158 ();
 FILLCELL_X8 FILLER_30_176 ();
 FILLCELL_X4 FILLER_30_184 ();
 FILLCELL_X1 FILLER_30_188 ();
 FILLCELL_X16 FILLER_30_202 ();
 FILLCELL_X8 FILLER_30_218 ();
 FILLCELL_X4 FILLER_30_226 ();
 FILLCELL_X1 FILLER_30_230 ();
 FILLCELL_X2 FILLER_30_238 ();
 FILLCELL_X1 FILLER_30_240 ();
 FILLCELL_X1 FILLER_30_250 ();
 FILLCELL_X16 FILLER_30_269 ();
 FILLCELL_X8 FILLER_30_285 ();
 FILLCELL_X1 FILLER_30_293 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X8 FILLER_31_33 ();
 FILLCELL_X4 FILLER_31_41 ();
 FILLCELL_X1 FILLER_31_45 ();
 FILLCELL_X8 FILLER_31_53 ();
 FILLCELL_X2 FILLER_31_61 ();
 FILLCELL_X1 FILLER_31_63 ();
 FILLCELL_X4 FILLER_31_81 ();
 FILLCELL_X2 FILLER_31_85 ();
 FILLCELL_X8 FILLER_31_104 ();
 FILLCELL_X2 FILLER_31_112 ();
 FILLCELL_X1 FILLER_31_114 ();
 FILLCELL_X1 FILLER_31_139 ();
 FILLCELL_X2 FILLER_31_147 ();
 FILLCELL_X1 FILLER_31_166 ();
 FILLCELL_X8 FILLER_31_174 ();
 FILLCELL_X4 FILLER_31_182 ();
 FILLCELL_X8 FILLER_31_213 ();
 FILLCELL_X4 FILLER_31_221 ();
 FILLCELL_X2 FILLER_31_225 ();
 FILLCELL_X8 FILLER_31_256 ();
 FILLCELL_X4 FILLER_31_264 ();
 FILLCELL_X1 FILLER_31_268 ();
 FILLCELL_X16 FILLER_31_276 ();
 FILLCELL_X2 FILLER_31_292 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_33 ();
 FILLCELL_X1 FILLER_32_58 ();
 FILLCELL_X8 FILLER_32_66 ();
 FILLCELL_X4 FILLER_32_74 ();
 FILLCELL_X1 FILLER_32_78 ();
 FILLCELL_X1 FILLER_32_96 ();
 FILLCELL_X2 FILLER_32_100 ();
 FILLCELL_X8 FILLER_32_108 ();
 FILLCELL_X2 FILLER_32_116 ();
 FILLCELL_X1 FILLER_32_118 ();
 FILLCELL_X8 FILLER_32_143 ();
 FILLCELL_X4 FILLER_32_151 ();
 FILLCELL_X2 FILLER_32_155 ();
 FILLCELL_X2 FILLER_32_174 ();
 FILLCELL_X2 FILLER_32_182 ();
 FILLCELL_X1 FILLER_32_184 ();
 FILLCELL_X8 FILLER_32_196 ();
 FILLCELL_X2 FILLER_32_204 ();
 FILLCELL_X1 FILLER_32_206 ();
 FILLCELL_X32 FILLER_32_209 ();
 FILLCELL_X4 FILLER_32_241 ();
 FILLCELL_X2 FILLER_32_245 ();
 FILLCELL_X1 FILLER_32_250 ();
 FILLCELL_X1 FILLER_32_257 ();
 FILLCELL_X1 FILLER_32_271 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X4 FILLER_33_33 ();
 FILLCELL_X2 FILLER_33_37 ();
 FILLCELL_X16 FILLER_33_56 ();
 FILLCELL_X4 FILLER_33_72 ();
 FILLCELL_X2 FILLER_33_76 ();
 FILLCELL_X1 FILLER_33_78 ();
 FILLCELL_X4 FILLER_33_86 ();
 FILLCELL_X2 FILLER_33_90 ();
 FILLCELL_X4 FILLER_33_99 ();
 FILLCELL_X16 FILLER_33_110 ();
 FILLCELL_X2 FILLER_33_126 ();
 FILLCELL_X16 FILLER_33_139 ();
 FILLCELL_X8 FILLER_33_155 ();
 FILLCELL_X2 FILLER_33_163 ();
 FILLCELL_X2 FILLER_33_182 ();
 FILLCELL_X1 FILLER_33_184 ();
 FILLCELL_X32 FILLER_33_209 ();
 FILLCELL_X2 FILLER_33_241 ();
 FILLCELL_X1 FILLER_33_243 ();
 FILLCELL_X2 FILLER_33_292 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X4 FILLER_34_33 ();
 FILLCELL_X2 FILLER_34_37 ();
 FILLCELL_X16 FILLER_34_60 ();
 FILLCELL_X4 FILLER_34_76 ();
 FILLCELL_X1 FILLER_34_80 ();
 FILLCELL_X2 FILLER_34_107 ();
 FILLCELL_X1 FILLER_34_109 ();
 FILLCELL_X4 FILLER_34_113 ();
 FILLCELL_X1 FILLER_34_117 ();
 FILLCELL_X8 FILLER_34_151 ();
 FILLCELL_X2 FILLER_34_173 ();
 FILLCELL_X8 FILLER_34_182 ();
 FILLCELL_X1 FILLER_34_190 ();
 FILLCELL_X32 FILLER_34_231 ();
 FILLCELL_X16 FILLER_34_263 ();
 FILLCELL_X8 FILLER_34_279 ();
 FILLCELL_X4 FILLER_34_287 ();
 FILLCELL_X2 FILLER_34_291 ();
 FILLCELL_X1 FILLER_34_293 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X4 FILLER_35_33 ();
 FILLCELL_X4 FILLER_35_71 ();
 FILLCELL_X2 FILLER_35_75 ();
 FILLCELL_X1 FILLER_35_77 ();
 FILLCELL_X4 FILLER_35_102 ();
 FILLCELL_X2 FILLER_35_106 ();
 FILLCELL_X4 FILLER_35_112 ();
 FILLCELL_X4 FILLER_35_133 ();
 FILLCELL_X1 FILLER_35_137 ();
 FILLCELL_X8 FILLER_35_142 ();
 FILLCELL_X2 FILLER_35_150 ();
 FILLCELL_X8 FILLER_35_169 ();
 FILLCELL_X2 FILLER_35_177 ();
 FILLCELL_X1 FILLER_35_227 ();
 FILLCELL_X32 FILLER_35_245 ();
 FILLCELL_X16 FILLER_35_277 ();
 FILLCELL_X1 FILLER_35_293 ();
 FILLCELL_X4 FILLER_36_1 ();
 FILLCELL_X8 FILLER_36_30 ();
 FILLCELL_X2 FILLER_36_38 ();
 FILLCELL_X1 FILLER_36_40 ();
 FILLCELL_X2 FILLER_36_58 ();
 FILLCELL_X4 FILLER_36_67 ();
 FILLCELL_X2 FILLER_36_71 ();
 FILLCELL_X1 FILLER_36_80 ();
 FILLCELL_X2 FILLER_36_98 ();
 FILLCELL_X1 FILLER_36_100 ();
 FILLCELL_X2 FILLER_36_120 ();
 FILLCELL_X2 FILLER_36_126 ();
 FILLCELL_X1 FILLER_36_128 ();
 FILLCELL_X2 FILLER_36_133 ();
 FILLCELL_X1 FILLER_36_135 ();
 FILLCELL_X2 FILLER_36_155 ();
 FILLCELL_X4 FILLER_36_163 ();
 FILLCELL_X2 FILLER_36_167 ();
 FILLCELL_X8 FILLER_36_173 ();
 FILLCELL_X2 FILLER_36_181 ();
 FILLCELL_X2 FILLER_36_187 ();
 FILLCELL_X1 FILLER_36_189 ();
 FILLCELL_X2 FILLER_36_214 ();
 FILLCELL_X2 FILLER_36_223 ();
 FILLCELL_X1 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_233 ();
 FILLCELL_X16 FILLER_36_265 ();
 FILLCELL_X8 FILLER_36_281 ();
 FILLCELL_X4 FILLER_36_289 ();
 FILLCELL_X1 FILLER_36_293 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X8 FILLER_37_33 ();
 FILLCELL_X4 FILLER_37_41 ();
 FILLCELL_X1 FILLER_37_45 ();
 FILLCELL_X8 FILLER_37_70 ();
 FILLCELL_X4 FILLER_37_78 ();
 FILLCELL_X1 FILLER_37_82 ();
 FILLCELL_X8 FILLER_37_97 ();
 FILLCELL_X1 FILLER_37_124 ();
 FILLCELL_X2 FILLER_37_142 ();
 FILLCELL_X2 FILLER_37_161 ();
 FILLCELL_X4 FILLER_37_197 ();
 FILLCELL_X2 FILLER_37_201 ();
 FILLCELL_X1 FILLER_37_203 ();
 FILLCELL_X8 FILLER_37_211 ();
 FILLCELL_X4 FILLER_37_219 ();
 FILLCELL_X2 FILLER_37_223 ();
 FILLCELL_X32 FILLER_37_249 ();
 FILLCELL_X8 FILLER_37_281 ();
 FILLCELL_X4 FILLER_37_289 ();
 FILLCELL_X1 FILLER_37_293 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X2 FILLER_38_97 ();
 FILLCELL_X4 FILLER_38_102 ();
 FILLCELL_X2 FILLER_38_106 ();
 FILLCELL_X16 FILLER_38_111 ();
 FILLCELL_X2 FILLER_38_127 ();
 FILLCELL_X1 FILLER_38_129 ();
 FILLCELL_X1 FILLER_38_132 ();
 FILLCELL_X2 FILLER_38_136 ();
 FILLCELL_X4 FILLER_38_141 ();
 FILLCELL_X2 FILLER_38_145 ();
 FILLCELL_X1 FILLER_38_147 ();
 FILLCELL_X4 FILLER_38_154 ();
 FILLCELL_X2 FILLER_38_158 ();
 FILLCELL_X4 FILLER_38_163 ();
 FILLCELL_X1 FILLER_38_167 ();
 FILLCELL_X8 FILLER_38_170 ();
 FILLCELL_X4 FILLER_38_178 ();
 FILLCELL_X32 FILLER_38_184 ();
 FILLCELL_X32 FILLER_38_216 ();
 FILLCELL_X32 FILLER_38_248 ();
 FILLCELL_X8 FILLER_38_280 ();
 FILLCELL_X4 FILLER_38_288 ();
 FILLCELL_X2 FILLER_38_292 ();
endmodule
