module configurable_carry_select_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [63:0] a;
 input [63:0] b;
 output [63:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire \first_block.full_adders[0].fa.sum ;
 wire \first_block.full_adders[1].fa.sum ;
 wire \first_block.full_adders[2].fa.sum ;
 wire \first_block.full_adders[3].fa.sum ;
 wire \first_block.full_adders[4].fa.sum ;
 wire \first_block.full_adders[5].fa.sum ;
 wire \first_block.full_adders[6].fa.sum ;
 wire \first_block.full_adders[7].fa.sum ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;

 INV_X1 _465_ (.A(net1),
    .ZN(_306_));
 INV_X1 _466_ (.A(net65),
    .ZN(_307_));
 INV_X1 _467_ (.A(net129),
    .ZN(_308_));
 INV_X1 _468_ (.A(_309_),
    .ZN(_310_));
 INV_X1 _469_ (.A(_312_),
    .ZN(\first_block.full_adders[1].fa.sum ));
 INV_X1 _470_ (.A(_314_),
    .ZN(\first_block.full_adders[2].fa.sum ));
 INV_X1 _471_ (.A(_316_),
    .ZN(\first_block.full_adders[3].fa.sum ));
 INV_X1 _472_ (.A(_318_),
    .ZN(\first_block.full_adders[4].fa.sum ));
 INV_X1 _473_ (.A(_320_),
    .ZN(\first_block.full_adders[5].fa.sum ));
 INV_X1 _474_ (.A(_322_),
    .ZN(\first_block.full_adders[6].fa.sum ));
 INV_X1 _475_ (.A(_324_),
    .ZN(\first_block.full_adders[7].fa.sum ));
 INV_X1 _476_ (.A(net43),
    .ZN(_325_));
 INV_X1 _477_ (.A(net52),
    .ZN(_331_));
 INV_X1 _478_ (.A(net8),
    .ZN(_337_));
 INV_X1 _479_ (.A(net17),
    .ZN(_343_));
 INV_X1 _480_ (.A(net26),
    .ZN(_349_));
 INV_X1 _481_ (.A(net35),
    .ZN(_355_));
 INV_X1 _482_ (.A(net63),
    .ZN(_459_));
 INV_X1 _483_ (.A(net107),
    .ZN(_326_));
 INV_X1 _484_ (.A(net116),
    .ZN(_332_));
 INV_X1 _485_ (.A(net72),
    .ZN(_338_));
 INV_X1 _486_ (.A(net81),
    .ZN(_344_));
 INV_X1 _487_ (.A(net90),
    .ZN(_350_));
 INV_X1 _488_ (.A(net99),
    .ZN(_356_));
 INV_X1 _489_ (.A(net127),
    .ZN(_460_));
 OR2_X1 _490_ (.A1(_447_),
    .A2(_449_),
    .ZN(_000_));
 OAI33_X1 _491_ (.A1(net59),
    .A2(net123),
    .A3(_447_),
    .B1(_000_),
    .B2(net58),
    .B3(net122),
    .ZN(_001_));
 INV_X1 _492_ (.A(_453_),
    .ZN(_002_));
 NOR2_X1 _493_ (.A1(net55),
    .A2(net119),
    .ZN(_003_));
 OR2_X1 _494_ (.A1(net54),
    .A2(net118),
    .ZN(_004_));
 INV_X1 _495_ (.A(_457_),
    .ZN(_005_));
 NOR2_X1 _496_ (.A1(net53),
    .A2(net117),
    .ZN(_006_));
 INV_X1 _497_ (.A(_335_),
    .ZN(_007_));
 OAI21_X1 _498_ (.A(_005_),
    .B1(_006_),
    .B2(_007_),
    .ZN(_008_));
 AOI21_X1 _499_ (.A(_455_),
    .B1(_004_),
    .B2(_008_),
    .ZN(_009_));
 OAI21_X1 _500_ (.A(_002_),
    .B1(_003_),
    .B2(_009_),
    .ZN(_010_));
 OAI21_X1 _501_ (.A(_010_),
    .B1(net121),
    .B2(net57),
    .ZN(_011_));
 OAI21_X1 _502_ (.A(_005_),
    .B1(_006_),
    .B2(_333_),
    .ZN(_012_));
 AOI21_X1 _503_ (.A(_455_),
    .B1(_004_),
    .B2(_012_),
    .ZN(_013_));
 OAI21_X1 _504_ (.A(_002_),
    .B1(_003_),
    .B2(_013_),
    .ZN(_014_));
 OAI21_X1 _505_ (.A(_014_),
    .B1(net121),
    .B2(net57),
    .ZN(_015_));
 NOR3_X1 _506_ (.A1(net51),
    .A2(net115),
    .A3(_431_),
    .ZN(_016_));
 INV_X1 _507_ (.A(_433_),
    .ZN(_017_));
 NOR2_X1 _508_ (.A1(net50),
    .A2(net114),
    .ZN(_018_));
 NOR2_X1 _509_ (.A1(net49),
    .A2(net113),
    .ZN(_019_));
 OR2_X1 _510_ (.A1(net48),
    .A2(net112),
    .ZN(_020_));
 INV_X1 _511_ (.A(_439_),
    .ZN(_021_));
 OR2_X1 _512_ (.A1(net47),
    .A2(net111),
    .ZN(_022_));
 NOR2_X1 _513_ (.A1(net46),
    .A2(net110),
    .ZN(_023_));
 OAI21_X1 _514_ (.A(_329_),
    .B1(net108),
    .B2(net44),
    .ZN(_024_));
 INV_X1 _515_ (.A(_443_),
    .ZN(_025_));
 AOI21_X1 _516_ (.A(_023_),
    .B1(_024_),
    .B2(_025_),
    .ZN(_026_));
 OAI21_X1 _517_ (.A(_022_),
    .B1(_026_),
    .B2(_441_),
    .ZN(_027_));
 NAND2_X1 _518_ (.A1(_021_),
    .A2(_027_),
    .ZN(_028_));
 AOI21_X1 _519_ (.A(_437_),
    .B1(_020_),
    .B2(_028_),
    .ZN(_029_));
 NOR2_X1 _520_ (.A1(_019_),
    .A2(_029_),
    .ZN(_030_));
 NOR2_X1 _521_ (.A1(_435_),
    .A2(_030_),
    .ZN(_031_));
 OAI21_X1 _522_ (.A(_017_),
    .B1(_018_),
    .B2(_031_),
    .ZN(_032_));
 NOR3_X1 _523_ (.A1(_417_),
    .A2(_431_),
    .A3(_032_),
    .ZN(_033_));
 OR2_X2 _524_ (.A1(net42),
    .A2(net106),
    .ZN(_034_));
 OR2_X2 _525_ (.A1(net41),
    .A2(net105),
    .ZN(_035_));
 AOI21_X4 _526_ (.A(_419_),
    .B1(_421_),
    .B2(_035_),
    .ZN(_036_));
 OAI21_X4 _527_ (.A(_035_),
    .B1(net104),
    .B2(net40),
    .ZN(_037_));
 NOR2_X1 _528_ (.A1(net39),
    .A2(net103),
    .ZN(_038_));
 OR2_X1 _529_ (.A1(net38),
    .A2(net102),
    .ZN(_039_));
 NOR2_X1 _530_ (.A1(net37),
    .A2(net101),
    .ZN(_040_));
 OAI21_X1 _531_ (.A(_359_),
    .B1(net100),
    .B2(net36),
    .ZN(_041_));
 INV_X1 _532_ (.A(_429_),
    .ZN(_042_));
 AOI21_X1 _533_ (.A(_040_),
    .B1(_041_),
    .B2(_042_),
    .ZN(_043_));
 OAI21_X1 _534_ (.A(_039_),
    .B1(_043_),
    .B2(_427_),
    .ZN(_044_));
 INV_X1 _535_ (.A(_425_),
    .ZN(_045_));
 AOI21_X1 _536_ (.A(_038_),
    .B1(_044_),
    .B2(_045_),
    .ZN(_046_));
 NOR2_X2 _537_ (.A1(_423_),
    .A2(_046_),
    .ZN(_047_));
 OAI21_X4 _538_ (.A(_036_),
    .B1(_037_),
    .B2(_047_),
    .ZN(_048_));
 NAND2_X1 _539_ (.A1(_034_),
    .A2(_048_),
    .ZN(_049_));
 NOR4_X2 _540_ (.A1(net22),
    .A2(net86),
    .A3(_391_),
    .A4(_393_),
    .ZN(_050_));
 NOR2_X1 _541_ (.A1(net24),
    .A2(net88),
    .ZN(_051_));
 INV_X1 _542_ (.A(_391_),
    .ZN(_052_));
 INV_X1 _543_ (.A(net25),
    .ZN(_053_));
 INV_X1 _544_ (.A(net89),
    .ZN(_054_));
 AOI221_X2 _545_ (.A(_050_),
    .B1(_051_),
    .B2(_052_),
    .C1(_053_),
    .C2(_054_),
    .ZN(_055_));
 OAI22_X2 _546_ (.A1(net20),
    .A2(net84),
    .B1(net21),
    .B2(net85),
    .ZN(_056_));
 NOR2_X1 _547_ (.A1(net19),
    .A2(net83),
    .ZN(_057_));
 INV_X1 _548_ (.A(_399_),
    .ZN(_058_));
 NOR2_X1 _549_ (.A1(_399_),
    .A2(_401_),
    .ZN(_059_));
 OAI21_X1 _550_ (.A(_347_),
    .B1(net82),
    .B2(net18),
    .ZN(_060_));
 AOI221_X2 _551_ (.A(_056_),
    .B1(_057_),
    .B2(_058_),
    .C1(_059_),
    .C2(_060_),
    .ZN(_061_));
 INV_X2 _552_ (.A(_395_),
    .ZN(_062_));
 NOR3_X2 _553_ (.A1(_389_),
    .A2(_391_),
    .A3(_393_),
    .ZN(_063_));
 OAI21_X4 _554_ (.A(_397_),
    .B1(net85),
    .B2(net21),
    .ZN(_064_));
 NAND3_X2 _555_ (.A1(_062_),
    .A2(_063_),
    .A3(_064_),
    .ZN(_065_));
 OAI22_X4 _556_ (.A1(_389_),
    .A2(_055_),
    .B1(_061_),
    .B2(_065_),
    .ZN(_066_));
 OR2_X1 _557_ (.A1(net20),
    .A2(net84),
    .ZN(_067_));
 OAI22_X4 _558_ (.A1(net21),
    .A2(net85),
    .B1(_397_),
    .B2(_067_),
    .ZN(_068_));
 OR3_X1 _559_ (.A1(net18),
    .A2(net82),
    .A3(_401_),
    .ZN(_069_));
 INV_X1 _560_ (.A(_345_),
    .ZN(_070_));
 OAI221_X2 _561_ (.A(_069_),
    .B1(_401_),
    .B2(_070_),
    .C1(net19),
    .C2(net83),
    .ZN(_071_));
 NOR3_X2 _562_ (.A1(_395_),
    .A2(_397_),
    .A3(_399_),
    .ZN(_072_));
 AOI22_X4 _563_ (.A1(_062_),
    .A2(_068_),
    .B1(_071_),
    .B2(_072_),
    .ZN(_073_));
 NOR4_X4 _564_ (.A1(_389_),
    .A2(_391_),
    .A3(_393_),
    .A4(_073_),
    .ZN(_074_));
 NOR2_X1 _565_ (.A1(_066_),
    .A2(_074_),
    .ZN(_075_));
 OR2_X2 _566_ (.A1(_361_),
    .A2(_363_),
    .ZN(_076_));
 NOR2_X2 _567_ (.A1(net6),
    .A2(net70),
    .ZN(_077_));
 OAI21_X2 _568_ (.A(_367_),
    .B1(net69),
    .B2(net5),
    .ZN(_078_));
 INV_X1 _569_ (.A(_365_),
    .ZN(_079_));
 AOI21_X4 _570_ (.A(_077_),
    .B1(_078_),
    .B2(_079_),
    .ZN(_080_));
 NOR2_X1 _571_ (.A1(_076_),
    .A2(_080_),
    .ZN(_081_));
 NOR2_X1 _572_ (.A1(net4),
    .A2(net68),
    .ZN(_082_));
 NOR4_X4 _573_ (.A1(net2),
    .A2(net66),
    .A3(_369_),
    .A4(_371_),
    .ZN(_083_));
 OR2_X1 _574_ (.A1(net3),
    .A2(net67),
    .ZN(_084_));
 NOR2_X1 _575_ (.A1(_369_),
    .A2(_084_),
    .ZN(_085_));
 NOR3_X4 _576_ (.A1(_082_),
    .A2(_083_),
    .A3(_085_),
    .ZN(_086_));
 NOR3_X2 _577_ (.A1(_369_),
    .A2(_371_),
    .A3(_373_),
    .ZN(_087_));
 NOR2_X2 _578_ (.A1(net64),
    .A2(net128),
    .ZN(_088_));
 INV_X1 _579_ (.A(_463_),
    .ZN(_089_));
 MUX2_X2 _580_ (.A(_089_),
    .B(_461_),
    .S(_323_),
    .Z(_090_));
 OAI21_X4 _581_ (.A(_087_),
    .B1(_088_),
    .B2(_090_),
    .ZN(_091_));
 NOR2_X2 _582_ (.A1(net5),
    .A2(net69),
    .ZN(_092_));
 NOR2_X4 _583_ (.A1(_077_),
    .A2(_092_),
    .ZN(_093_));
 NAND3_X2 _584_ (.A1(_086_),
    .A2(_091_),
    .A3(_093_),
    .ZN(_094_));
 AOI21_X1 _585_ (.A(_066_),
    .B1(_081_),
    .B2(_094_),
    .ZN(_095_));
 OR3_X4 _586_ (.A1(net7),
    .A2(net71),
    .A3(_361_),
    .ZN(_096_));
 OR2_X1 _587_ (.A1(net16),
    .A2(net80),
    .ZN(_097_));
 AOI21_X2 _588_ (.A(_375_),
    .B1(_377_),
    .B2(_097_),
    .ZN(_098_));
 OAI22_X4 _589_ (.A1(net15),
    .A2(net79),
    .B1(net16),
    .B2(net80),
    .ZN(_099_));
 INV_X1 _590_ (.A(_379_),
    .ZN(_100_));
 OAI21_X4 _591_ (.A(_098_),
    .B1(_099_),
    .B2(_100_),
    .ZN(_101_));
 NOR4_X2 _592_ (.A1(net11),
    .A2(net75),
    .A3(_381_),
    .A4(_383_),
    .ZN(_102_));
 NOR3_X2 _593_ (.A1(net13),
    .A2(net77),
    .A3(_381_),
    .ZN(_103_));
 NOR2_X1 _594_ (.A1(net14),
    .A2(net78),
    .ZN(_104_));
 OR4_X4 _595_ (.A1(_099_),
    .A2(_102_),
    .A3(_103_),
    .A4(_104_),
    .ZN(_105_));
 OAI21_X1 _596_ (.A(_387_),
    .B1(net74),
    .B2(net10),
    .ZN(_106_));
 NOR3_X1 _597_ (.A1(_381_),
    .A2(_383_),
    .A3(_385_),
    .ZN(_107_));
 AND2_X2 _598_ (.A1(_106_),
    .A2(_107_),
    .ZN(_108_));
 NOR2_X1 _599_ (.A1(net10),
    .A2(net74),
    .ZN(_109_));
 NOR2_X1 _600_ (.A1(net9),
    .A2(net73),
    .ZN(_110_));
 OR3_X2 _601_ (.A1(_339_),
    .A2(_109_),
    .A3(_110_),
    .ZN(_111_));
 AOI21_X4 _602_ (.A(_105_),
    .B1(_108_),
    .B2(_111_),
    .ZN(_112_));
 NOR2_X2 _603_ (.A1(_101_),
    .A2(_112_),
    .ZN(_113_));
 AND2_X1 _604_ (.A1(_096_),
    .A2(_113_),
    .ZN(_114_));
 OAI221_X2 _605_ (.A(_341_),
    .B1(net74),
    .B2(net10),
    .C1(net9),
    .C2(net73),
    .ZN(_115_));
 AOI21_X4 _606_ (.A(_105_),
    .B1(_108_),
    .B2(_115_),
    .ZN(_116_));
 NOR3_X1 _607_ (.A1(_066_),
    .A2(_101_),
    .A3(_116_),
    .ZN(_117_));
 OR2_X1 _608_ (.A1(_076_),
    .A2(_080_),
    .ZN(_118_));
 AND2_X2 _609_ (.A1(_096_),
    .A2(_118_),
    .ZN(_119_));
 AND4_X2 _610_ (.A1(_096_),
    .A2(_086_),
    .A3(_091_),
    .A4(_093_),
    .ZN(_120_));
 NOR2_X4 _611_ (.A1(_119_),
    .A2(_120_),
    .ZN(_121_));
 AOI221_X4 _612_ (.A(_075_),
    .B1(_095_),
    .B2(_114_),
    .C1(_117_),
    .C2(_121_),
    .ZN(_122_));
 NOR2_X1 _613_ (.A1(_389_),
    .A2(_055_),
    .ZN(_123_));
 NOR2_X2 _614_ (.A1(_123_),
    .A2(_074_),
    .ZN(_124_));
 NOR2_X1 _615_ (.A1(_101_),
    .A2(_116_),
    .ZN(_125_));
 NAND2_X4 _616_ (.A1(_096_),
    .A2(_118_),
    .ZN(_126_));
 NAND4_X4 _617_ (.A1(_096_),
    .A2(_086_),
    .A3(_091_),
    .A4(_093_),
    .ZN(_127_));
 NAND3_X2 _618_ (.A1(_125_),
    .A2(_126_),
    .A3(_127_),
    .ZN(_128_));
 OAI21_X4 _619_ (.A(_113_),
    .B1(_120_),
    .B2(_119_),
    .ZN(_129_));
 NAND3_X4 _620_ (.A1(_124_),
    .A2(_128_),
    .A3(_129_),
    .ZN(_130_));
 INV_X1 _621_ (.A(_403_),
    .ZN(_131_));
 NOR2_X1 _622_ (.A1(net32),
    .A2(net96),
    .ZN(_132_));
 OR2_X1 _623_ (.A1(net31),
    .A2(net95),
    .ZN(_133_));
 AOI21_X1 _624_ (.A(_407_),
    .B1(_409_),
    .B2(_133_),
    .ZN(_134_));
 NOR2_X1 _625_ (.A1(_132_),
    .A2(_134_),
    .ZN(_135_));
 NOR2_X2 _626_ (.A1(_405_),
    .A2(_135_),
    .ZN(_136_));
 NOR2_X2 _627_ (.A1(net33),
    .A2(net97),
    .ZN(_137_));
 OAI21_X4 _628_ (.A(_131_),
    .B1(_136_),
    .B2(_137_),
    .ZN(_138_));
 OAI221_X2 _629_ (.A(_133_),
    .B1(net96),
    .B2(net32),
    .C1(net30),
    .C2(net94),
    .ZN(_139_));
 NOR2_X4 _630_ (.A1(_137_),
    .A2(_139_),
    .ZN(_140_));
 INV_X2 _631_ (.A(_411_),
    .ZN(_141_));
 NOR2_X2 _632_ (.A1(net29),
    .A2(net93),
    .ZN(_142_));
 INV_X1 _633_ (.A(_142_),
    .ZN(_143_));
 INV_X1 _634_ (.A(_413_),
    .ZN(_144_));
 NOR2_X1 _635_ (.A1(net28),
    .A2(net92),
    .ZN(_145_));
 OR2_X1 _636_ (.A1(net27),
    .A2(net91),
    .ZN(_146_));
 AOI21_X1 _637_ (.A(_415_),
    .B1(_146_),
    .B2(_353_),
    .ZN(_147_));
 OAI21_X1 _638_ (.A(_144_),
    .B1(_145_),
    .B2(_147_),
    .ZN(_148_));
 NAND2_X1 _639_ (.A1(_143_),
    .A2(_148_),
    .ZN(_149_));
 NAND2_X2 _640_ (.A1(_141_),
    .A2(_149_),
    .ZN(_150_));
 AOI21_X2 _641_ (.A(_138_),
    .B1(_140_),
    .B2(_150_),
    .ZN(_151_));
 NAND3_X4 _642_ (.A1(_122_),
    .A2(_130_),
    .A3(_151_),
    .ZN(_152_));
 OR2_X1 _643_ (.A1(net28),
    .A2(net92),
    .ZN(_153_));
 INV_X1 _644_ (.A(_415_),
    .ZN(_154_));
 NOR2_X1 _645_ (.A1(net27),
    .A2(net91),
    .ZN(_155_));
 OAI21_X1 _646_ (.A(_154_),
    .B1(_155_),
    .B2(_351_),
    .ZN(_156_));
 AOI21_X1 _647_ (.A(_413_),
    .B1(_153_),
    .B2(_156_),
    .ZN(_157_));
 OAI21_X2 _648_ (.A(_141_),
    .B1(_142_),
    .B2(_157_),
    .ZN(_158_));
 AOI21_X2 _649_ (.A(_138_),
    .B1(_140_),
    .B2(_158_),
    .ZN(_159_));
 INV_X1 _650_ (.A(_064_),
    .ZN(_160_));
 NOR3_X2 _651_ (.A1(_395_),
    .A2(_061_),
    .A3(_160_),
    .ZN(_161_));
 AOI21_X1 _652_ (.A(_123_),
    .B1(_063_),
    .B2(_161_),
    .ZN(_162_));
 NAND4_X1 _653_ (.A1(_162_),
    .A2(_125_),
    .A3(_126_),
    .A4(_127_),
    .ZN(_163_));
 AND2_X1 _654_ (.A1(_081_),
    .A2(_094_),
    .ZN(_164_));
 NAND3_X1 _655_ (.A1(_162_),
    .A2(_096_),
    .A3(_113_),
    .ZN(_165_));
 OAI221_X2 _656_ (.A(_163_),
    .B1(_164_),
    .B2(_165_),
    .C1(_074_),
    .C2(_066_),
    .ZN(_166_));
 AND3_X2 _657_ (.A1(_124_),
    .A2(_128_),
    .A3(_129_),
    .ZN(_167_));
 OAI21_X4 _658_ (.A(_159_),
    .B1(_166_),
    .B2(_167_),
    .ZN(_168_));
 AOI21_X4 _659_ (.A(_049_),
    .B1(_152_),
    .B2(_168_),
    .ZN(_169_));
 INV_X1 _660_ (.A(_038_),
    .ZN(_170_));
 NOR2_X1 _661_ (.A1(net38),
    .A2(net102),
    .ZN(_171_));
 INV_X1 _662_ (.A(_040_),
    .ZN(_172_));
 NOR2_X1 _663_ (.A1(net36),
    .A2(net100),
    .ZN(_173_));
 OAI21_X1 _664_ (.A(_042_),
    .B1(_173_),
    .B2(_357_),
    .ZN(_174_));
 AOI21_X1 _665_ (.A(_427_),
    .B1(_172_),
    .B2(_174_),
    .ZN(_175_));
 OAI21_X1 _666_ (.A(_045_),
    .B1(_171_),
    .B2(_175_),
    .ZN(_176_));
 AOI21_X2 _667_ (.A(_423_),
    .B1(_170_),
    .B2(_176_),
    .ZN(_177_));
 OAI21_X4 _668_ (.A(_036_),
    .B1(_037_),
    .B2(_177_),
    .ZN(_178_));
 AND4_X2 _669_ (.A1(_034_),
    .A2(_168_),
    .A3(_152_),
    .A4(_178_),
    .ZN(_179_));
 NOR2_X4 _670_ (.A1(_169_),
    .A2(_179_),
    .ZN(_180_));
 INV_X1 _671_ (.A(_018_),
    .ZN(_181_));
 INV_X1 _672_ (.A(_437_),
    .ZN(_182_));
 INV_X1 _673_ (.A(_441_),
    .ZN(_183_));
 OR2_X1 _674_ (.A1(net44),
    .A2(net108),
    .ZN(_184_));
 INV_X1 _675_ (.A(_327_),
    .ZN(_185_));
 AOI21_X1 _676_ (.A(_443_),
    .B1(_184_),
    .B2(_185_),
    .ZN(_186_));
 OAI21_X1 _677_ (.A(_183_),
    .B1(_023_),
    .B2(_186_),
    .ZN(_187_));
 AOI21_X1 _678_ (.A(_439_),
    .B1(_022_),
    .B2(_187_),
    .ZN(_188_));
 NOR2_X1 _679_ (.A1(net48),
    .A2(net112),
    .ZN(_189_));
 OAI21_X1 _680_ (.A(_182_),
    .B1(_188_),
    .B2(_189_),
    .ZN(_190_));
 NOR2_X1 _681_ (.A1(_018_),
    .A2(_019_),
    .ZN(_191_));
 AOI221_X2 _682_ (.A(_433_),
    .B1(_435_),
    .B2(_181_),
    .C1(_190_),
    .C2(_191_),
    .ZN(_192_));
 AND3_X1 _683_ (.A1(_192_),
    .A2(_034_),
    .A3(_048_),
    .ZN(_193_));
 AND3_X1 _684_ (.A1(_122_),
    .A2(_130_),
    .A3(_151_),
    .ZN(_194_));
 AOI221_X2 _685_ (.A(_138_),
    .B1(_140_),
    .B2(_158_),
    .C1(_122_),
    .C2(_130_),
    .ZN(_195_));
 OAI21_X2 _686_ (.A(_193_),
    .B1(_194_),
    .B2(_195_),
    .ZN(_196_));
 AND3_X1 _687_ (.A1(_192_),
    .A2(_034_),
    .A3(_178_),
    .ZN(_197_));
 NAND3_X2 _688_ (.A1(_168_),
    .A2(_152_),
    .A3(_197_),
    .ZN(_198_));
 NAND2_X1 _689_ (.A1(_417_),
    .A2(_192_),
    .ZN(_199_));
 NAND3_X4 _690_ (.A1(_196_),
    .A2(_198_),
    .A3(_199_),
    .ZN(_200_));
 INV_X1 _691_ (.A(_431_),
    .ZN(_201_));
 AOI221_X2 _692_ (.A(_016_),
    .B1(_033_),
    .B2(_180_),
    .C1(_200_),
    .C2(_201_),
    .ZN(_202_));
 MUX2_X1 _693_ (.A(_011_),
    .B(_015_),
    .S(_202_),
    .Z(_203_));
 NOR2_X1 _694_ (.A1(_451_),
    .A2(_000_),
    .ZN(_204_));
 INV_X1 _695_ (.A(net124),
    .ZN(_205_));
 INV_X1 _696_ (.A(net60),
    .ZN(_206_));
 AOI221_X1 _697_ (.A(_001_),
    .B1(_203_),
    .B2(_204_),
    .C1(_205_),
    .C2(_206_),
    .ZN(_207_));
 OR2_X1 _698_ (.A1(_445_),
    .A2(_207_),
    .ZN(net130));
 NOR2_X1 _699_ (.A1(_090_),
    .A2(_088_),
    .ZN(_208_));
 NOR2_X1 _700_ (.A1(_373_),
    .A2(_208_),
    .ZN(_209_));
 XNOR2_X1 _701_ (.A(_372_),
    .B(_209_),
    .ZN(net132));
 INV_X1 _702_ (.A(_371_),
    .ZN(_210_));
 NOR2_X1 _703_ (.A1(net2),
    .A2(net66),
    .ZN(_211_));
 OAI21_X1 _704_ (.A(_210_),
    .B1(_211_),
    .B2(_209_),
    .ZN(_212_));
 XOR2_X1 _705_ (.A(_370_),
    .B(_212_),
    .Z(net133));
 AOI21_X1 _706_ (.A(_369_),
    .B1(_084_),
    .B2(_212_),
    .ZN(_213_));
 XNOR2_X1 _707_ (.A(_368_),
    .B(_213_),
    .ZN(net134));
 AOI21_X1 _708_ (.A(_367_),
    .B1(_086_),
    .B2(_091_),
    .ZN(_214_));
 XNOR2_X1 _709_ (.A(_366_),
    .B(_214_),
    .ZN(net135));
 AND2_X1 _710_ (.A1(_079_),
    .A2(_078_),
    .ZN(_215_));
 NAND2_X1 _711_ (.A1(_086_),
    .A2(_091_),
    .ZN(_216_));
 OAI21_X1 _712_ (.A(_215_),
    .B1(_216_),
    .B2(_092_),
    .ZN(_217_));
 XOR2_X1 _713_ (.A(_364_),
    .B(_217_),
    .Z(net136));
 OR2_X1 _714_ (.A1(net6),
    .A2(net70),
    .ZN(_218_));
 AOI21_X1 _715_ (.A(_363_),
    .B1(_218_),
    .B2(_217_),
    .ZN(_219_));
 XNOR2_X1 _716_ (.A(_362_),
    .B(_219_),
    .ZN(net137));
 XNOR2_X1 _717_ (.A(_340_),
    .B(_121_),
    .ZN(net138));
 AOI21_X1 _718_ (.A(_339_),
    .B1(_126_),
    .B2(_127_),
    .ZN(_220_));
 AOI21_X2 _719_ (.A(_220_),
    .B1(_121_),
    .B2(_341_),
    .ZN(_221_));
 XNOR2_X1 _720_ (.A(_388_),
    .B(_221_),
    .ZN(net139));
 NOR2_X1 _721_ (.A1(_110_),
    .A2(_221_),
    .ZN(_222_));
 NOR2_X1 _722_ (.A1(_387_),
    .A2(_222_),
    .ZN(_223_));
 XNOR2_X1 _723_ (.A(_386_),
    .B(_223_),
    .ZN(net140));
 INV_X1 _724_ (.A(_385_),
    .ZN(_224_));
 OAI21_X2 _725_ (.A(_224_),
    .B1(_109_),
    .B2(_223_),
    .ZN(_225_));
 XOR2_X1 _726_ (.A(_384_),
    .B(_225_),
    .Z(net141));
 OR2_X1 _727_ (.A1(net11),
    .A2(net75),
    .ZN(_226_));
 AOI21_X1 _728_ (.A(_383_),
    .B1(_226_),
    .B2(_225_),
    .ZN(_227_));
 XNOR2_X1 _729_ (.A(_382_),
    .B(_227_),
    .ZN(net143));
 NOR2_X1 _730_ (.A1(_102_),
    .A2(_103_),
    .ZN(_228_));
 OR2_X1 _731_ (.A1(_381_),
    .A2(_383_),
    .ZN(_229_));
 OAI21_X1 _732_ (.A(_228_),
    .B1(_225_),
    .B2(_229_),
    .ZN(_230_));
 XNOR2_X1 _733_ (.A(_380_),
    .B(_230_),
    .ZN(net144));
 OAI21_X1 _734_ (.A(_100_),
    .B1(_104_),
    .B2(_230_),
    .ZN(_231_));
 XOR2_X1 _735_ (.A(_378_),
    .B(_231_),
    .Z(net145));
 OR2_X1 _736_ (.A1(net15),
    .A2(net79),
    .ZN(_232_));
 AOI21_X1 _737_ (.A(_377_),
    .B1(_232_),
    .B2(_231_),
    .ZN(_233_));
 XNOR2_X1 _738_ (.A(_376_),
    .B(_233_),
    .ZN(net146));
 AND2_X4 _739_ (.A1(_128_),
    .A2(_129_),
    .ZN(_234_));
 XOR2_X1 _740_ (.A(_346_),
    .B(_234_),
    .Z(net147));
 INV_X1 _741_ (.A(_347_),
    .ZN(_235_));
 MUX2_X1 _742_ (.A(_235_),
    .B(_345_),
    .S(_234_),
    .Z(_236_));
 XNOR2_X1 _743_ (.A(_402_),
    .B(_236_),
    .ZN(net148));
 NOR2_X1 _744_ (.A1(net18),
    .A2(net82),
    .ZN(_237_));
 NOR2_X1 _745_ (.A1(_237_),
    .A2(_236_),
    .ZN(_238_));
 NOR2_X1 _746_ (.A1(_401_),
    .A2(_238_),
    .ZN(_239_));
 XNOR2_X1 _747_ (.A(_400_),
    .B(_239_),
    .ZN(net149));
 OAI21_X1 _748_ (.A(_058_),
    .B1(_057_),
    .B2(_239_),
    .ZN(_240_));
 XOR2_X1 _749_ (.A(_398_),
    .B(_240_),
    .Z(net150));
 AOI21_X1 _750_ (.A(_397_),
    .B1(_067_),
    .B2(_240_),
    .ZN(_241_));
 XNOR2_X1 _751_ (.A(_396_),
    .B(_241_),
    .ZN(net151));
 NAND2_X1 _752_ (.A1(_073_),
    .A2(_234_),
    .ZN(_242_));
 OAI21_X4 _753_ (.A(_242_),
    .B1(_234_),
    .B2(_161_),
    .ZN(_243_));
 XOR2_X1 _754_ (.A(_394_),
    .B(_243_),
    .Z(net152));
 OR2_X1 _755_ (.A1(net22),
    .A2(net86),
    .ZN(_244_));
 AOI21_X2 _756_ (.A(_393_),
    .B1(_244_),
    .B2(_243_),
    .ZN(_245_));
 XNOR2_X1 _757_ (.A(_392_),
    .B(_245_),
    .ZN(net154));
 OAI21_X1 _758_ (.A(_052_),
    .B1(_051_),
    .B2(_245_),
    .ZN(_246_));
 XOR2_X1 _759_ (.A(_390_),
    .B(_246_),
    .Z(net155));
 NAND2_X2 _760_ (.A1(_122_),
    .A2(_130_),
    .ZN(_247_));
 XOR2_X2 _761_ (.A(_352_),
    .B(_247_),
    .Z(net156));
 OAI21_X2 _762_ (.A(_351_),
    .B1(_166_),
    .B2(_167_),
    .ZN(_248_));
 OAI21_X4 _763_ (.A(_248_),
    .B1(_247_),
    .B2(_353_),
    .ZN(_249_));
 XNOR2_X2 _764_ (.A(_416_),
    .B(_249_),
    .ZN(net157));
 NOR3_X1 _765_ (.A1(_353_),
    .A2(_166_),
    .A3(_167_),
    .ZN(_250_));
 AOI21_X2 _766_ (.A(_250_),
    .B1(_247_),
    .B2(_351_),
    .ZN(_251_));
 AOI21_X2 _767_ (.A(_415_),
    .B1(_146_),
    .B2(_251_),
    .ZN(_252_));
 XNOR2_X2 _768_ (.A(_414_),
    .B(_252_),
    .ZN(net158));
 OAI21_X2 _769_ (.A(_154_),
    .B1(_155_),
    .B2(_249_),
    .ZN(_253_));
 AOI21_X4 _770_ (.A(_413_),
    .B1(_153_),
    .B2(_253_),
    .ZN(_254_));
 XNOR2_X2 _771_ (.A(_412_),
    .B(_254_),
    .ZN(net159));
 OAI21_X2 _772_ (.A(_144_),
    .B1(_145_),
    .B2(_252_),
    .ZN(_255_));
 AOI21_X4 _773_ (.A(_411_),
    .B1(_143_),
    .B2(_255_),
    .ZN(_256_));
 XNOR2_X1 _774_ (.A(_410_),
    .B(_256_),
    .ZN(net160));
 INV_X1 _775_ (.A(_409_),
    .ZN(_257_));
 NOR2_X1 _776_ (.A1(net30),
    .A2(net94),
    .ZN(_258_));
 OAI21_X2 _777_ (.A(_257_),
    .B1(_258_),
    .B2(_256_),
    .ZN(_259_));
 XOR2_X1 _778_ (.A(_408_),
    .B(_259_),
    .Z(net161));
 OR2_X1 _779_ (.A1(_406_),
    .A2(_407_),
    .ZN(_260_));
 OAI21_X4 _780_ (.A(_141_),
    .B1(_142_),
    .B2(_254_),
    .ZN(_261_));
 INV_X1 _781_ (.A(_258_),
    .ZN(_262_));
 AOI211_X2 _782_ (.A(_409_),
    .B(_260_),
    .C1(_261_),
    .C2(_262_),
    .ZN(_263_));
 NAND2_X1 _783_ (.A1(_406_),
    .A2(_407_),
    .ZN(_264_));
 OAI21_X1 _784_ (.A(_264_),
    .B1(_260_),
    .B2(_133_),
    .ZN(_265_));
 AND2_X1 _785_ (.A1(_406_),
    .A2(_133_),
    .ZN(_266_));
 AOI211_X2 _786_ (.A(_263_),
    .B(_265_),
    .C1(_259_),
    .C2(_266_),
    .ZN(net162));
 OAI21_X1 _787_ (.A(_136_),
    .B1(_139_),
    .B2(_256_),
    .ZN(_267_));
 XOR2_X1 _788_ (.A(_404_),
    .B(_267_),
    .Z(net163));
 NAND2_X4 _789_ (.A1(_168_),
    .A2(_152_),
    .ZN(_268_));
 XNOR2_X1 _790_ (.A(_358_),
    .B(_268_),
    .ZN(net165));
 OAI21_X4 _791_ (.A(_359_),
    .B1(_195_),
    .B2(_194_),
    .ZN(_269_));
 OAI21_X2 _792_ (.A(_269_),
    .B1(_268_),
    .B2(_357_),
    .ZN(_270_));
 XOR2_X1 _793_ (.A(_430_),
    .B(_270_),
    .Z(net166));
 OR2_X1 _794_ (.A1(net36),
    .A2(net100),
    .ZN(_271_));
 AOI21_X2 _795_ (.A(_429_),
    .B1(_271_),
    .B2(_270_),
    .ZN(_272_));
 XNOR2_X1 _796_ (.A(_428_),
    .B(_272_),
    .ZN(net167));
 INV_X1 _797_ (.A(_427_),
    .ZN(_273_));
 OAI21_X1 _798_ (.A(_273_),
    .B1(_040_),
    .B2(_272_),
    .ZN(_274_));
 XOR2_X1 _799_ (.A(_426_),
    .B(_274_),
    .Z(net168));
 AOI21_X1 _800_ (.A(_425_),
    .B1(_039_),
    .B2(_274_),
    .ZN(_275_));
 XNOR2_X1 _801_ (.A(_424_),
    .B(_275_),
    .ZN(net169));
 MUX2_X1 _802_ (.A(_177_),
    .B(_047_),
    .S(_268_),
    .Z(_276_));
 XNOR2_X1 _803_ (.A(_422_),
    .B(_276_),
    .ZN(net170));
 INV_X1 _804_ (.A(_421_),
    .ZN(_277_));
 NOR2_X1 _805_ (.A1(net40),
    .A2(net104),
    .ZN(_278_));
 OAI21_X1 _806_ (.A(_277_),
    .B1(_278_),
    .B2(_276_),
    .ZN(_279_));
 XOR2_X1 _807_ (.A(_420_),
    .B(_279_),
    .Z(net171));
 MUX2_X1 _808_ (.A(_178_),
    .B(_048_),
    .S(_268_),
    .Z(_280_));
 XOR2_X1 _809_ (.A(_418_),
    .B(_280_),
    .Z(net172));
 NOR3_X4 _810_ (.A1(_417_),
    .A2(_169_),
    .A3(_179_),
    .ZN(_281_));
 XNOR2_X2 _811_ (.A(_328_),
    .B(_281_),
    .ZN(net173));
 MUX2_X1 _812_ (.A(_185_),
    .B(_329_),
    .S(_281_),
    .Z(_282_));
 XOR2_X2 _813_ (.A(_444_),
    .B(_282_),
    .Z(net174));
 AOI21_X2 _814_ (.A(_443_),
    .B1(_184_),
    .B2(_282_),
    .ZN(_283_));
 XNOR2_X1 _815_ (.A(_442_),
    .B(_283_),
    .ZN(net176));
 OAI21_X1 _816_ (.A(_183_),
    .B1(_023_),
    .B2(_283_),
    .ZN(_284_));
 XOR2_X1 _817_ (.A(_440_),
    .B(_284_),
    .Z(net177));
 NAND2_X1 _818_ (.A1(_022_),
    .A2(_187_),
    .ZN(_285_));
 NAND2_X1 _819_ (.A1(_021_),
    .A2(_285_),
    .ZN(_286_));
 MUX2_X1 _820_ (.A(_286_),
    .B(_028_),
    .S(_281_),
    .Z(_287_));
 XOR2_X1 _821_ (.A(_438_),
    .B(_287_),
    .Z(net178));
 AOI21_X1 _822_ (.A(_437_),
    .B1(_286_),
    .B2(_020_),
    .ZN(_288_));
 MUX2_X1 _823_ (.A(_288_),
    .B(_029_),
    .S(_281_),
    .Z(_289_));
 XNOR2_X1 _824_ (.A(_436_),
    .B(_289_),
    .ZN(net179));
 NAND2_X1 _825_ (.A1(_281_),
    .A2(_031_),
    .ZN(_290_));
 INV_X1 _826_ (.A(_435_),
    .ZN(_291_));
 OAI21_X1 _827_ (.A(_291_),
    .B1(_288_),
    .B2(_019_),
    .ZN(_292_));
 OAI21_X1 _828_ (.A(_290_),
    .B1(_281_),
    .B2(_292_),
    .ZN(_293_));
 XNOR2_X1 _829_ (.A(_434_),
    .B(_293_),
    .ZN(net180));
 INV_X1 _830_ (.A(_032_),
    .ZN(_294_));
 AOI21_X1 _831_ (.A(_200_),
    .B1(_294_),
    .B2(_281_),
    .ZN(_295_));
 XOR2_X1 _832_ (.A(_432_),
    .B(_295_),
    .Z(net181));
 XOR2_X1 _833_ (.A(_334_),
    .B(_202_),
    .Z(net182));
 MUX2_X1 _834_ (.A(_007_),
    .B(_333_),
    .S(_202_),
    .Z(_296_));
 XNOR2_X1 _835_ (.A(_458_),
    .B(_296_),
    .ZN(net183));
 MUX2_X1 _836_ (.A(_008_),
    .B(_012_),
    .S(_202_),
    .Z(_297_));
 XOR2_X1 _837_ (.A(_456_),
    .B(_297_),
    .Z(net184));
 AOI21_X1 _838_ (.A(_455_),
    .B1(_004_),
    .B2(_297_),
    .ZN(_298_));
 XNOR2_X1 _839_ (.A(_454_),
    .B(_298_),
    .ZN(net185));
 MUX2_X1 _840_ (.A(_010_),
    .B(_014_),
    .S(_202_),
    .Z(_299_));
 XOR2_X1 _841_ (.A(_452_),
    .B(_299_),
    .Z(net187));
 INV_X1 _842_ (.A(_451_),
    .ZN(_300_));
 NAND2_X1 _843_ (.A1(_300_),
    .A2(_203_),
    .ZN(_301_));
 XOR2_X1 _844_ (.A(_450_),
    .B(_301_),
    .Z(net188));
 NOR3_X1 _845_ (.A1(net58),
    .A2(net122),
    .A3(_449_),
    .ZN(_302_));
 NOR2_X1 _846_ (.A1(_449_),
    .A2(_451_),
    .ZN(_303_));
 AOI21_X1 _847_ (.A(_302_),
    .B1(_203_),
    .B2(_303_),
    .ZN(_304_));
 XOR2_X1 _848_ (.A(_448_),
    .B(_304_),
    .Z(net189));
 AOI21_X1 _849_ (.A(_001_),
    .B1(_203_),
    .B2(_204_),
    .ZN(_305_));
 XOR2_X1 _850_ (.A(_446_),
    .B(_305_),
    .Z(net190));
 XOR2_X1 _851_ (.A(_323_),
    .B(_462_),
    .Z(net193));
 XNOR2_X1 _852_ (.A(_374_),
    .B(_090_),
    .ZN(net194));
 FA_X1 _853_ (.A(_306_),
    .B(_307_),
    .CI(_308_),
    .CO(_309_),
    .S(\first_block.full_adders[0].fa.sum ));
 FA_X1 _854_ (.A(net12),
    .B(net76),
    .CI(_310_),
    .CO(_311_),
    .S(_312_));
 FA_X1 _855_ (.A(net23),
    .B(net87),
    .CI(_311_),
    .CO(_313_),
    .S(_314_));
 FA_X1 _856_ (.A(net34),
    .B(net98),
    .CI(_313_),
    .CO(_315_),
    .S(_316_));
 FA_X1 _857_ (.A(net45),
    .B(net109),
    .CI(_315_),
    .CO(_317_),
    .S(_318_));
 FA_X1 _858_ (.A(net56),
    .B(net120),
    .CI(_317_),
    .CO(_319_),
    .S(_320_));
 FA_X1 _859_ (.A(net61),
    .B(net125),
    .CI(_319_),
    .CO(_321_),
    .S(_322_));
 FA_X1 _860_ (.A(net62),
    .B(net126),
    .CI(_321_),
    .CO(_323_),
    .S(_324_));
 HA_X1 _861_ (.A(_325_),
    .B(_326_),
    .CO(_327_),
    .S(_328_));
 HA_X1 _862_ (.A(net43),
    .B(net107),
    .CO(_329_),
    .S(_330_));
 HA_X1 _863_ (.A(_331_),
    .B(_332_),
    .CO(_333_),
    .S(_334_));
 HA_X1 _864_ (.A(net52),
    .B(net116),
    .CO(_335_),
    .S(_336_));
 HA_X1 _865_ (.A(_337_),
    .B(_338_),
    .CO(_339_),
    .S(_340_));
 HA_X1 _866_ (.A(net8),
    .B(net72),
    .CO(_341_),
    .S(_342_));
 HA_X1 _867_ (.A(_343_),
    .B(_344_),
    .CO(_345_),
    .S(_346_));
 HA_X1 _868_ (.A(net17),
    .B(net81),
    .CO(_347_),
    .S(_348_));
 HA_X1 _869_ (.A(_349_),
    .B(_350_),
    .CO(_351_),
    .S(_352_));
 HA_X1 _870_ (.A(net26),
    .B(net90),
    .CO(_353_),
    .S(_354_));
 HA_X1 _871_ (.A(_355_),
    .B(_356_),
    .CO(_357_),
    .S(_358_));
 HA_X1 _872_ (.A(net35),
    .B(net99),
    .CO(_359_),
    .S(_360_));
 HA_X1 _873_ (.A(net7),
    .B(net71),
    .CO(_361_),
    .S(_362_));
 HA_X1 _874_ (.A(net6),
    .B(net70),
    .CO(_363_),
    .S(_364_));
 HA_X1 _875_ (.A(net5),
    .B(net69),
    .CO(_365_),
    .S(_366_));
 HA_X1 _876_ (.A(net4),
    .B(net68),
    .CO(_367_),
    .S(_368_));
 HA_X1 _877_ (.A(net3),
    .B(net67),
    .CO(_369_),
    .S(_370_));
 HA_X1 _878_ (.A(net2),
    .B(net66),
    .CO(_371_),
    .S(_372_));
 HA_X1 _879_ (.A(net64),
    .B(net128),
    .CO(_373_),
    .S(_374_));
 HA_X1 _880_ (.A(net16),
    .B(net80),
    .CO(_375_),
    .S(_376_));
 HA_X1 _881_ (.A(net15),
    .B(net79),
    .CO(_377_),
    .S(_378_));
 HA_X1 _882_ (.A(net14),
    .B(net78),
    .CO(_379_),
    .S(_380_));
 HA_X1 _883_ (.A(net13),
    .B(net77),
    .CO(_381_),
    .S(_382_));
 HA_X1 _884_ (.A(net11),
    .B(net75),
    .CO(_383_),
    .S(_384_));
 HA_X1 _885_ (.A(net10),
    .B(net74),
    .CO(_385_),
    .S(_386_));
 HA_X1 _886_ (.A(net9),
    .B(net73),
    .CO(_387_),
    .S(_388_));
 HA_X1 _887_ (.A(net25),
    .B(net89),
    .CO(_389_),
    .S(_390_));
 HA_X1 _888_ (.A(net24),
    .B(net88),
    .CO(_391_),
    .S(_392_));
 HA_X1 _889_ (.A(net22),
    .B(net86),
    .CO(_393_),
    .S(_394_));
 HA_X1 _890_ (.A(net21),
    .B(net85),
    .CO(_395_),
    .S(_396_));
 HA_X1 _891_ (.A(net20),
    .B(net84),
    .CO(_397_),
    .S(_398_));
 HA_X1 _892_ (.A(net19),
    .B(net83),
    .CO(_399_),
    .S(_400_));
 HA_X1 _893_ (.A(net18),
    .B(net82),
    .CO(_401_),
    .S(_402_));
 HA_X1 _894_ (.A(net33),
    .B(net97),
    .CO(_403_),
    .S(_404_));
 HA_X1 _895_ (.A(net32),
    .B(net96),
    .CO(_405_),
    .S(_406_));
 HA_X1 _896_ (.A(net31),
    .B(net95),
    .CO(_407_),
    .S(_408_));
 HA_X1 _897_ (.A(net30),
    .B(net94),
    .CO(_409_),
    .S(_410_));
 HA_X1 _898_ (.A(net29),
    .B(net93),
    .CO(_411_),
    .S(_412_));
 HA_X1 _899_ (.A(net28),
    .B(net92),
    .CO(_413_),
    .S(_414_));
 HA_X1 _900_ (.A(net27),
    .B(net91),
    .CO(_415_),
    .S(_416_));
 HA_X1 _901_ (.A(net42),
    .B(net106),
    .CO(_417_),
    .S(_418_));
 HA_X1 _902_ (.A(net41),
    .B(net105),
    .CO(_419_),
    .S(_420_));
 HA_X1 _903_ (.A(net40),
    .B(net104),
    .CO(_421_),
    .S(_422_));
 HA_X1 _904_ (.A(net39),
    .B(net103),
    .CO(_423_),
    .S(_424_));
 HA_X1 _905_ (.A(net38),
    .B(net102),
    .CO(_425_),
    .S(_426_));
 HA_X1 _906_ (.A(net37),
    .B(net101),
    .CO(_427_),
    .S(_428_));
 HA_X1 _907_ (.A(net36),
    .B(net100),
    .CO(_429_),
    .S(_430_));
 HA_X1 _908_ (.A(net51),
    .B(net115),
    .CO(_431_),
    .S(_432_));
 HA_X1 _909_ (.A(net50),
    .B(net114),
    .CO(_433_),
    .S(_434_));
 HA_X1 _910_ (.A(net49),
    .B(net113),
    .CO(_435_),
    .S(_436_));
 HA_X1 _911_ (.A(net48),
    .B(net112),
    .CO(_437_),
    .S(_438_));
 HA_X1 _912_ (.A(net47),
    .B(net111),
    .CO(_439_),
    .S(_440_));
 HA_X1 _913_ (.A(net46),
    .B(net110),
    .CO(_441_),
    .S(_442_));
 HA_X1 _914_ (.A(net44),
    .B(net108),
    .CO(_443_),
    .S(_444_));
 HA_X1 _915_ (.A(net60),
    .B(net124),
    .CO(_445_),
    .S(_446_));
 HA_X1 _916_ (.A(net59),
    .B(net123),
    .CO(_447_),
    .S(_448_));
 HA_X1 _917_ (.A(net58),
    .B(net122),
    .CO(_449_),
    .S(_450_));
 HA_X1 _918_ (.A(net57),
    .B(net121),
    .CO(_451_),
    .S(_452_));
 HA_X1 _919_ (.A(net55),
    .B(net119),
    .CO(_453_),
    .S(_454_));
 HA_X1 _920_ (.A(net54),
    .B(net118),
    .CO(_455_),
    .S(_456_));
 HA_X1 _921_ (.A(net53),
    .B(net117),
    .CO(_457_),
    .S(_458_));
 HA_X1 _922_ (.A(_459_),
    .B(_460_),
    .CO(_461_),
    .S(_462_));
 HA_X1 _923_ (.A(net63),
    .B(net127),
    .CO(_463_),
    .S(_464_));
 BUF_X1 _924_ (.A(\first_block.full_adders[0].fa.sum ),
    .Z(net131));
 BUF_X1 _925_ (.A(\first_block.full_adders[1].fa.sum ),
    .Z(net142));
 BUF_X1 _926_ (.A(\first_block.full_adders[2].fa.sum ),
    .Z(net153));
 BUF_X1 _927_ (.A(\first_block.full_adders[3].fa.sum ),
    .Z(net164));
 BUF_X1 _928_ (.A(\first_block.full_adders[4].fa.sum ),
    .Z(net175));
 BUF_X1 _929_ (.A(\first_block.full_adders[5].fa.sum ),
    .Z(net186));
 BUF_X1 _930_ (.A(\first_block.full_adders[6].fa.sum ),
    .Z(net191));
 BUF_X1 _931_ (.A(\first_block.full_adders[7].fa.sum ),
    .Z(net192));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_730 ();
 BUF_X1 input1 (.A(a[0]),
    .Z(net1));
 CLKBUF_X2 input2 (.A(a[10]),
    .Z(net2));
 BUF_X1 input3 (.A(a[11]),
    .Z(net3));
 BUF_X1 input4 (.A(a[12]),
    .Z(net4));
 CLKBUF_X2 input5 (.A(a[13]),
    .Z(net5));
 BUF_X1 input6 (.A(a[14]),
    .Z(net6));
 BUF_X1 input7 (.A(a[15]),
    .Z(net7));
 BUF_X1 input8 (.A(a[16]),
    .Z(net8));
 BUF_X1 input9 (.A(a[17]),
    .Z(net9));
 CLKBUF_X2 input10 (.A(a[18]),
    .Z(net10));
 BUF_X1 input11 (.A(a[19]),
    .Z(net11));
 BUF_X1 input12 (.A(a[1]),
    .Z(net12));
 BUF_X1 input13 (.A(a[20]),
    .Z(net13));
 BUF_X1 input14 (.A(a[21]),
    .Z(net14));
 CLKBUF_X2 input15 (.A(a[22]),
    .Z(net15));
 CLKBUF_X2 input16 (.A(a[23]),
    .Z(net16));
 BUF_X1 input17 (.A(a[24]),
    .Z(net17));
 BUF_X1 input18 (.A(a[25]),
    .Z(net18));
 BUF_X1 input19 (.A(a[26]),
    .Z(net19));
 BUF_X1 input20 (.A(a[27]),
    .Z(net20));
 CLKBUF_X3 input21 (.A(a[28]),
    .Z(net21));
 BUF_X1 input22 (.A(a[29]),
    .Z(net22));
 BUF_X1 input23 (.A(a[2]),
    .Z(net23));
 BUF_X1 input24 (.A(a[30]),
    .Z(net24));
 BUF_X1 input25 (.A(a[31]),
    .Z(net25));
 CLKBUF_X3 input26 (.A(a[32]),
    .Z(net26));
 BUF_X2 input27 (.A(a[33]),
    .Z(net27));
 BUF_X2 input28 (.A(a[34]),
    .Z(net28));
 BUF_X2 input29 (.A(a[35]),
    .Z(net29));
 BUF_X1 input30 (.A(a[36]),
    .Z(net30));
 BUF_X1 input31 (.A(a[37]),
    .Z(net31));
 BUF_X1 input32 (.A(a[38]),
    .Z(net32));
 BUF_X1 input33 (.A(a[39]),
    .Z(net33));
 BUF_X1 input34 (.A(a[3]),
    .Z(net34));
 BUF_X1 input35 (.A(a[40]),
    .Z(net35));
 BUF_X1 input36 (.A(a[41]),
    .Z(net36));
 BUF_X1 input37 (.A(a[42]),
    .Z(net37));
 BUF_X1 input38 (.A(a[43]),
    .Z(net38));
 BUF_X1 input39 (.A(a[44]),
    .Z(net39));
 CLKBUF_X2 input40 (.A(a[45]),
    .Z(net40));
 BUF_X1 input41 (.A(a[46]),
    .Z(net41));
 BUF_X1 input42 (.A(a[47]),
    .Z(net42));
 BUF_X1 input43 (.A(a[48]),
    .Z(net43));
 BUF_X4 input44 (.A(a[49]),
    .Z(net44));
 BUF_X1 input45 (.A(a[4]),
    .Z(net45));
 BUF_X1 input46 (.A(a[50]),
    .Z(net46));
 BUF_X1 input47 (.A(a[51]),
    .Z(net47));
 BUF_X1 input48 (.A(a[52]),
    .Z(net48));
 BUF_X1 input49 (.A(a[53]),
    .Z(net49));
 BUF_X1 input50 (.A(a[54]),
    .Z(net50));
 BUF_X1 input51 (.A(a[55]),
    .Z(net51));
 BUF_X1 input52 (.A(a[56]),
    .Z(net52));
 BUF_X1 input53 (.A(a[57]),
    .Z(net53));
 BUF_X1 input54 (.A(a[58]),
    .Z(net54));
 BUF_X1 input55 (.A(a[59]),
    .Z(net55));
 BUF_X1 input56 (.A(a[5]),
    .Z(net56));
 BUF_X1 input57 (.A(a[60]),
    .Z(net57));
 BUF_X1 input58 (.A(a[61]),
    .Z(net58));
 BUF_X1 input59 (.A(a[62]),
    .Z(net59));
 BUF_X1 input60 (.A(a[63]),
    .Z(net60));
 BUF_X1 input61 (.A(a[6]),
    .Z(net61));
 BUF_X1 input62 (.A(a[7]),
    .Z(net62));
 BUF_X1 input63 (.A(a[8]),
    .Z(net63));
 BUF_X1 input64 (.A(a[9]),
    .Z(net64));
 BUF_X1 input65 (.A(b[0]),
    .Z(net65));
 CLKBUF_X2 input66 (.A(b[10]),
    .Z(net66));
 BUF_X1 input67 (.A(b[11]),
    .Z(net67));
 BUF_X1 input68 (.A(b[12]),
    .Z(net68));
 CLKBUF_X2 input69 (.A(b[13]),
    .Z(net69));
 BUF_X1 input70 (.A(b[14]),
    .Z(net70));
 BUF_X1 input71 (.A(b[15]),
    .Z(net71));
 BUF_X1 input72 (.A(b[16]),
    .Z(net72));
 BUF_X1 input73 (.A(b[17]),
    .Z(net73));
 CLKBUF_X2 input74 (.A(b[18]),
    .Z(net74));
 BUF_X1 input75 (.A(b[19]),
    .Z(net75));
 BUF_X1 input76 (.A(b[1]),
    .Z(net76));
 BUF_X1 input77 (.A(b[20]),
    .Z(net77));
 BUF_X1 input78 (.A(b[21]),
    .Z(net78));
 CLKBUF_X2 input79 (.A(b[22]),
    .Z(net79));
 CLKBUF_X2 input80 (.A(b[23]),
    .Z(net80));
 BUF_X1 input81 (.A(b[24]),
    .Z(net81));
 BUF_X1 input82 (.A(b[25]),
    .Z(net82));
 BUF_X1 input83 (.A(b[26]),
    .Z(net83));
 BUF_X1 input84 (.A(b[27]),
    .Z(net84));
 CLKBUF_X3 input85 (.A(b[28]),
    .Z(net85));
 BUF_X1 input86 (.A(b[29]),
    .Z(net86));
 BUF_X1 input87 (.A(b[2]),
    .Z(net87));
 BUF_X1 input88 (.A(b[30]),
    .Z(net88));
 BUF_X1 input89 (.A(b[31]),
    .Z(net89));
 CLKBUF_X3 input90 (.A(b[32]),
    .Z(net90));
 BUF_X2 input91 (.A(b[33]),
    .Z(net91));
 BUF_X2 input92 (.A(b[34]),
    .Z(net92));
 BUF_X2 input93 (.A(b[35]),
    .Z(net93));
 BUF_X1 input94 (.A(b[36]),
    .Z(net94));
 BUF_X1 input95 (.A(b[37]),
    .Z(net95));
 BUF_X1 input96 (.A(b[38]),
    .Z(net96));
 BUF_X1 input97 (.A(b[39]),
    .Z(net97));
 BUF_X1 input98 (.A(b[3]),
    .Z(net98));
 BUF_X1 input99 (.A(b[40]),
    .Z(net99));
 BUF_X1 input100 (.A(b[41]),
    .Z(net100));
 BUF_X1 input101 (.A(b[42]),
    .Z(net101));
 BUF_X1 input102 (.A(b[43]),
    .Z(net102));
 BUF_X1 input103 (.A(b[44]),
    .Z(net103));
 BUF_X2 input104 (.A(b[45]),
    .Z(net104));
 BUF_X1 input105 (.A(b[46]),
    .Z(net105));
 BUF_X1 input106 (.A(b[47]),
    .Z(net106));
 BUF_X1 input107 (.A(b[48]),
    .Z(net107));
 BUF_X4 input108 (.A(b[49]),
    .Z(net108));
 BUF_X1 input109 (.A(b[4]),
    .Z(net109));
 BUF_X1 input110 (.A(b[50]),
    .Z(net110));
 BUF_X1 input111 (.A(b[51]),
    .Z(net111));
 BUF_X1 input112 (.A(b[52]),
    .Z(net112));
 BUF_X1 input113 (.A(b[53]),
    .Z(net113));
 BUF_X1 input114 (.A(b[54]),
    .Z(net114));
 BUF_X1 input115 (.A(b[55]),
    .Z(net115));
 BUF_X1 input116 (.A(b[56]),
    .Z(net116));
 BUF_X1 input117 (.A(b[57]),
    .Z(net117));
 BUF_X1 input118 (.A(b[58]),
    .Z(net118));
 BUF_X1 input119 (.A(b[59]),
    .Z(net119));
 BUF_X1 input120 (.A(b[5]),
    .Z(net120));
 BUF_X1 input121 (.A(b[60]),
    .Z(net121));
 BUF_X1 input122 (.A(b[61]),
    .Z(net122));
 BUF_X1 input123 (.A(b[62]),
    .Z(net123));
 BUF_X1 input124 (.A(b[63]),
    .Z(net124));
 BUF_X1 input125 (.A(b[6]),
    .Z(net125));
 BUF_X1 input126 (.A(b[7]),
    .Z(net126));
 BUF_X1 input127 (.A(b[8]),
    .Z(net127));
 BUF_X1 input128 (.A(b[9]),
    .Z(net128));
 BUF_X1 input129 (.A(cin),
    .Z(net129));
 BUF_X1 output130 (.A(net130),
    .Z(cout));
 BUF_X1 output131 (.A(net131),
    .Z(sum[0]));
 BUF_X1 output132 (.A(net132),
    .Z(sum[10]));
 BUF_X1 output133 (.A(net133),
    .Z(sum[11]));
 BUF_X1 output134 (.A(net134),
    .Z(sum[12]));
 BUF_X1 output135 (.A(net135),
    .Z(sum[13]));
 BUF_X1 output136 (.A(net136),
    .Z(sum[14]));
 BUF_X1 output137 (.A(net137),
    .Z(sum[15]));
 BUF_X1 output138 (.A(net138),
    .Z(sum[16]));
 BUF_X1 output139 (.A(net139),
    .Z(sum[17]));
 BUF_X1 output140 (.A(net140),
    .Z(sum[18]));
 BUF_X1 output141 (.A(net141),
    .Z(sum[19]));
 BUF_X1 output142 (.A(net142),
    .Z(sum[1]));
 BUF_X1 output143 (.A(net143),
    .Z(sum[20]));
 BUF_X1 output144 (.A(net144),
    .Z(sum[21]));
 BUF_X1 output145 (.A(net145),
    .Z(sum[22]));
 BUF_X1 output146 (.A(net146),
    .Z(sum[23]));
 BUF_X1 output147 (.A(net147),
    .Z(sum[24]));
 BUF_X1 output148 (.A(net148),
    .Z(sum[25]));
 BUF_X1 output149 (.A(net149),
    .Z(sum[26]));
 BUF_X1 output150 (.A(net150),
    .Z(sum[27]));
 BUF_X1 output151 (.A(net151),
    .Z(sum[28]));
 BUF_X1 output152 (.A(net152),
    .Z(sum[29]));
 BUF_X1 output153 (.A(net153),
    .Z(sum[2]));
 BUF_X1 output154 (.A(net154),
    .Z(sum[30]));
 BUF_X1 output155 (.A(net155),
    .Z(sum[31]));
 BUF_X1 output156 (.A(net156),
    .Z(sum[32]));
 BUF_X1 output157 (.A(net157),
    .Z(sum[33]));
 BUF_X1 output158 (.A(net158),
    .Z(sum[34]));
 BUF_X1 output159 (.A(net159),
    .Z(sum[35]));
 BUF_X1 output160 (.A(net160),
    .Z(sum[36]));
 BUF_X1 output161 (.A(net161),
    .Z(sum[37]));
 BUF_X1 output162 (.A(net162),
    .Z(sum[38]));
 BUF_X1 output163 (.A(net163),
    .Z(sum[39]));
 BUF_X1 output164 (.A(net164),
    .Z(sum[3]));
 BUF_X1 output165 (.A(net165),
    .Z(sum[40]));
 BUF_X1 output166 (.A(net166),
    .Z(sum[41]));
 BUF_X1 output167 (.A(net167),
    .Z(sum[42]));
 BUF_X1 output168 (.A(net168),
    .Z(sum[43]));
 BUF_X1 output169 (.A(net169),
    .Z(sum[44]));
 BUF_X1 output170 (.A(net170),
    .Z(sum[45]));
 BUF_X1 output171 (.A(net171),
    .Z(sum[46]));
 BUF_X1 output172 (.A(net172),
    .Z(sum[47]));
 BUF_X1 output173 (.A(net173),
    .Z(sum[48]));
 BUF_X1 output174 (.A(net174),
    .Z(sum[49]));
 BUF_X1 output175 (.A(net175),
    .Z(sum[4]));
 BUF_X1 output176 (.A(net176),
    .Z(sum[50]));
 BUF_X1 output177 (.A(net177),
    .Z(sum[51]));
 BUF_X1 output178 (.A(net178),
    .Z(sum[52]));
 BUF_X1 output179 (.A(net179),
    .Z(sum[53]));
 BUF_X1 output180 (.A(net180),
    .Z(sum[54]));
 BUF_X1 output181 (.A(net181),
    .Z(sum[55]));
 BUF_X1 output182 (.A(net182),
    .Z(sum[56]));
 BUF_X1 output183 (.A(net183),
    .Z(sum[57]));
 BUF_X1 output184 (.A(net184),
    .Z(sum[58]));
 BUF_X1 output185 (.A(net185),
    .Z(sum[59]));
 BUF_X1 output186 (.A(net186),
    .Z(sum[5]));
 BUF_X1 output187 (.A(net187),
    .Z(sum[60]));
 BUF_X1 output188 (.A(net188),
    .Z(sum[61]));
 BUF_X1 output189 (.A(net189),
    .Z(sum[62]));
 BUF_X1 output190 (.A(net190),
    .Z(sum[63]));
 BUF_X1 output191 (.A(net191),
    .Z(sum[6]));
 BUF_X1 output192 (.A(net192),
    .Z(sum[7]));
 BUF_X1 output193 (.A(net193),
    .Z(sum[8]));
 BUF_X1 output194 (.A(net194),
    .Z(sum[9]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X1 FILLER_0_792 ();
 FILLCELL_X1 FILLER_0_818 ();
 FILLCELL_X2 FILLER_0_823 ();
 FILLCELL_X1 FILLER_0_842 ();
 FILLCELL_X2 FILLER_0_873 ();
 FILLCELL_X1 FILLER_0_879 ();
 FILLCELL_X1 FILLER_0_883 ();
 FILLCELL_X2 FILLER_0_903 ();
 FILLCELL_X1 FILLER_0_905 ();
 FILLCELL_X1 FILLER_0_912 ();
 FILLCELL_X1 FILLER_0_917 ();
 FILLCELL_X2 FILLER_0_927 ();
 FILLCELL_X1 FILLER_0_929 ();
 FILLCELL_X4 FILLER_0_934 ();
 FILLCELL_X1 FILLER_0_938 ();
 FILLCELL_X4 FILLER_0_951 ();
 FILLCELL_X1 FILLER_0_955 ();
 FILLCELL_X2 FILLER_0_959 ();
 FILLCELL_X2 FILLER_0_967 ();
 FILLCELL_X1 FILLER_0_969 ();
 FILLCELL_X8 FILLER_0_982 ();
 FILLCELL_X1 FILLER_0_990 ();
 FILLCELL_X32 FILLER_0_1006 ();
 FILLCELL_X32 FILLER_0_1038 ();
 FILLCELL_X32 FILLER_0_1070 ();
 FILLCELL_X32 FILLER_0_1102 ();
 FILLCELL_X32 FILLER_0_1134 ();
 FILLCELL_X32 FILLER_0_1166 ();
 FILLCELL_X32 FILLER_0_1198 ();
 FILLCELL_X32 FILLER_0_1230 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X32 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_0_1679 ();
 FILLCELL_X32 FILLER_0_1711 ();
 FILLCELL_X32 FILLER_0_1743 ();
 FILLCELL_X16 FILLER_0_1775 ();
 FILLCELL_X4 FILLER_0_1791 ();
 FILLCELL_X2 FILLER_0_1795 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X16 FILLER_1_769 ();
 FILLCELL_X2 FILLER_1_785 ();
 FILLCELL_X1 FILLER_1_807 ();
 FILLCELL_X1 FILLER_1_833 ();
 FILLCELL_X2 FILLER_1_841 ();
 FILLCELL_X4 FILLER_1_864 ();
 FILLCELL_X1 FILLER_1_868 ();
 FILLCELL_X2 FILLER_1_902 ();
 FILLCELL_X8 FILLER_1_908 ();
 FILLCELL_X1 FILLER_1_916 ();
 FILLCELL_X2 FILLER_1_922 ();
 FILLCELL_X1 FILLER_1_924 ();
 FILLCELL_X2 FILLER_1_931 ();
 FILLCELL_X1 FILLER_1_933 ();
 FILLCELL_X8 FILLER_1_939 ();
 FILLCELL_X1 FILLER_1_947 ();
 FILLCELL_X4 FILLER_1_950 ();
 FILLCELL_X2 FILLER_1_954 ();
 FILLCELL_X4 FILLER_1_959 ();
 FILLCELL_X32 FILLER_1_1005 ();
 FILLCELL_X32 FILLER_1_1037 ();
 FILLCELL_X32 FILLER_1_1069 ();
 FILLCELL_X32 FILLER_1_1101 ();
 FILLCELL_X32 FILLER_1_1133 ();
 FILLCELL_X32 FILLER_1_1165 ();
 FILLCELL_X32 FILLER_1_1197 ();
 FILLCELL_X32 FILLER_1_1229 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X32 FILLER_1_1648 ();
 FILLCELL_X32 FILLER_1_1680 ();
 FILLCELL_X32 FILLER_1_1712 ();
 FILLCELL_X32 FILLER_1_1744 ();
 FILLCELL_X16 FILLER_1_1776 ();
 FILLCELL_X4 FILLER_1_1792 ();
 FILLCELL_X1 FILLER_1_1796 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X8 FILLER_2_792 ();
 FILLCELL_X1 FILLER_2_800 ();
 FILLCELL_X4 FILLER_2_805 ();
 FILLCELL_X2 FILLER_2_809 ();
 FILLCELL_X2 FILLER_2_814 ();
 FILLCELL_X2 FILLER_2_850 ();
 FILLCELL_X4 FILLER_2_855 ();
 FILLCELL_X1 FILLER_2_859 ();
 FILLCELL_X16 FILLER_2_866 ();
 FILLCELL_X4 FILLER_2_882 ();
 FILLCELL_X1 FILLER_2_918 ();
 FILLCELL_X16 FILLER_2_967 ();
 FILLCELL_X8 FILLER_2_983 ();
 FILLCELL_X32 FILLER_2_993 ();
 FILLCELL_X32 FILLER_2_1025 ();
 FILLCELL_X32 FILLER_2_1057 ();
 FILLCELL_X32 FILLER_2_1089 ();
 FILLCELL_X32 FILLER_2_1121 ();
 FILLCELL_X32 FILLER_2_1153 ();
 FILLCELL_X32 FILLER_2_1185 ();
 FILLCELL_X32 FILLER_2_1217 ();
 FILLCELL_X32 FILLER_2_1249 ();
 FILLCELL_X32 FILLER_2_1281 ();
 FILLCELL_X32 FILLER_2_1313 ();
 FILLCELL_X32 FILLER_2_1345 ();
 FILLCELL_X32 FILLER_2_1377 ();
 FILLCELL_X32 FILLER_2_1409 ();
 FILLCELL_X32 FILLER_2_1441 ();
 FILLCELL_X32 FILLER_2_1473 ();
 FILLCELL_X32 FILLER_2_1505 ();
 FILLCELL_X32 FILLER_2_1537 ();
 FILLCELL_X32 FILLER_2_1569 ();
 FILLCELL_X32 FILLER_2_1601 ();
 FILLCELL_X32 FILLER_2_1633 ();
 FILLCELL_X32 FILLER_2_1665 ();
 FILLCELL_X32 FILLER_2_1697 ();
 FILLCELL_X32 FILLER_2_1729 ();
 FILLCELL_X32 FILLER_2_1761 ();
 FILLCELL_X4 FILLER_2_1793 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X16 FILLER_3_769 ();
 FILLCELL_X8 FILLER_3_785 ();
 FILLCELL_X4 FILLER_3_793 ();
 FILLCELL_X1 FILLER_3_797 ();
 FILLCELL_X2 FILLER_3_804 ();
 FILLCELL_X2 FILLER_3_809 ();
 FILLCELL_X16 FILLER_3_825 ();
 FILLCELL_X2 FILLER_3_841 ();
 FILLCELL_X2 FILLER_3_846 ();
 FILLCELL_X32 FILLER_3_869 ();
 FILLCELL_X32 FILLER_3_901 ();
 FILLCELL_X32 FILLER_3_933 ();
 FILLCELL_X32 FILLER_3_965 ();
 FILLCELL_X32 FILLER_3_997 ();
 FILLCELL_X32 FILLER_3_1029 ();
 FILLCELL_X32 FILLER_3_1061 ();
 FILLCELL_X32 FILLER_3_1093 ();
 FILLCELL_X32 FILLER_3_1125 ();
 FILLCELL_X32 FILLER_3_1157 ();
 FILLCELL_X32 FILLER_3_1189 ();
 FILLCELL_X32 FILLER_3_1221 ();
 FILLCELL_X8 FILLER_3_1253 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X32 FILLER_3_1648 ();
 FILLCELL_X32 FILLER_3_1680 ();
 FILLCELL_X32 FILLER_3_1712 ();
 FILLCELL_X32 FILLER_3_1744 ();
 FILLCELL_X16 FILLER_3_1776 ();
 FILLCELL_X4 FILLER_3_1792 ();
 FILLCELL_X1 FILLER_3_1796 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X8 FILLER_4_792 ();
 FILLCELL_X4 FILLER_4_800 ();
 FILLCELL_X16 FILLER_4_814 ();
 FILLCELL_X8 FILLER_4_830 ();
 FILLCELL_X4 FILLER_4_838 ();
 FILLCELL_X1 FILLER_4_842 ();
 FILLCELL_X2 FILLER_4_855 ();
 FILLCELL_X32 FILLER_4_859 ();
 FILLCELL_X32 FILLER_4_891 ();
 FILLCELL_X32 FILLER_4_923 ();
 FILLCELL_X32 FILLER_4_955 ();
 FILLCELL_X32 FILLER_4_987 ();
 FILLCELL_X32 FILLER_4_1019 ();
 FILLCELL_X32 FILLER_4_1051 ();
 FILLCELL_X32 FILLER_4_1083 ();
 FILLCELL_X32 FILLER_4_1115 ();
 FILLCELL_X32 FILLER_4_1147 ();
 FILLCELL_X32 FILLER_4_1179 ();
 FILLCELL_X32 FILLER_4_1211 ();
 FILLCELL_X32 FILLER_4_1243 ();
 FILLCELL_X32 FILLER_4_1275 ();
 FILLCELL_X32 FILLER_4_1307 ();
 FILLCELL_X32 FILLER_4_1339 ();
 FILLCELL_X32 FILLER_4_1371 ();
 FILLCELL_X32 FILLER_4_1403 ();
 FILLCELL_X32 FILLER_4_1435 ();
 FILLCELL_X32 FILLER_4_1467 ();
 FILLCELL_X32 FILLER_4_1499 ();
 FILLCELL_X32 FILLER_4_1531 ();
 FILLCELL_X32 FILLER_4_1563 ();
 FILLCELL_X32 FILLER_4_1595 ();
 FILLCELL_X32 FILLER_4_1627 ();
 FILLCELL_X32 FILLER_4_1659 ();
 FILLCELL_X32 FILLER_4_1691 ();
 FILLCELL_X32 FILLER_4_1723 ();
 FILLCELL_X32 FILLER_4_1755 ();
 FILLCELL_X8 FILLER_4_1787 ();
 FILLCELL_X2 FILLER_4_1795 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X16 FILLER_5_801 ();
 FILLCELL_X4 FILLER_5_817 ();
 FILLCELL_X32 FILLER_5_838 ();
 FILLCELL_X32 FILLER_5_870 ();
 FILLCELL_X32 FILLER_5_902 ();
 FILLCELL_X32 FILLER_5_934 ();
 FILLCELL_X32 FILLER_5_966 ();
 FILLCELL_X32 FILLER_5_998 ();
 FILLCELL_X32 FILLER_5_1030 ();
 FILLCELL_X32 FILLER_5_1062 ();
 FILLCELL_X32 FILLER_5_1094 ();
 FILLCELL_X32 FILLER_5_1126 ();
 FILLCELL_X32 FILLER_5_1158 ();
 FILLCELL_X32 FILLER_5_1190 ();
 FILLCELL_X32 FILLER_5_1222 ();
 FILLCELL_X8 FILLER_5_1254 ();
 FILLCELL_X1 FILLER_5_1262 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X32 FILLER_5_1648 ();
 FILLCELL_X32 FILLER_5_1680 ();
 FILLCELL_X32 FILLER_5_1712 ();
 FILLCELL_X32 FILLER_5_1744 ();
 FILLCELL_X16 FILLER_5_1776 ();
 FILLCELL_X4 FILLER_5_1792 ();
 FILLCELL_X1 FILLER_5_1796 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X1 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_835 ();
 FILLCELL_X32 FILLER_6_867 ();
 FILLCELL_X32 FILLER_6_899 ();
 FILLCELL_X32 FILLER_6_931 ();
 FILLCELL_X32 FILLER_6_963 ();
 FILLCELL_X32 FILLER_6_995 ();
 FILLCELL_X32 FILLER_6_1027 ();
 FILLCELL_X32 FILLER_6_1059 ();
 FILLCELL_X32 FILLER_6_1091 ();
 FILLCELL_X32 FILLER_6_1123 ();
 FILLCELL_X32 FILLER_6_1155 ();
 FILLCELL_X32 FILLER_6_1187 ();
 FILLCELL_X32 FILLER_6_1219 ();
 FILLCELL_X32 FILLER_6_1251 ();
 FILLCELL_X32 FILLER_6_1283 ();
 FILLCELL_X32 FILLER_6_1315 ();
 FILLCELL_X32 FILLER_6_1347 ();
 FILLCELL_X32 FILLER_6_1379 ();
 FILLCELL_X32 FILLER_6_1411 ();
 FILLCELL_X32 FILLER_6_1443 ();
 FILLCELL_X32 FILLER_6_1475 ();
 FILLCELL_X32 FILLER_6_1507 ();
 FILLCELL_X32 FILLER_6_1539 ();
 FILLCELL_X32 FILLER_6_1571 ();
 FILLCELL_X32 FILLER_6_1603 ();
 FILLCELL_X32 FILLER_6_1635 ();
 FILLCELL_X32 FILLER_6_1667 ();
 FILLCELL_X32 FILLER_6_1699 ();
 FILLCELL_X32 FILLER_6_1731 ();
 FILLCELL_X32 FILLER_6_1763 ();
 FILLCELL_X2 FILLER_6_1795 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X16 FILLER_7_801 ();
 FILLCELL_X8 FILLER_7_817 ();
 FILLCELL_X2 FILLER_7_825 ();
 FILLCELL_X1 FILLER_7_827 ();
 FILLCELL_X32 FILLER_7_835 ();
 FILLCELL_X32 FILLER_7_867 ();
 FILLCELL_X32 FILLER_7_899 ();
 FILLCELL_X32 FILLER_7_931 ();
 FILLCELL_X32 FILLER_7_963 ();
 FILLCELL_X32 FILLER_7_995 ();
 FILLCELL_X32 FILLER_7_1027 ();
 FILLCELL_X32 FILLER_7_1059 ();
 FILLCELL_X32 FILLER_7_1091 ();
 FILLCELL_X32 FILLER_7_1123 ();
 FILLCELL_X32 FILLER_7_1155 ();
 FILLCELL_X32 FILLER_7_1187 ();
 FILLCELL_X32 FILLER_7_1219 ();
 FILLCELL_X8 FILLER_7_1251 ();
 FILLCELL_X4 FILLER_7_1259 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X32 FILLER_7_1648 ();
 FILLCELL_X32 FILLER_7_1680 ();
 FILLCELL_X32 FILLER_7_1712 ();
 FILLCELL_X32 FILLER_7_1744 ();
 FILLCELL_X16 FILLER_7_1776 ();
 FILLCELL_X4 FILLER_7_1792 ();
 FILLCELL_X1 FILLER_7_1796 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X4 FILLER_8_824 ();
 FILLCELL_X2 FILLER_8_837 ();
 FILLCELL_X2 FILLER_8_844 ();
 FILLCELL_X1 FILLER_8_846 ();
 FILLCELL_X32 FILLER_8_867 ();
 FILLCELL_X32 FILLER_8_899 ();
 FILLCELL_X32 FILLER_8_931 ();
 FILLCELL_X32 FILLER_8_963 ();
 FILLCELL_X32 FILLER_8_995 ();
 FILLCELL_X32 FILLER_8_1027 ();
 FILLCELL_X32 FILLER_8_1059 ();
 FILLCELL_X32 FILLER_8_1091 ();
 FILLCELL_X32 FILLER_8_1123 ();
 FILLCELL_X32 FILLER_8_1155 ();
 FILLCELL_X32 FILLER_8_1187 ();
 FILLCELL_X32 FILLER_8_1219 ();
 FILLCELL_X32 FILLER_8_1251 ();
 FILLCELL_X32 FILLER_8_1283 ();
 FILLCELL_X32 FILLER_8_1315 ();
 FILLCELL_X32 FILLER_8_1347 ();
 FILLCELL_X32 FILLER_8_1379 ();
 FILLCELL_X32 FILLER_8_1411 ();
 FILLCELL_X32 FILLER_8_1443 ();
 FILLCELL_X32 FILLER_8_1475 ();
 FILLCELL_X32 FILLER_8_1507 ();
 FILLCELL_X32 FILLER_8_1539 ();
 FILLCELL_X32 FILLER_8_1571 ();
 FILLCELL_X32 FILLER_8_1603 ();
 FILLCELL_X32 FILLER_8_1635 ();
 FILLCELL_X32 FILLER_8_1667 ();
 FILLCELL_X32 FILLER_8_1699 ();
 FILLCELL_X32 FILLER_8_1731 ();
 FILLCELL_X32 FILLER_8_1763 ();
 FILLCELL_X2 FILLER_8_1795 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X16 FILLER_9_801 ();
 FILLCELL_X8 FILLER_9_817 ();
 FILLCELL_X4 FILLER_9_825 ();
 FILLCELL_X8 FILLER_9_840 ();
 FILLCELL_X32 FILLER_9_858 ();
 FILLCELL_X32 FILLER_9_890 ();
 FILLCELL_X32 FILLER_9_922 ();
 FILLCELL_X32 FILLER_9_954 ();
 FILLCELL_X32 FILLER_9_986 ();
 FILLCELL_X32 FILLER_9_1018 ();
 FILLCELL_X32 FILLER_9_1050 ();
 FILLCELL_X32 FILLER_9_1082 ();
 FILLCELL_X32 FILLER_9_1114 ();
 FILLCELL_X32 FILLER_9_1146 ();
 FILLCELL_X32 FILLER_9_1178 ();
 FILLCELL_X32 FILLER_9_1210 ();
 FILLCELL_X16 FILLER_9_1242 ();
 FILLCELL_X4 FILLER_9_1258 ();
 FILLCELL_X1 FILLER_9_1262 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X32 FILLER_9_1648 ();
 FILLCELL_X32 FILLER_9_1680 ();
 FILLCELL_X32 FILLER_9_1712 ();
 FILLCELL_X32 FILLER_9_1744 ();
 FILLCELL_X16 FILLER_9_1776 ();
 FILLCELL_X4 FILLER_9_1792 ();
 FILLCELL_X1 FILLER_9_1796 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X2 FILLER_10_824 ();
 FILLCELL_X1 FILLER_10_826 ();
 FILLCELL_X8 FILLER_10_840 ();
 FILLCELL_X1 FILLER_10_848 ();
 FILLCELL_X32 FILLER_10_859 ();
 FILLCELL_X32 FILLER_10_891 ();
 FILLCELL_X32 FILLER_10_923 ();
 FILLCELL_X32 FILLER_10_955 ();
 FILLCELL_X32 FILLER_10_987 ();
 FILLCELL_X32 FILLER_10_1019 ();
 FILLCELL_X32 FILLER_10_1051 ();
 FILLCELL_X32 FILLER_10_1083 ();
 FILLCELL_X32 FILLER_10_1115 ();
 FILLCELL_X32 FILLER_10_1147 ();
 FILLCELL_X32 FILLER_10_1179 ();
 FILLCELL_X32 FILLER_10_1211 ();
 FILLCELL_X32 FILLER_10_1243 ();
 FILLCELL_X32 FILLER_10_1275 ();
 FILLCELL_X32 FILLER_10_1307 ();
 FILLCELL_X32 FILLER_10_1339 ();
 FILLCELL_X32 FILLER_10_1371 ();
 FILLCELL_X32 FILLER_10_1403 ();
 FILLCELL_X32 FILLER_10_1435 ();
 FILLCELL_X32 FILLER_10_1467 ();
 FILLCELL_X32 FILLER_10_1499 ();
 FILLCELL_X32 FILLER_10_1531 ();
 FILLCELL_X32 FILLER_10_1563 ();
 FILLCELL_X32 FILLER_10_1595 ();
 FILLCELL_X32 FILLER_10_1627 ();
 FILLCELL_X32 FILLER_10_1659 ();
 FILLCELL_X32 FILLER_10_1691 ();
 FILLCELL_X32 FILLER_10_1723 ();
 FILLCELL_X32 FILLER_10_1755 ();
 FILLCELL_X8 FILLER_10_1787 ();
 FILLCELL_X2 FILLER_10_1795 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X8 FILLER_11_833 ();
 FILLCELL_X4 FILLER_11_841 ();
 FILLCELL_X2 FILLER_11_845 ();
 FILLCELL_X1 FILLER_11_847 ();
 FILLCELL_X32 FILLER_11_864 ();
 FILLCELL_X32 FILLER_11_896 ();
 FILLCELL_X32 FILLER_11_928 ();
 FILLCELL_X32 FILLER_11_960 ();
 FILLCELL_X32 FILLER_11_992 ();
 FILLCELL_X32 FILLER_11_1024 ();
 FILLCELL_X32 FILLER_11_1056 ();
 FILLCELL_X32 FILLER_11_1088 ();
 FILLCELL_X32 FILLER_11_1120 ();
 FILLCELL_X32 FILLER_11_1152 ();
 FILLCELL_X32 FILLER_11_1184 ();
 FILLCELL_X32 FILLER_11_1216 ();
 FILLCELL_X8 FILLER_11_1248 ();
 FILLCELL_X4 FILLER_11_1256 ();
 FILLCELL_X2 FILLER_11_1260 ();
 FILLCELL_X1 FILLER_11_1262 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X32 FILLER_11_1648 ();
 FILLCELL_X32 FILLER_11_1680 ();
 FILLCELL_X32 FILLER_11_1712 ();
 FILLCELL_X32 FILLER_11_1744 ();
 FILLCELL_X16 FILLER_11_1776 ();
 FILLCELL_X4 FILLER_11_1792 ();
 FILLCELL_X1 FILLER_11_1796 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X32 FILLER_12_1592 ();
 FILLCELL_X32 FILLER_12_1624 ();
 FILLCELL_X32 FILLER_12_1656 ();
 FILLCELL_X32 FILLER_12_1688 ();
 FILLCELL_X32 FILLER_12_1720 ();
 FILLCELL_X32 FILLER_12_1752 ();
 FILLCELL_X8 FILLER_12_1784 ();
 FILLCELL_X4 FILLER_12_1792 ();
 FILLCELL_X1 FILLER_12_1796 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X32 FILLER_13_1648 ();
 FILLCELL_X32 FILLER_13_1680 ();
 FILLCELL_X32 FILLER_13_1712 ();
 FILLCELL_X32 FILLER_13_1744 ();
 FILLCELL_X16 FILLER_13_1776 ();
 FILLCELL_X4 FILLER_13_1792 ();
 FILLCELL_X1 FILLER_13_1796 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X32 FILLER_14_1688 ();
 FILLCELL_X32 FILLER_14_1720 ();
 FILLCELL_X32 FILLER_14_1752 ();
 FILLCELL_X8 FILLER_14_1784 ();
 FILLCELL_X4 FILLER_14_1792 ();
 FILLCELL_X1 FILLER_14_1796 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X32 FILLER_15_1584 ();
 FILLCELL_X32 FILLER_15_1616 ();
 FILLCELL_X32 FILLER_15_1648 ();
 FILLCELL_X32 FILLER_15_1680 ();
 FILLCELL_X32 FILLER_15_1712 ();
 FILLCELL_X32 FILLER_15_1744 ();
 FILLCELL_X16 FILLER_15_1776 ();
 FILLCELL_X4 FILLER_15_1792 ();
 FILLCELL_X1 FILLER_15_1796 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X32 FILLER_16_1592 ();
 FILLCELL_X32 FILLER_16_1624 ();
 FILLCELL_X32 FILLER_16_1656 ();
 FILLCELL_X32 FILLER_16_1688 ();
 FILLCELL_X32 FILLER_16_1720 ();
 FILLCELL_X32 FILLER_16_1752 ();
 FILLCELL_X8 FILLER_16_1784 ();
 FILLCELL_X4 FILLER_16_1792 ();
 FILLCELL_X1 FILLER_16_1796 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X32 FILLER_17_1584 ();
 FILLCELL_X32 FILLER_17_1616 ();
 FILLCELL_X32 FILLER_17_1648 ();
 FILLCELL_X32 FILLER_17_1680 ();
 FILLCELL_X32 FILLER_17_1712 ();
 FILLCELL_X32 FILLER_17_1744 ();
 FILLCELL_X16 FILLER_17_1776 ();
 FILLCELL_X4 FILLER_17_1792 ();
 FILLCELL_X1 FILLER_17_1796 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X32 FILLER_18_1752 ();
 FILLCELL_X8 FILLER_18_1784 ();
 FILLCELL_X4 FILLER_18_1792 ();
 FILLCELL_X1 FILLER_18_1796 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X32 FILLER_19_1584 ();
 FILLCELL_X32 FILLER_19_1616 ();
 FILLCELL_X32 FILLER_19_1648 ();
 FILLCELL_X32 FILLER_19_1680 ();
 FILLCELL_X32 FILLER_19_1712 ();
 FILLCELL_X32 FILLER_19_1744 ();
 FILLCELL_X16 FILLER_19_1776 ();
 FILLCELL_X4 FILLER_19_1792 ();
 FILLCELL_X1 FILLER_19_1796 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X32 FILLER_20_1592 ();
 FILLCELL_X32 FILLER_20_1624 ();
 FILLCELL_X32 FILLER_20_1656 ();
 FILLCELL_X32 FILLER_20_1688 ();
 FILLCELL_X32 FILLER_20_1720 ();
 FILLCELL_X32 FILLER_20_1752 ();
 FILLCELL_X8 FILLER_20_1784 ();
 FILLCELL_X4 FILLER_20_1792 ();
 FILLCELL_X1 FILLER_20_1796 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X32 FILLER_21_1744 ();
 FILLCELL_X16 FILLER_21_1776 ();
 FILLCELL_X4 FILLER_21_1792 ();
 FILLCELL_X1 FILLER_21_1796 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X32 FILLER_22_1752 ();
 FILLCELL_X8 FILLER_22_1784 ();
 FILLCELL_X4 FILLER_22_1792 ();
 FILLCELL_X1 FILLER_22_1796 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X32 FILLER_23_1584 ();
 FILLCELL_X32 FILLER_23_1616 ();
 FILLCELL_X32 FILLER_23_1648 ();
 FILLCELL_X32 FILLER_23_1680 ();
 FILLCELL_X32 FILLER_23_1712 ();
 FILLCELL_X32 FILLER_23_1744 ();
 FILLCELL_X16 FILLER_23_1776 ();
 FILLCELL_X4 FILLER_23_1792 ();
 FILLCELL_X1 FILLER_23_1796 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X32 FILLER_24_1592 ();
 FILLCELL_X32 FILLER_24_1624 ();
 FILLCELL_X32 FILLER_24_1656 ();
 FILLCELL_X32 FILLER_24_1688 ();
 FILLCELL_X32 FILLER_24_1720 ();
 FILLCELL_X32 FILLER_24_1752 ();
 FILLCELL_X8 FILLER_24_1784 ();
 FILLCELL_X4 FILLER_24_1792 ();
 FILLCELL_X1 FILLER_24_1796 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X32 FILLER_25_1584 ();
 FILLCELL_X32 FILLER_25_1616 ();
 FILLCELL_X32 FILLER_25_1648 ();
 FILLCELL_X32 FILLER_25_1680 ();
 FILLCELL_X32 FILLER_25_1712 ();
 FILLCELL_X32 FILLER_25_1744 ();
 FILLCELL_X16 FILLER_25_1776 ();
 FILLCELL_X4 FILLER_25_1792 ();
 FILLCELL_X1 FILLER_25_1796 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X32 FILLER_26_1592 ();
 FILLCELL_X32 FILLER_26_1624 ();
 FILLCELL_X32 FILLER_26_1656 ();
 FILLCELL_X32 FILLER_26_1688 ();
 FILLCELL_X32 FILLER_26_1720 ();
 FILLCELL_X32 FILLER_26_1752 ();
 FILLCELL_X8 FILLER_26_1784 ();
 FILLCELL_X4 FILLER_26_1792 ();
 FILLCELL_X1 FILLER_26_1796 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X32 FILLER_27_1584 ();
 FILLCELL_X32 FILLER_27_1616 ();
 FILLCELL_X32 FILLER_27_1648 ();
 FILLCELL_X32 FILLER_27_1680 ();
 FILLCELL_X32 FILLER_27_1712 ();
 FILLCELL_X32 FILLER_27_1744 ();
 FILLCELL_X16 FILLER_27_1776 ();
 FILLCELL_X4 FILLER_27_1792 ();
 FILLCELL_X1 FILLER_27_1796 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X32 FILLER_28_1592 ();
 FILLCELL_X32 FILLER_28_1624 ();
 FILLCELL_X32 FILLER_28_1656 ();
 FILLCELL_X32 FILLER_28_1688 ();
 FILLCELL_X32 FILLER_28_1720 ();
 FILLCELL_X32 FILLER_28_1752 ();
 FILLCELL_X8 FILLER_28_1784 ();
 FILLCELL_X4 FILLER_28_1792 ();
 FILLCELL_X1 FILLER_28_1796 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X32 FILLER_29_1584 ();
 FILLCELL_X32 FILLER_29_1616 ();
 FILLCELL_X32 FILLER_29_1648 ();
 FILLCELL_X32 FILLER_29_1680 ();
 FILLCELL_X32 FILLER_29_1712 ();
 FILLCELL_X32 FILLER_29_1744 ();
 FILLCELL_X16 FILLER_29_1776 ();
 FILLCELL_X4 FILLER_29_1792 ();
 FILLCELL_X1 FILLER_29_1796 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X32 FILLER_30_1592 ();
 FILLCELL_X32 FILLER_30_1624 ();
 FILLCELL_X32 FILLER_30_1656 ();
 FILLCELL_X32 FILLER_30_1688 ();
 FILLCELL_X32 FILLER_30_1720 ();
 FILLCELL_X32 FILLER_30_1752 ();
 FILLCELL_X8 FILLER_30_1784 ();
 FILLCELL_X4 FILLER_30_1792 ();
 FILLCELL_X1 FILLER_30_1796 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X32 FILLER_31_1584 ();
 FILLCELL_X32 FILLER_31_1616 ();
 FILLCELL_X32 FILLER_31_1648 ();
 FILLCELL_X32 FILLER_31_1680 ();
 FILLCELL_X32 FILLER_31_1712 ();
 FILLCELL_X32 FILLER_31_1744 ();
 FILLCELL_X16 FILLER_31_1776 ();
 FILLCELL_X4 FILLER_31_1792 ();
 FILLCELL_X1 FILLER_31_1796 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X32 FILLER_32_1592 ();
 FILLCELL_X32 FILLER_32_1624 ();
 FILLCELL_X32 FILLER_32_1656 ();
 FILLCELL_X32 FILLER_32_1688 ();
 FILLCELL_X32 FILLER_32_1720 ();
 FILLCELL_X32 FILLER_32_1752 ();
 FILLCELL_X8 FILLER_32_1784 ();
 FILLCELL_X4 FILLER_32_1792 ();
 FILLCELL_X1 FILLER_32_1796 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X32 FILLER_33_1584 ();
 FILLCELL_X32 FILLER_33_1616 ();
 FILLCELL_X32 FILLER_33_1648 ();
 FILLCELL_X32 FILLER_33_1680 ();
 FILLCELL_X32 FILLER_33_1712 ();
 FILLCELL_X32 FILLER_33_1744 ();
 FILLCELL_X16 FILLER_33_1776 ();
 FILLCELL_X4 FILLER_33_1792 ();
 FILLCELL_X1 FILLER_33_1796 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X32 FILLER_34_1592 ();
 FILLCELL_X32 FILLER_34_1624 ();
 FILLCELL_X32 FILLER_34_1656 ();
 FILLCELL_X32 FILLER_34_1688 ();
 FILLCELL_X32 FILLER_34_1720 ();
 FILLCELL_X32 FILLER_34_1752 ();
 FILLCELL_X8 FILLER_34_1784 ();
 FILLCELL_X4 FILLER_34_1792 ();
 FILLCELL_X1 FILLER_34_1796 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X32 FILLER_35_1584 ();
 FILLCELL_X32 FILLER_35_1616 ();
 FILLCELL_X32 FILLER_35_1648 ();
 FILLCELL_X32 FILLER_35_1680 ();
 FILLCELL_X32 FILLER_35_1712 ();
 FILLCELL_X32 FILLER_35_1744 ();
 FILLCELL_X16 FILLER_35_1776 ();
 FILLCELL_X4 FILLER_35_1792 ();
 FILLCELL_X1 FILLER_35_1796 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X32 FILLER_36_1592 ();
 FILLCELL_X32 FILLER_36_1624 ();
 FILLCELL_X32 FILLER_36_1656 ();
 FILLCELL_X32 FILLER_36_1688 ();
 FILLCELL_X32 FILLER_36_1720 ();
 FILLCELL_X32 FILLER_36_1752 ();
 FILLCELL_X8 FILLER_36_1784 ();
 FILLCELL_X4 FILLER_36_1792 ();
 FILLCELL_X1 FILLER_36_1796 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X32 FILLER_37_1584 ();
 FILLCELL_X32 FILLER_37_1616 ();
 FILLCELL_X32 FILLER_37_1648 ();
 FILLCELL_X32 FILLER_37_1680 ();
 FILLCELL_X32 FILLER_37_1712 ();
 FILLCELL_X32 FILLER_37_1744 ();
 FILLCELL_X16 FILLER_37_1776 ();
 FILLCELL_X4 FILLER_37_1792 ();
 FILLCELL_X1 FILLER_37_1796 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X32 FILLER_38_1592 ();
 FILLCELL_X32 FILLER_38_1624 ();
 FILLCELL_X32 FILLER_38_1656 ();
 FILLCELL_X32 FILLER_38_1688 ();
 FILLCELL_X32 FILLER_38_1720 ();
 FILLCELL_X32 FILLER_38_1752 ();
 FILLCELL_X8 FILLER_38_1784 ();
 FILLCELL_X4 FILLER_38_1792 ();
 FILLCELL_X1 FILLER_38_1796 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X32 FILLER_39_1584 ();
 FILLCELL_X32 FILLER_39_1616 ();
 FILLCELL_X32 FILLER_39_1648 ();
 FILLCELL_X32 FILLER_39_1680 ();
 FILLCELL_X32 FILLER_39_1712 ();
 FILLCELL_X32 FILLER_39_1744 ();
 FILLCELL_X16 FILLER_39_1776 ();
 FILLCELL_X4 FILLER_39_1792 ();
 FILLCELL_X1 FILLER_39_1796 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X32 FILLER_40_1592 ();
 FILLCELL_X32 FILLER_40_1624 ();
 FILLCELL_X32 FILLER_40_1656 ();
 FILLCELL_X32 FILLER_40_1688 ();
 FILLCELL_X32 FILLER_40_1720 ();
 FILLCELL_X32 FILLER_40_1752 ();
 FILLCELL_X8 FILLER_40_1784 ();
 FILLCELL_X4 FILLER_40_1792 ();
 FILLCELL_X1 FILLER_40_1796 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X32 FILLER_41_1584 ();
 FILLCELL_X32 FILLER_41_1616 ();
 FILLCELL_X32 FILLER_41_1648 ();
 FILLCELL_X32 FILLER_41_1680 ();
 FILLCELL_X32 FILLER_41_1712 ();
 FILLCELL_X32 FILLER_41_1744 ();
 FILLCELL_X16 FILLER_41_1776 ();
 FILLCELL_X4 FILLER_41_1792 ();
 FILLCELL_X1 FILLER_41_1796 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X32 FILLER_42_1592 ();
 FILLCELL_X32 FILLER_42_1624 ();
 FILLCELL_X32 FILLER_42_1656 ();
 FILLCELL_X32 FILLER_42_1688 ();
 FILLCELL_X32 FILLER_42_1720 ();
 FILLCELL_X32 FILLER_42_1752 ();
 FILLCELL_X8 FILLER_42_1784 ();
 FILLCELL_X4 FILLER_42_1792 ();
 FILLCELL_X1 FILLER_42_1796 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X32 FILLER_43_1584 ();
 FILLCELL_X32 FILLER_43_1616 ();
 FILLCELL_X32 FILLER_43_1648 ();
 FILLCELL_X32 FILLER_43_1680 ();
 FILLCELL_X32 FILLER_43_1712 ();
 FILLCELL_X32 FILLER_43_1744 ();
 FILLCELL_X16 FILLER_43_1776 ();
 FILLCELL_X4 FILLER_43_1792 ();
 FILLCELL_X1 FILLER_43_1796 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X32 FILLER_44_1592 ();
 FILLCELL_X32 FILLER_44_1624 ();
 FILLCELL_X32 FILLER_44_1656 ();
 FILLCELL_X32 FILLER_44_1688 ();
 FILLCELL_X32 FILLER_44_1720 ();
 FILLCELL_X32 FILLER_44_1752 ();
 FILLCELL_X8 FILLER_44_1784 ();
 FILLCELL_X4 FILLER_44_1792 ();
 FILLCELL_X1 FILLER_44_1796 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X32 FILLER_45_1584 ();
 FILLCELL_X32 FILLER_45_1616 ();
 FILLCELL_X32 FILLER_45_1648 ();
 FILLCELL_X32 FILLER_45_1680 ();
 FILLCELL_X32 FILLER_45_1712 ();
 FILLCELL_X32 FILLER_45_1744 ();
 FILLCELL_X16 FILLER_45_1776 ();
 FILLCELL_X4 FILLER_45_1792 ();
 FILLCELL_X1 FILLER_45_1796 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X32 FILLER_46_1592 ();
 FILLCELL_X32 FILLER_46_1624 ();
 FILLCELL_X32 FILLER_46_1656 ();
 FILLCELL_X32 FILLER_46_1688 ();
 FILLCELL_X32 FILLER_46_1720 ();
 FILLCELL_X32 FILLER_46_1752 ();
 FILLCELL_X8 FILLER_46_1784 ();
 FILLCELL_X4 FILLER_46_1792 ();
 FILLCELL_X1 FILLER_46_1796 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X32 FILLER_47_1584 ();
 FILLCELL_X32 FILLER_47_1616 ();
 FILLCELL_X32 FILLER_47_1648 ();
 FILLCELL_X32 FILLER_47_1680 ();
 FILLCELL_X32 FILLER_47_1712 ();
 FILLCELL_X32 FILLER_47_1744 ();
 FILLCELL_X16 FILLER_47_1776 ();
 FILLCELL_X4 FILLER_47_1792 ();
 FILLCELL_X1 FILLER_47_1796 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X32 FILLER_48_1592 ();
 FILLCELL_X32 FILLER_48_1624 ();
 FILLCELL_X32 FILLER_48_1656 ();
 FILLCELL_X32 FILLER_48_1688 ();
 FILLCELL_X32 FILLER_48_1720 ();
 FILLCELL_X32 FILLER_48_1752 ();
 FILLCELL_X8 FILLER_48_1784 ();
 FILLCELL_X4 FILLER_48_1792 ();
 FILLCELL_X1 FILLER_48_1796 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X32 FILLER_49_1584 ();
 FILLCELL_X32 FILLER_49_1616 ();
 FILLCELL_X32 FILLER_49_1648 ();
 FILLCELL_X32 FILLER_49_1680 ();
 FILLCELL_X32 FILLER_49_1712 ();
 FILLCELL_X32 FILLER_49_1744 ();
 FILLCELL_X16 FILLER_49_1776 ();
 FILLCELL_X4 FILLER_49_1792 ();
 FILLCELL_X1 FILLER_49_1796 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X32 FILLER_50_1592 ();
 FILLCELL_X32 FILLER_50_1624 ();
 FILLCELL_X32 FILLER_50_1656 ();
 FILLCELL_X32 FILLER_50_1688 ();
 FILLCELL_X32 FILLER_50_1720 ();
 FILLCELL_X32 FILLER_50_1752 ();
 FILLCELL_X8 FILLER_50_1784 ();
 FILLCELL_X4 FILLER_50_1792 ();
 FILLCELL_X1 FILLER_50_1796 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X32 FILLER_51_1584 ();
 FILLCELL_X32 FILLER_51_1616 ();
 FILLCELL_X32 FILLER_51_1648 ();
 FILLCELL_X32 FILLER_51_1680 ();
 FILLCELL_X32 FILLER_51_1712 ();
 FILLCELL_X32 FILLER_51_1744 ();
 FILLCELL_X16 FILLER_51_1776 ();
 FILLCELL_X4 FILLER_51_1792 ();
 FILLCELL_X1 FILLER_51_1796 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X32 FILLER_52_1592 ();
 FILLCELL_X32 FILLER_52_1624 ();
 FILLCELL_X32 FILLER_52_1656 ();
 FILLCELL_X32 FILLER_52_1688 ();
 FILLCELL_X32 FILLER_52_1720 ();
 FILLCELL_X32 FILLER_52_1752 ();
 FILLCELL_X8 FILLER_52_1784 ();
 FILLCELL_X4 FILLER_52_1792 ();
 FILLCELL_X1 FILLER_52_1796 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X32 FILLER_53_1584 ();
 FILLCELL_X32 FILLER_53_1616 ();
 FILLCELL_X32 FILLER_53_1648 ();
 FILLCELL_X32 FILLER_53_1680 ();
 FILLCELL_X32 FILLER_53_1712 ();
 FILLCELL_X32 FILLER_53_1744 ();
 FILLCELL_X16 FILLER_53_1776 ();
 FILLCELL_X4 FILLER_53_1792 ();
 FILLCELL_X1 FILLER_53_1796 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X32 FILLER_54_1592 ();
 FILLCELL_X32 FILLER_54_1624 ();
 FILLCELL_X32 FILLER_54_1656 ();
 FILLCELL_X32 FILLER_54_1688 ();
 FILLCELL_X32 FILLER_54_1720 ();
 FILLCELL_X32 FILLER_54_1752 ();
 FILLCELL_X8 FILLER_54_1784 ();
 FILLCELL_X4 FILLER_54_1792 ();
 FILLCELL_X1 FILLER_54_1796 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X32 FILLER_55_1584 ();
 FILLCELL_X32 FILLER_55_1616 ();
 FILLCELL_X32 FILLER_55_1648 ();
 FILLCELL_X32 FILLER_55_1680 ();
 FILLCELL_X32 FILLER_55_1712 ();
 FILLCELL_X32 FILLER_55_1744 ();
 FILLCELL_X16 FILLER_55_1776 ();
 FILLCELL_X4 FILLER_55_1792 ();
 FILLCELL_X1 FILLER_55_1796 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X32 FILLER_56_1592 ();
 FILLCELL_X32 FILLER_56_1624 ();
 FILLCELL_X32 FILLER_56_1656 ();
 FILLCELL_X32 FILLER_56_1688 ();
 FILLCELL_X32 FILLER_56_1720 ();
 FILLCELL_X32 FILLER_56_1752 ();
 FILLCELL_X8 FILLER_56_1784 ();
 FILLCELL_X4 FILLER_56_1792 ();
 FILLCELL_X1 FILLER_56_1796 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X32 FILLER_57_1584 ();
 FILLCELL_X32 FILLER_57_1616 ();
 FILLCELL_X32 FILLER_57_1648 ();
 FILLCELL_X32 FILLER_57_1680 ();
 FILLCELL_X32 FILLER_57_1712 ();
 FILLCELL_X32 FILLER_57_1744 ();
 FILLCELL_X16 FILLER_57_1776 ();
 FILLCELL_X4 FILLER_57_1792 ();
 FILLCELL_X1 FILLER_57_1796 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X32 FILLER_58_1592 ();
 FILLCELL_X32 FILLER_58_1624 ();
 FILLCELL_X32 FILLER_58_1656 ();
 FILLCELL_X32 FILLER_58_1688 ();
 FILLCELL_X32 FILLER_58_1720 ();
 FILLCELL_X32 FILLER_58_1752 ();
 FILLCELL_X8 FILLER_58_1784 ();
 FILLCELL_X4 FILLER_58_1792 ();
 FILLCELL_X1 FILLER_58_1796 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X32 FILLER_59_1584 ();
 FILLCELL_X32 FILLER_59_1616 ();
 FILLCELL_X32 FILLER_59_1648 ();
 FILLCELL_X32 FILLER_59_1680 ();
 FILLCELL_X32 FILLER_59_1712 ();
 FILLCELL_X32 FILLER_59_1744 ();
 FILLCELL_X16 FILLER_59_1776 ();
 FILLCELL_X4 FILLER_59_1792 ();
 FILLCELL_X1 FILLER_59_1796 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X32 FILLER_60_1592 ();
 FILLCELL_X32 FILLER_60_1624 ();
 FILLCELL_X32 FILLER_60_1656 ();
 FILLCELL_X32 FILLER_60_1688 ();
 FILLCELL_X32 FILLER_60_1720 ();
 FILLCELL_X32 FILLER_60_1752 ();
 FILLCELL_X8 FILLER_60_1784 ();
 FILLCELL_X4 FILLER_60_1792 ();
 FILLCELL_X1 FILLER_60_1796 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X32 FILLER_61_1584 ();
 FILLCELL_X32 FILLER_61_1616 ();
 FILLCELL_X32 FILLER_61_1648 ();
 FILLCELL_X32 FILLER_61_1680 ();
 FILLCELL_X32 FILLER_61_1712 ();
 FILLCELL_X32 FILLER_61_1744 ();
 FILLCELL_X16 FILLER_61_1776 ();
 FILLCELL_X4 FILLER_61_1792 ();
 FILLCELL_X1 FILLER_61_1796 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X32 FILLER_62_1592 ();
 FILLCELL_X32 FILLER_62_1624 ();
 FILLCELL_X32 FILLER_62_1656 ();
 FILLCELL_X32 FILLER_62_1688 ();
 FILLCELL_X32 FILLER_62_1720 ();
 FILLCELL_X32 FILLER_62_1752 ();
 FILLCELL_X8 FILLER_62_1784 ();
 FILLCELL_X4 FILLER_62_1792 ();
 FILLCELL_X1 FILLER_62_1796 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X32 FILLER_63_1584 ();
 FILLCELL_X32 FILLER_63_1616 ();
 FILLCELL_X32 FILLER_63_1648 ();
 FILLCELL_X32 FILLER_63_1680 ();
 FILLCELL_X32 FILLER_63_1712 ();
 FILLCELL_X32 FILLER_63_1744 ();
 FILLCELL_X16 FILLER_63_1776 ();
 FILLCELL_X4 FILLER_63_1792 ();
 FILLCELL_X1 FILLER_63_1796 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X32 FILLER_64_1592 ();
 FILLCELL_X32 FILLER_64_1624 ();
 FILLCELL_X32 FILLER_64_1656 ();
 FILLCELL_X32 FILLER_64_1688 ();
 FILLCELL_X32 FILLER_64_1720 ();
 FILLCELL_X32 FILLER_64_1752 ();
 FILLCELL_X8 FILLER_64_1784 ();
 FILLCELL_X4 FILLER_64_1792 ();
 FILLCELL_X1 FILLER_64_1796 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X32 FILLER_65_1584 ();
 FILLCELL_X32 FILLER_65_1616 ();
 FILLCELL_X32 FILLER_65_1648 ();
 FILLCELL_X32 FILLER_65_1680 ();
 FILLCELL_X32 FILLER_65_1712 ();
 FILLCELL_X32 FILLER_65_1744 ();
 FILLCELL_X16 FILLER_65_1776 ();
 FILLCELL_X4 FILLER_65_1792 ();
 FILLCELL_X1 FILLER_65_1796 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X32 FILLER_66_1592 ();
 FILLCELL_X32 FILLER_66_1624 ();
 FILLCELL_X32 FILLER_66_1656 ();
 FILLCELL_X32 FILLER_66_1688 ();
 FILLCELL_X32 FILLER_66_1720 ();
 FILLCELL_X32 FILLER_66_1752 ();
 FILLCELL_X8 FILLER_66_1784 ();
 FILLCELL_X4 FILLER_66_1792 ();
 FILLCELL_X1 FILLER_66_1796 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X16 FILLER_67_801 ();
 FILLCELL_X8 FILLER_67_817 ();
 FILLCELL_X32 FILLER_67_832 ();
 FILLCELL_X32 FILLER_67_864 ();
 FILLCELL_X32 FILLER_67_896 ();
 FILLCELL_X32 FILLER_67_928 ();
 FILLCELL_X32 FILLER_67_960 ();
 FILLCELL_X32 FILLER_67_992 ();
 FILLCELL_X32 FILLER_67_1024 ();
 FILLCELL_X32 FILLER_67_1056 ();
 FILLCELL_X32 FILLER_67_1088 ();
 FILLCELL_X32 FILLER_67_1120 ();
 FILLCELL_X32 FILLER_67_1152 ();
 FILLCELL_X32 FILLER_67_1184 ();
 FILLCELL_X32 FILLER_67_1216 ();
 FILLCELL_X8 FILLER_67_1248 ();
 FILLCELL_X4 FILLER_67_1256 ();
 FILLCELL_X2 FILLER_67_1260 ();
 FILLCELL_X1 FILLER_67_1262 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X32 FILLER_67_1584 ();
 FILLCELL_X32 FILLER_67_1616 ();
 FILLCELL_X32 FILLER_67_1648 ();
 FILLCELL_X32 FILLER_67_1680 ();
 FILLCELL_X32 FILLER_67_1712 ();
 FILLCELL_X32 FILLER_67_1744 ();
 FILLCELL_X16 FILLER_67_1776 ();
 FILLCELL_X4 FILLER_67_1792 ();
 FILLCELL_X1 FILLER_67_1796 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X16 FILLER_68_792 ();
 FILLCELL_X8 FILLER_68_808 ();
 FILLCELL_X4 FILLER_68_816 ();
 FILLCELL_X1 FILLER_68_820 ();
 FILLCELL_X32 FILLER_68_839 ();
 FILLCELL_X32 FILLER_68_871 ();
 FILLCELL_X32 FILLER_68_903 ();
 FILLCELL_X32 FILLER_68_935 ();
 FILLCELL_X32 FILLER_68_967 ();
 FILLCELL_X32 FILLER_68_999 ();
 FILLCELL_X32 FILLER_68_1031 ();
 FILLCELL_X32 FILLER_68_1063 ();
 FILLCELL_X32 FILLER_68_1095 ();
 FILLCELL_X32 FILLER_68_1127 ();
 FILLCELL_X32 FILLER_68_1159 ();
 FILLCELL_X32 FILLER_68_1191 ();
 FILLCELL_X32 FILLER_68_1223 ();
 FILLCELL_X32 FILLER_68_1255 ();
 FILLCELL_X32 FILLER_68_1287 ();
 FILLCELL_X32 FILLER_68_1319 ();
 FILLCELL_X32 FILLER_68_1351 ();
 FILLCELL_X32 FILLER_68_1383 ();
 FILLCELL_X32 FILLER_68_1415 ();
 FILLCELL_X32 FILLER_68_1447 ();
 FILLCELL_X32 FILLER_68_1479 ();
 FILLCELL_X32 FILLER_68_1511 ();
 FILLCELL_X32 FILLER_68_1543 ();
 FILLCELL_X32 FILLER_68_1575 ();
 FILLCELL_X32 FILLER_68_1607 ();
 FILLCELL_X32 FILLER_68_1639 ();
 FILLCELL_X32 FILLER_68_1671 ();
 FILLCELL_X32 FILLER_68_1703 ();
 FILLCELL_X32 FILLER_68_1735 ();
 FILLCELL_X16 FILLER_68_1767 ();
 FILLCELL_X8 FILLER_68_1783 ();
 FILLCELL_X4 FILLER_68_1791 ();
 FILLCELL_X2 FILLER_68_1795 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X16 FILLER_69_801 ();
 FILLCELL_X4 FILLER_69_817 ();
 FILLCELL_X1 FILLER_69_821 ();
 FILLCELL_X32 FILLER_69_829 ();
 FILLCELL_X32 FILLER_69_861 ();
 FILLCELL_X32 FILLER_69_893 ();
 FILLCELL_X32 FILLER_69_925 ();
 FILLCELL_X32 FILLER_69_957 ();
 FILLCELL_X32 FILLER_69_989 ();
 FILLCELL_X32 FILLER_69_1021 ();
 FILLCELL_X32 FILLER_69_1053 ();
 FILLCELL_X32 FILLER_69_1085 ();
 FILLCELL_X32 FILLER_69_1117 ();
 FILLCELL_X32 FILLER_69_1149 ();
 FILLCELL_X32 FILLER_69_1181 ();
 FILLCELL_X32 FILLER_69_1213 ();
 FILLCELL_X16 FILLER_69_1245 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X32 FILLER_69_1584 ();
 FILLCELL_X32 FILLER_69_1616 ();
 FILLCELL_X32 FILLER_69_1648 ();
 FILLCELL_X32 FILLER_69_1680 ();
 FILLCELL_X32 FILLER_69_1712 ();
 FILLCELL_X32 FILLER_69_1744 ();
 FILLCELL_X16 FILLER_69_1776 ();
 FILLCELL_X4 FILLER_69_1792 ();
 FILLCELL_X1 FILLER_69_1796 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X32 FILLER_70_1592 ();
 FILLCELL_X32 FILLER_70_1624 ();
 FILLCELL_X32 FILLER_70_1656 ();
 FILLCELL_X32 FILLER_70_1688 ();
 FILLCELL_X32 FILLER_70_1720 ();
 FILLCELL_X32 FILLER_70_1752 ();
 FILLCELL_X8 FILLER_70_1784 ();
 FILLCELL_X4 FILLER_70_1792 ();
 FILLCELL_X1 FILLER_70_1796 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1584 ();
 FILLCELL_X32 FILLER_71_1616 ();
 FILLCELL_X32 FILLER_71_1648 ();
 FILLCELL_X32 FILLER_71_1680 ();
 FILLCELL_X32 FILLER_71_1712 ();
 FILLCELL_X32 FILLER_71_1744 ();
 FILLCELL_X16 FILLER_71_1776 ();
 FILLCELL_X4 FILLER_71_1792 ();
 FILLCELL_X1 FILLER_71_1796 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X32 FILLER_72_1592 ();
 FILLCELL_X32 FILLER_72_1624 ();
 FILLCELL_X32 FILLER_72_1656 ();
 FILLCELL_X32 FILLER_72_1688 ();
 FILLCELL_X32 FILLER_72_1720 ();
 FILLCELL_X32 FILLER_72_1752 ();
 FILLCELL_X8 FILLER_72_1784 ();
 FILLCELL_X4 FILLER_72_1792 ();
 FILLCELL_X1 FILLER_72_1796 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X32 FILLER_73_1584 ();
 FILLCELL_X32 FILLER_73_1616 ();
 FILLCELL_X32 FILLER_73_1648 ();
 FILLCELL_X32 FILLER_73_1680 ();
 FILLCELL_X32 FILLER_73_1712 ();
 FILLCELL_X32 FILLER_73_1744 ();
 FILLCELL_X16 FILLER_73_1776 ();
 FILLCELL_X4 FILLER_73_1792 ();
 FILLCELL_X1 FILLER_73_1796 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X32 FILLER_74_1592 ();
 FILLCELL_X32 FILLER_74_1624 ();
 FILLCELL_X32 FILLER_74_1656 ();
 FILLCELL_X32 FILLER_74_1688 ();
 FILLCELL_X32 FILLER_74_1720 ();
 FILLCELL_X32 FILLER_74_1752 ();
 FILLCELL_X8 FILLER_74_1784 ();
 FILLCELL_X4 FILLER_74_1792 ();
 FILLCELL_X1 FILLER_74_1796 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X16 FILLER_75_865 ();
 FILLCELL_X8 FILLER_75_881 ();
 FILLCELL_X2 FILLER_75_889 ();
 FILLCELL_X1 FILLER_75_891 ();
 FILLCELL_X32 FILLER_75_902 ();
 FILLCELL_X32 FILLER_75_934 ();
 FILLCELL_X32 FILLER_75_966 ();
 FILLCELL_X32 FILLER_75_998 ();
 FILLCELL_X32 FILLER_75_1030 ();
 FILLCELL_X32 FILLER_75_1062 ();
 FILLCELL_X32 FILLER_75_1094 ();
 FILLCELL_X32 FILLER_75_1126 ();
 FILLCELL_X32 FILLER_75_1158 ();
 FILLCELL_X32 FILLER_75_1190 ();
 FILLCELL_X32 FILLER_75_1222 ();
 FILLCELL_X8 FILLER_75_1254 ();
 FILLCELL_X1 FILLER_75_1262 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X32 FILLER_75_1584 ();
 FILLCELL_X32 FILLER_75_1616 ();
 FILLCELL_X32 FILLER_75_1648 ();
 FILLCELL_X32 FILLER_75_1680 ();
 FILLCELL_X32 FILLER_75_1712 ();
 FILLCELL_X32 FILLER_75_1744 ();
 FILLCELL_X16 FILLER_75_1776 ();
 FILLCELL_X4 FILLER_75_1792 ();
 FILLCELL_X1 FILLER_75_1796 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X8 FILLER_76_856 ();
 FILLCELL_X4 FILLER_76_864 ();
 FILLCELL_X1 FILLER_76_868 ();
 FILLCELL_X16 FILLER_76_879 ();
 FILLCELL_X1 FILLER_76_895 ();
 FILLCELL_X4 FILLER_76_906 ();
 FILLCELL_X2 FILLER_76_910 ();
 FILLCELL_X1 FILLER_76_912 ();
 FILLCELL_X32 FILLER_76_923 ();
 FILLCELL_X32 FILLER_76_955 ();
 FILLCELL_X32 FILLER_76_987 ();
 FILLCELL_X32 FILLER_76_1019 ();
 FILLCELL_X32 FILLER_76_1051 ();
 FILLCELL_X32 FILLER_76_1083 ();
 FILLCELL_X32 FILLER_76_1115 ();
 FILLCELL_X32 FILLER_76_1147 ();
 FILLCELL_X32 FILLER_76_1179 ();
 FILLCELL_X32 FILLER_76_1211 ();
 FILLCELL_X32 FILLER_76_1243 ();
 FILLCELL_X32 FILLER_76_1275 ();
 FILLCELL_X32 FILLER_76_1307 ();
 FILLCELL_X32 FILLER_76_1339 ();
 FILLCELL_X32 FILLER_76_1371 ();
 FILLCELL_X32 FILLER_76_1403 ();
 FILLCELL_X32 FILLER_76_1435 ();
 FILLCELL_X32 FILLER_76_1467 ();
 FILLCELL_X32 FILLER_76_1499 ();
 FILLCELL_X32 FILLER_76_1531 ();
 FILLCELL_X32 FILLER_76_1563 ();
 FILLCELL_X32 FILLER_76_1595 ();
 FILLCELL_X32 FILLER_76_1627 ();
 FILLCELL_X32 FILLER_76_1659 ();
 FILLCELL_X32 FILLER_76_1691 ();
 FILLCELL_X32 FILLER_76_1723 ();
 FILLCELL_X32 FILLER_76_1755 ();
 FILLCELL_X8 FILLER_76_1787 ();
 FILLCELL_X2 FILLER_76_1795 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X4 FILLER_77_865 ();
 FILLCELL_X1 FILLER_77_869 ();
 FILLCELL_X32 FILLER_77_880 ();
 FILLCELL_X4 FILLER_77_912 ();
 FILLCELL_X2 FILLER_77_916 ();
 FILLCELL_X1 FILLER_77_918 ();
 FILLCELL_X1 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_935 ();
 FILLCELL_X32 FILLER_77_967 ();
 FILLCELL_X32 FILLER_77_999 ();
 FILLCELL_X32 FILLER_77_1031 ();
 FILLCELL_X32 FILLER_77_1063 ();
 FILLCELL_X32 FILLER_77_1095 ();
 FILLCELL_X32 FILLER_77_1127 ();
 FILLCELL_X32 FILLER_77_1159 ();
 FILLCELL_X32 FILLER_77_1191 ();
 FILLCELL_X32 FILLER_77_1223 ();
 FILLCELL_X8 FILLER_77_1255 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X32 FILLER_77_1584 ();
 FILLCELL_X32 FILLER_77_1616 ();
 FILLCELL_X32 FILLER_77_1648 ();
 FILLCELL_X32 FILLER_77_1680 ();
 FILLCELL_X32 FILLER_77_1712 ();
 FILLCELL_X32 FILLER_77_1744 ();
 FILLCELL_X16 FILLER_77_1776 ();
 FILLCELL_X4 FILLER_77_1792 ();
 FILLCELL_X1 FILLER_77_1796 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X16 FILLER_78_856 ();
 FILLCELL_X2 FILLER_78_872 ();
 FILLCELL_X16 FILLER_78_881 ();
 FILLCELL_X1 FILLER_78_897 ();
 FILLCELL_X32 FILLER_78_905 ();
 FILLCELL_X32 FILLER_78_937 ();
 FILLCELL_X32 FILLER_78_969 ();
 FILLCELL_X32 FILLER_78_1001 ();
 FILLCELL_X32 FILLER_78_1033 ();
 FILLCELL_X32 FILLER_78_1065 ();
 FILLCELL_X32 FILLER_78_1097 ();
 FILLCELL_X32 FILLER_78_1129 ();
 FILLCELL_X32 FILLER_78_1161 ();
 FILLCELL_X32 FILLER_78_1193 ();
 FILLCELL_X32 FILLER_78_1225 ();
 FILLCELL_X32 FILLER_78_1257 ();
 FILLCELL_X32 FILLER_78_1289 ();
 FILLCELL_X32 FILLER_78_1321 ();
 FILLCELL_X32 FILLER_78_1353 ();
 FILLCELL_X32 FILLER_78_1385 ();
 FILLCELL_X32 FILLER_78_1417 ();
 FILLCELL_X32 FILLER_78_1449 ();
 FILLCELL_X32 FILLER_78_1481 ();
 FILLCELL_X32 FILLER_78_1513 ();
 FILLCELL_X32 FILLER_78_1545 ();
 FILLCELL_X32 FILLER_78_1577 ();
 FILLCELL_X32 FILLER_78_1609 ();
 FILLCELL_X32 FILLER_78_1641 ();
 FILLCELL_X32 FILLER_78_1673 ();
 FILLCELL_X32 FILLER_78_1705 ();
 FILLCELL_X32 FILLER_78_1737 ();
 FILLCELL_X16 FILLER_78_1769 ();
 FILLCELL_X8 FILLER_78_1785 ();
 FILLCELL_X4 FILLER_78_1793 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X8 FILLER_79_865 ();
 FILLCELL_X1 FILLER_79_873 ();
 FILLCELL_X1 FILLER_79_884 ();
 FILLCELL_X4 FILLER_79_892 ();
 FILLCELL_X1 FILLER_79_900 ();
 FILLCELL_X4 FILLER_79_914 ();
 FILLCELL_X2 FILLER_79_918 ();
 FILLCELL_X32 FILLER_79_938 ();
 FILLCELL_X32 FILLER_79_970 ();
 FILLCELL_X32 FILLER_79_1002 ();
 FILLCELL_X32 FILLER_79_1034 ();
 FILLCELL_X32 FILLER_79_1066 ();
 FILLCELL_X32 FILLER_79_1098 ();
 FILLCELL_X32 FILLER_79_1130 ();
 FILLCELL_X32 FILLER_79_1162 ();
 FILLCELL_X32 FILLER_79_1194 ();
 FILLCELL_X32 FILLER_79_1226 ();
 FILLCELL_X4 FILLER_79_1258 ();
 FILLCELL_X1 FILLER_79_1262 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X32 FILLER_79_1584 ();
 FILLCELL_X32 FILLER_79_1616 ();
 FILLCELL_X32 FILLER_79_1648 ();
 FILLCELL_X32 FILLER_79_1680 ();
 FILLCELL_X32 FILLER_79_1712 ();
 FILLCELL_X32 FILLER_79_1744 ();
 FILLCELL_X16 FILLER_79_1776 ();
 FILLCELL_X4 FILLER_79_1792 ();
 FILLCELL_X1 FILLER_79_1796 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X16 FILLER_80_856 ();
 FILLCELL_X4 FILLER_80_872 ();
 FILLCELL_X2 FILLER_80_876 ();
 FILLCELL_X8 FILLER_80_885 ();
 FILLCELL_X1 FILLER_80_893 ();
 FILLCELL_X2 FILLER_80_903 ();
 FILLCELL_X8 FILLER_80_909 ();
 FILLCELL_X1 FILLER_80_917 ();
 FILLCELL_X1 FILLER_80_925 ();
 FILLCELL_X32 FILLER_80_942 ();
 FILLCELL_X32 FILLER_80_974 ();
 FILLCELL_X32 FILLER_80_1006 ();
 FILLCELL_X32 FILLER_80_1038 ();
 FILLCELL_X32 FILLER_80_1070 ();
 FILLCELL_X32 FILLER_80_1102 ();
 FILLCELL_X32 FILLER_80_1134 ();
 FILLCELL_X32 FILLER_80_1166 ();
 FILLCELL_X32 FILLER_80_1198 ();
 FILLCELL_X32 FILLER_80_1230 ();
 FILLCELL_X32 FILLER_80_1262 ();
 FILLCELL_X32 FILLER_80_1294 ();
 FILLCELL_X32 FILLER_80_1326 ();
 FILLCELL_X32 FILLER_80_1358 ();
 FILLCELL_X32 FILLER_80_1390 ();
 FILLCELL_X32 FILLER_80_1422 ();
 FILLCELL_X32 FILLER_80_1454 ();
 FILLCELL_X32 FILLER_80_1486 ();
 FILLCELL_X32 FILLER_80_1518 ();
 FILLCELL_X32 FILLER_80_1550 ();
 FILLCELL_X32 FILLER_80_1582 ();
 FILLCELL_X32 FILLER_80_1614 ();
 FILLCELL_X32 FILLER_80_1646 ();
 FILLCELL_X32 FILLER_80_1678 ();
 FILLCELL_X32 FILLER_80_1710 ();
 FILLCELL_X32 FILLER_80_1742 ();
 FILLCELL_X16 FILLER_80_1774 ();
 FILLCELL_X4 FILLER_80_1790 ();
 FILLCELL_X2 FILLER_80_1794 ();
 FILLCELL_X1 FILLER_80_1796 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X16 FILLER_81_897 ();
 FILLCELL_X8 FILLER_81_913 ();
 FILLCELL_X2 FILLER_81_921 ();
 FILLCELL_X1 FILLER_81_923 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X32 FILLER_81_1584 ();
 FILLCELL_X32 FILLER_81_1616 ();
 FILLCELL_X32 FILLER_81_1648 ();
 FILLCELL_X32 FILLER_81_1680 ();
 FILLCELL_X32 FILLER_81_1712 ();
 FILLCELL_X32 FILLER_81_1744 ();
 FILLCELL_X16 FILLER_81_1776 ();
 FILLCELL_X4 FILLER_81_1792 ();
 FILLCELL_X1 FILLER_81_1796 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X32 FILLER_82_1592 ();
 FILLCELL_X32 FILLER_82_1624 ();
 FILLCELL_X32 FILLER_82_1656 ();
 FILLCELL_X32 FILLER_82_1688 ();
 FILLCELL_X32 FILLER_82_1720 ();
 FILLCELL_X32 FILLER_82_1752 ();
 FILLCELL_X8 FILLER_82_1784 ();
 FILLCELL_X4 FILLER_82_1792 ();
 FILLCELL_X1 FILLER_82_1796 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X32 FILLER_83_1584 ();
 FILLCELL_X32 FILLER_83_1616 ();
 FILLCELL_X32 FILLER_83_1648 ();
 FILLCELL_X32 FILLER_83_1680 ();
 FILLCELL_X32 FILLER_83_1712 ();
 FILLCELL_X32 FILLER_83_1744 ();
 FILLCELL_X16 FILLER_83_1776 ();
 FILLCELL_X4 FILLER_83_1792 ();
 FILLCELL_X1 FILLER_83_1796 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X32 FILLER_84_1592 ();
 FILLCELL_X32 FILLER_84_1624 ();
 FILLCELL_X32 FILLER_84_1656 ();
 FILLCELL_X32 FILLER_84_1688 ();
 FILLCELL_X32 FILLER_84_1720 ();
 FILLCELL_X32 FILLER_84_1752 ();
 FILLCELL_X8 FILLER_84_1784 ();
 FILLCELL_X4 FILLER_84_1792 ();
 FILLCELL_X1 FILLER_84_1796 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X32 FILLER_85_1584 ();
 FILLCELL_X32 FILLER_85_1616 ();
 FILLCELL_X32 FILLER_85_1648 ();
 FILLCELL_X32 FILLER_85_1680 ();
 FILLCELL_X32 FILLER_85_1712 ();
 FILLCELL_X32 FILLER_85_1744 ();
 FILLCELL_X16 FILLER_85_1776 ();
 FILLCELL_X4 FILLER_85_1792 ();
 FILLCELL_X1 FILLER_85_1796 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X32 FILLER_86_1592 ();
 FILLCELL_X32 FILLER_86_1624 ();
 FILLCELL_X32 FILLER_86_1656 ();
 FILLCELL_X32 FILLER_86_1688 ();
 FILLCELL_X32 FILLER_86_1720 ();
 FILLCELL_X32 FILLER_86_1752 ();
 FILLCELL_X8 FILLER_86_1784 ();
 FILLCELL_X4 FILLER_86_1792 ();
 FILLCELL_X1 FILLER_86_1796 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X32 FILLER_87_1584 ();
 FILLCELL_X32 FILLER_87_1616 ();
 FILLCELL_X32 FILLER_87_1648 ();
 FILLCELL_X32 FILLER_87_1680 ();
 FILLCELL_X32 FILLER_87_1712 ();
 FILLCELL_X32 FILLER_87_1744 ();
 FILLCELL_X16 FILLER_87_1776 ();
 FILLCELL_X4 FILLER_87_1792 ();
 FILLCELL_X1 FILLER_87_1796 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X32 FILLER_88_1592 ();
 FILLCELL_X32 FILLER_88_1624 ();
 FILLCELL_X32 FILLER_88_1656 ();
 FILLCELL_X32 FILLER_88_1688 ();
 FILLCELL_X32 FILLER_88_1720 ();
 FILLCELL_X32 FILLER_88_1752 ();
 FILLCELL_X8 FILLER_88_1784 ();
 FILLCELL_X4 FILLER_88_1792 ();
 FILLCELL_X1 FILLER_88_1796 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X32 FILLER_89_1584 ();
 FILLCELL_X32 FILLER_89_1616 ();
 FILLCELL_X32 FILLER_89_1648 ();
 FILLCELL_X32 FILLER_89_1680 ();
 FILLCELL_X32 FILLER_89_1712 ();
 FILLCELL_X32 FILLER_89_1744 ();
 FILLCELL_X16 FILLER_89_1776 ();
 FILLCELL_X4 FILLER_89_1792 ();
 FILLCELL_X1 FILLER_89_1796 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X32 FILLER_90_1592 ();
 FILLCELL_X32 FILLER_90_1624 ();
 FILLCELL_X32 FILLER_90_1656 ();
 FILLCELL_X32 FILLER_90_1688 ();
 FILLCELL_X32 FILLER_90_1720 ();
 FILLCELL_X32 FILLER_90_1752 ();
 FILLCELL_X8 FILLER_90_1784 ();
 FILLCELL_X4 FILLER_90_1792 ();
 FILLCELL_X1 FILLER_90_1796 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X32 FILLER_91_1584 ();
 FILLCELL_X32 FILLER_91_1616 ();
 FILLCELL_X32 FILLER_91_1648 ();
 FILLCELL_X32 FILLER_91_1680 ();
 FILLCELL_X32 FILLER_91_1712 ();
 FILLCELL_X32 FILLER_91_1744 ();
 FILLCELL_X16 FILLER_91_1776 ();
 FILLCELL_X4 FILLER_91_1792 ();
 FILLCELL_X1 FILLER_91_1796 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X32 FILLER_92_1592 ();
 FILLCELL_X32 FILLER_92_1624 ();
 FILLCELL_X32 FILLER_92_1656 ();
 FILLCELL_X32 FILLER_92_1688 ();
 FILLCELL_X32 FILLER_92_1720 ();
 FILLCELL_X32 FILLER_92_1752 ();
 FILLCELL_X8 FILLER_92_1784 ();
 FILLCELL_X4 FILLER_92_1792 ();
 FILLCELL_X1 FILLER_92_1796 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X32 FILLER_93_1584 ();
 FILLCELL_X32 FILLER_93_1616 ();
 FILLCELL_X32 FILLER_93_1648 ();
 FILLCELL_X32 FILLER_93_1680 ();
 FILLCELL_X32 FILLER_93_1712 ();
 FILLCELL_X32 FILLER_93_1744 ();
 FILLCELL_X16 FILLER_93_1776 ();
 FILLCELL_X4 FILLER_93_1792 ();
 FILLCELL_X1 FILLER_93_1796 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X32 FILLER_94_1592 ();
 FILLCELL_X32 FILLER_94_1624 ();
 FILLCELL_X32 FILLER_94_1656 ();
 FILLCELL_X32 FILLER_94_1688 ();
 FILLCELL_X32 FILLER_94_1720 ();
 FILLCELL_X32 FILLER_94_1752 ();
 FILLCELL_X8 FILLER_94_1784 ();
 FILLCELL_X4 FILLER_94_1792 ();
 FILLCELL_X1 FILLER_94_1796 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X32 FILLER_95_961 ();
 FILLCELL_X32 FILLER_95_993 ();
 FILLCELL_X32 FILLER_95_1025 ();
 FILLCELL_X32 FILLER_95_1057 ();
 FILLCELL_X32 FILLER_95_1089 ();
 FILLCELL_X32 FILLER_95_1121 ();
 FILLCELL_X32 FILLER_95_1153 ();
 FILLCELL_X32 FILLER_95_1185 ();
 FILLCELL_X32 FILLER_95_1217 ();
 FILLCELL_X8 FILLER_95_1249 ();
 FILLCELL_X4 FILLER_95_1257 ();
 FILLCELL_X2 FILLER_95_1261 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X32 FILLER_95_1584 ();
 FILLCELL_X32 FILLER_95_1616 ();
 FILLCELL_X32 FILLER_95_1648 ();
 FILLCELL_X32 FILLER_95_1680 ();
 FILLCELL_X32 FILLER_95_1712 ();
 FILLCELL_X32 FILLER_95_1744 ();
 FILLCELL_X16 FILLER_95_1776 ();
 FILLCELL_X4 FILLER_95_1792 ();
 FILLCELL_X1 FILLER_95_1796 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X32 FILLER_96_1592 ();
 FILLCELL_X32 FILLER_96_1624 ();
 FILLCELL_X32 FILLER_96_1656 ();
 FILLCELL_X32 FILLER_96_1688 ();
 FILLCELL_X32 FILLER_96_1720 ();
 FILLCELL_X32 FILLER_96_1752 ();
 FILLCELL_X8 FILLER_96_1784 ();
 FILLCELL_X4 FILLER_96_1792 ();
 FILLCELL_X1 FILLER_96_1796 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X32 FILLER_97_961 ();
 FILLCELL_X32 FILLER_97_993 ();
 FILLCELL_X32 FILLER_97_1025 ();
 FILLCELL_X32 FILLER_97_1057 ();
 FILLCELL_X32 FILLER_97_1089 ();
 FILLCELL_X32 FILLER_97_1121 ();
 FILLCELL_X32 FILLER_97_1153 ();
 FILLCELL_X32 FILLER_97_1185 ();
 FILLCELL_X32 FILLER_97_1217 ();
 FILLCELL_X8 FILLER_97_1249 ();
 FILLCELL_X4 FILLER_97_1257 ();
 FILLCELL_X2 FILLER_97_1261 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X32 FILLER_97_1584 ();
 FILLCELL_X32 FILLER_97_1616 ();
 FILLCELL_X32 FILLER_97_1648 ();
 FILLCELL_X32 FILLER_97_1680 ();
 FILLCELL_X32 FILLER_97_1712 ();
 FILLCELL_X32 FILLER_97_1744 ();
 FILLCELL_X16 FILLER_97_1776 ();
 FILLCELL_X4 FILLER_97_1792 ();
 FILLCELL_X1 FILLER_97_1796 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X32 FILLER_98_1304 ();
 FILLCELL_X32 FILLER_98_1336 ();
 FILLCELL_X32 FILLER_98_1368 ();
 FILLCELL_X32 FILLER_98_1400 ();
 FILLCELL_X32 FILLER_98_1432 ();
 FILLCELL_X32 FILLER_98_1464 ();
 FILLCELL_X32 FILLER_98_1496 ();
 FILLCELL_X32 FILLER_98_1528 ();
 FILLCELL_X32 FILLER_98_1560 ();
 FILLCELL_X32 FILLER_98_1592 ();
 FILLCELL_X32 FILLER_98_1624 ();
 FILLCELL_X32 FILLER_98_1656 ();
 FILLCELL_X32 FILLER_98_1688 ();
 FILLCELL_X32 FILLER_98_1720 ();
 FILLCELL_X32 FILLER_98_1752 ();
 FILLCELL_X8 FILLER_98_1784 ();
 FILLCELL_X4 FILLER_98_1792 ();
 FILLCELL_X1 FILLER_98_1796 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X32 FILLER_99_1584 ();
 FILLCELL_X32 FILLER_99_1616 ();
 FILLCELL_X32 FILLER_99_1648 ();
 FILLCELL_X32 FILLER_99_1680 ();
 FILLCELL_X32 FILLER_99_1712 ();
 FILLCELL_X32 FILLER_99_1744 ();
 FILLCELL_X16 FILLER_99_1776 ();
 FILLCELL_X4 FILLER_99_1792 ();
 FILLCELL_X1 FILLER_99_1796 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X32 FILLER_100_952 ();
 FILLCELL_X32 FILLER_100_984 ();
 FILLCELL_X32 FILLER_100_1016 ();
 FILLCELL_X32 FILLER_100_1048 ();
 FILLCELL_X32 FILLER_100_1080 ();
 FILLCELL_X32 FILLER_100_1112 ();
 FILLCELL_X32 FILLER_100_1144 ();
 FILLCELL_X32 FILLER_100_1176 ();
 FILLCELL_X32 FILLER_100_1208 ();
 FILLCELL_X32 FILLER_100_1240 ();
 FILLCELL_X32 FILLER_100_1272 ();
 FILLCELL_X32 FILLER_100_1304 ();
 FILLCELL_X32 FILLER_100_1336 ();
 FILLCELL_X32 FILLER_100_1368 ();
 FILLCELL_X32 FILLER_100_1400 ();
 FILLCELL_X32 FILLER_100_1432 ();
 FILLCELL_X32 FILLER_100_1464 ();
 FILLCELL_X32 FILLER_100_1496 ();
 FILLCELL_X32 FILLER_100_1528 ();
 FILLCELL_X32 FILLER_100_1560 ();
 FILLCELL_X32 FILLER_100_1592 ();
 FILLCELL_X32 FILLER_100_1624 ();
 FILLCELL_X32 FILLER_100_1656 ();
 FILLCELL_X32 FILLER_100_1688 ();
 FILLCELL_X32 FILLER_100_1720 ();
 FILLCELL_X32 FILLER_100_1752 ();
 FILLCELL_X8 FILLER_100_1784 ();
 FILLCELL_X4 FILLER_100_1792 ();
 FILLCELL_X1 FILLER_100_1796 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X32 FILLER_101_1584 ();
 FILLCELL_X32 FILLER_101_1616 ();
 FILLCELL_X32 FILLER_101_1648 ();
 FILLCELL_X32 FILLER_101_1680 ();
 FILLCELL_X32 FILLER_101_1712 ();
 FILLCELL_X32 FILLER_101_1744 ();
 FILLCELL_X16 FILLER_101_1776 ();
 FILLCELL_X4 FILLER_101_1792 ();
 FILLCELL_X1 FILLER_101_1796 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X32 FILLER_102_1304 ();
 FILLCELL_X32 FILLER_102_1336 ();
 FILLCELL_X32 FILLER_102_1368 ();
 FILLCELL_X32 FILLER_102_1400 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X32 FILLER_102_1496 ();
 FILLCELL_X32 FILLER_102_1528 ();
 FILLCELL_X32 FILLER_102_1560 ();
 FILLCELL_X32 FILLER_102_1592 ();
 FILLCELL_X32 FILLER_102_1624 ();
 FILLCELL_X32 FILLER_102_1656 ();
 FILLCELL_X32 FILLER_102_1688 ();
 FILLCELL_X32 FILLER_102_1720 ();
 FILLCELL_X32 FILLER_102_1752 ();
 FILLCELL_X8 FILLER_102_1784 ();
 FILLCELL_X4 FILLER_102_1792 ();
 FILLCELL_X1 FILLER_102_1796 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X32 FILLER_103_1584 ();
 FILLCELL_X32 FILLER_103_1616 ();
 FILLCELL_X32 FILLER_103_1648 ();
 FILLCELL_X32 FILLER_103_1680 ();
 FILLCELL_X32 FILLER_103_1712 ();
 FILLCELL_X32 FILLER_103_1744 ();
 FILLCELL_X16 FILLER_103_1776 ();
 FILLCELL_X4 FILLER_103_1792 ();
 FILLCELL_X1 FILLER_103_1796 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X32 FILLER_104_1304 ();
 FILLCELL_X32 FILLER_104_1336 ();
 FILLCELL_X32 FILLER_104_1368 ();
 FILLCELL_X32 FILLER_104_1400 ();
 FILLCELL_X32 FILLER_104_1432 ();
 FILLCELL_X32 FILLER_104_1464 ();
 FILLCELL_X32 FILLER_104_1496 ();
 FILLCELL_X32 FILLER_104_1528 ();
 FILLCELL_X32 FILLER_104_1560 ();
 FILLCELL_X32 FILLER_104_1592 ();
 FILLCELL_X32 FILLER_104_1624 ();
 FILLCELL_X32 FILLER_104_1656 ();
 FILLCELL_X32 FILLER_104_1688 ();
 FILLCELL_X32 FILLER_104_1720 ();
 FILLCELL_X32 FILLER_104_1752 ();
 FILLCELL_X8 FILLER_104_1784 ();
 FILLCELL_X4 FILLER_104_1792 ();
 FILLCELL_X1 FILLER_104_1796 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X32 FILLER_105_961 ();
 FILLCELL_X32 FILLER_105_993 ();
 FILLCELL_X32 FILLER_105_1025 ();
 FILLCELL_X32 FILLER_105_1057 ();
 FILLCELL_X32 FILLER_105_1089 ();
 FILLCELL_X32 FILLER_105_1121 ();
 FILLCELL_X32 FILLER_105_1153 ();
 FILLCELL_X32 FILLER_105_1185 ();
 FILLCELL_X32 FILLER_105_1217 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X32 FILLER_105_1584 ();
 FILLCELL_X32 FILLER_105_1616 ();
 FILLCELL_X32 FILLER_105_1648 ();
 FILLCELL_X32 FILLER_105_1680 ();
 FILLCELL_X32 FILLER_105_1712 ();
 FILLCELL_X32 FILLER_105_1744 ();
 FILLCELL_X16 FILLER_105_1776 ();
 FILLCELL_X4 FILLER_105_1792 ();
 FILLCELL_X1 FILLER_105_1796 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X32 FILLER_106_1304 ();
 FILLCELL_X32 FILLER_106_1336 ();
 FILLCELL_X32 FILLER_106_1368 ();
 FILLCELL_X32 FILLER_106_1400 ();
 FILLCELL_X32 FILLER_106_1432 ();
 FILLCELL_X32 FILLER_106_1464 ();
 FILLCELL_X32 FILLER_106_1496 ();
 FILLCELL_X32 FILLER_106_1528 ();
 FILLCELL_X32 FILLER_106_1560 ();
 FILLCELL_X32 FILLER_106_1592 ();
 FILLCELL_X32 FILLER_106_1624 ();
 FILLCELL_X32 FILLER_106_1656 ();
 FILLCELL_X32 FILLER_106_1688 ();
 FILLCELL_X32 FILLER_106_1720 ();
 FILLCELL_X32 FILLER_106_1752 ();
 FILLCELL_X8 FILLER_106_1784 ();
 FILLCELL_X4 FILLER_106_1792 ();
 FILLCELL_X1 FILLER_106_1796 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X32 FILLER_107_961 ();
 FILLCELL_X32 FILLER_107_993 ();
 FILLCELL_X32 FILLER_107_1025 ();
 FILLCELL_X32 FILLER_107_1057 ();
 FILLCELL_X32 FILLER_107_1089 ();
 FILLCELL_X32 FILLER_107_1121 ();
 FILLCELL_X32 FILLER_107_1153 ();
 FILLCELL_X32 FILLER_107_1185 ();
 FILLCELL_X32 FILLER_107_1217 ();
 FILLCELL_X8 FILLER_107_1249 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X32 FILLER_107_1584 ();
 FILLCELL_X32 FILLER_107_1616 ();
 FILLCELL_X32 FILLER_107_1648 ();
 FILLCELL_X32 FILLER_107_1680 ();
 FILLCELL_X32 FILLER_107_1712 ();
 FILLCELL_X32 FILLER_107_1744 ();
 FILLCELL_X16 FILLER_107_1776 ();
 FILLCELL_X4 FILLER_107_1792 ();
 FILLCELL_X1 FILLER_107_1796 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X32 FILLER_108_856 ();
 FILLCELL_X32 FILLER_108_888 ();
 FILLCELL_X32 FILLER_108_920 ();
 FILLCELL_X32 FILLER_108_952 ();
 FILLCELL_X32 FILLER_108_984 ();
 FILLCELL_X32 FILLER_108_1016 ();
 FILLCELL_X32 FILLER_108_1048 ();
 FILLCELL_X32 FILLER_108_1080 ();
 FILLCELL_X32 FILLER_108_1112 ();
 FILLCELL_X32 FILLER_108_1144 ();
 FILLCELL_X32 FILLER_108_1176 ();
 FILLCELL_X32 FILLER_108_1208 ();
 FILLCELL_X32 FILLER_108_1240 ();
 FILLCELL_X32 FILLER_108_1272 ();
 FILLCELL_X32 FILLER_108_1304 ();
 FILLCELL_X32 FILLER_108_1336 ();
 FILLCELL_X32 FILLER_108_1368 ();
 FILLCELL_X32 FILLER_108_1400 ();
 FILLCELL_X32 FILLER_108_1432 ();
 FILLCELL_X32 FILLER_108_1464 ();
 FILLCELL_X32 FILLER_108_1496 ();
 FILLCELL_X32 FILLER_108_1528 ();
 FILLCELL_X32 FILLER_108_1560 ();
 FILLCELL_X32 FILLER_108_1592 ();
 FILLCELL_X32 FILLER_108_1624 ();
 FILLCELL_X32 FILLER_108_1656 ();
 FILLCELL_X32 FILLER_108_1688 ();
 FILLCELL_X32 FILLER_108_1720 ();
 FILLCELL_X32 FILLER_108_1752 ();
 FILLCELL_X8 FILLER_108_1784 ();
 FILLCELL_X4 FILLER_108_1792 ();
 FILLCELL_X1 FILLER_108_1796 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X32 FILLER_109_1584 ();
 FILLCELL_X32 FILLER_109_1616 ();
 FILLCELL_X32 FILLER_109_1648 ();
 FILLCELL_X32 FILLER_109_1680 ();
 FILLCELL_X16 FILLER_109_1712 ();
 FILLCELL_X8 FILLER_109_1728 ();
 FILLCELL_X4 FILLER_109_1736 ();
 FILLCELL_X4 FILLER_109_1749 ();
 FILLCELL_X2 FILLER_109_1753 ();
 FILLCELL_X2 FILLER_109_1757 ();
 FILLCELL_X1 FILLER_109_1759 ();
 FILLCELL_X16 FILLER_109_1769 ();
 FILLCELL_X8 FILLER_109_1785 ();
 FILLCELL_X4 FILLER_109_1793 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X32 FILLER_110_952 ();
 FILLCELL_X32 FILLER_110_984 ();
 FILLCELL_X32 FILLER_110_1016 ();
 FILLCELL_X32 FILLER_110_1048 ();
 FILLCELL_X32 FILLER_110_1080 ();
 FILLCELL_X32 FILLER_110_1112 ();
 FILLCELL_X32 FILLER_110_1144 ();
 FILLCELL_X32 FILLER_110_1176 ();
 FILLCELL_X32 FILLER_110_1208 ();
 FILLCELL_X32 FILLER_110_1240 ();
 FILLCELL_X32 FILLER_110_1272 ();
 FILLCELL_X32 FILLER_110_1304 ();
 FILLCELL_X32 FILLER_110_1336 ();
 FILLCELL_X32 FILLER_110_1368 ();
 FILLCELL_X32 FILLER_110_1400 ();
 FILLCELL_X32 FILLER_110_1432 ();
 FILLCELL_X32 FILLER_110_1464 ();
 FILLCELL_X32 FILLER_110_1496 ();
 FILLCELL_X32 FILLER_110_1528 ();
 FILLCELL_X32 FILLER_110_1560 ();
 FILLCELL_X32 FILLER_110_1592 ();
 FILLCELL_X32 FILLER_110_1624 ();
 FILLCELL_X32 FILLER_110_1656 ();
 FILLCELL_X32 FILLER_110_1688 ();
 FILLCELL_X8 FILLER_110_1720 ();
 FILLCELL_X4 FILLER_110_1728 ();
 FILLCELL_X1 FILLER_110_1732 ();
 FILLCELL_X1 FILLER_110_1753 ();
 FILLCELL_X8 FILLER_110_1767 ();
 FILLCELL_X2 FILLER_110_1775 ();
 FILLCELL_X1 FILLER_110_1796 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X32 FILLER_111_961 ();
 FILLCELL_X32 FILLER_111_993 ();
 FILLCELL_X32 FILLER_111_1025 ();
 FILLCELL_X32 FILLER_111_1057 ();
 FILLCELL_X32 FILLER_111_1089 ();
 FILLCELL_X32 FILLER_111_1121 ();
 FILLCELL_X32 FILLER_111_1153 ();
 FILLCELL_X32 FILLER_111_1185 ();
 FILLCELL_X32 FILLER_111_1217 ();
 FILLCELL_X8 FILLER_111_1249 ();
 FILLCELL_X4 FILLER_111_1257 ();
 FILLCELL_X2 FILLER_111_1261 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X32 FILLER_111_1584 ();
 FILLCELL_X32 FILLER_111_1616 ();
 FILLCELL_X32 FILLER_111_1648 ();
 FILLCELL_X32 FILLER_111_1680 ();
 FILLCELL_X16 FILLER_111_1712 ();
 FILLCELL_X8 FILLER_111_1728 ();
 FILLCELL_X2 FILLER_111_1736 ();
 FILLCELL_X4 FILLER_111_1742 ();
 FILLCELL_X16 FILLER_111_1750 ();
 FILLCELL_X2 FILLER_111_1766 ();
 FILLCELL_X1 FILLER_111_1768 ();
 FILLCELL_X8 FILLER_111_1772 ();
 FILLCELL_X4 FILLER_111_1780 ();
 FILLCELL_X2 FILLER_111_1788 ();
 FILLCELL_X1 FILLER_111_1790 ();
 FILLCELL_X32 FILLER_112_20 ();
 FILLCELL_X32 FILLER_112_52 ();
 FILLCELL_X32 FILLER_112_84 ();
 FILLCELL_X32 FILLER_112_116 ();
 FILLCELL_X32 FILLER_112_148 ();
 FILLCELL_X32 FILLER_112_180 ();
 FILLCELL_X32 FILLER_112_212 ();
 FILLCELL_X32 FILLER_112_244 ();
 FILLCELL_X32 FILLER_112_276 ();
 FILLCELL_X32 FILLER_112_308 ();
 FILLCELL_X32 FILLER_112_340 ();
 FILLCELL_X32 FILLER_112_372 ();
 FILLCELL_X32 FILLER_112_404 ();
 FILLCELL_X32 FILLER_112_436 ();
 FILLCELL_X32 FILLER_112_468 ();
 FILLCELL_X32 FILLER_112_500 ();
 FILLCELL_X32 FILLER_112_532 ();
 FILLCELL_X32 FILLER_112_564 ();
 FILLCELL_X32 FILLER_112_596 ();
 FILLCELL_X2 FILLER_112_628 ();
 FILLCELL_X1 FILLER_112_630 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X32 FILLER_112_952 ();
 FILLCELL_X32 FILLER_112_984 ();
 FILLCELL_X32 FILLER_112_1016 ();
 FILLCELL_X32 FILLER_112_1048 ();
 FILLCELL_X32 FILLER_112_1080 ();
 FILLCELL_X32 FILLER_112_1112 ();
 FILLCELL_X32 FILLER_112_1144 ();
 FILLCELL_X32 FILLER_112_1176 ();
 FILLCELL_X32 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_112_1240 ();
 FILLCELL_X32 FILLER_112_1272 ();
 FILLCELL_X32 FILLER_112_1304 ();
 FILLCELL_X32 FILLER_112_1336 ();
 FILLCELL_X32 FILLER_112_1368 ();
 FILLCELL_X32 FILLER_112_1400 ();
 FILLCELL_X32 FILLER_112_1432 ();
 FILLCELL_X32 FILLER_112_1464 ();
 FILLCELL_X32 FILLER_112_1496 ();
 FILLCELL_X32 FILLER_112_1528 ();
 FILLCELL_X32 FILLER_112_1560 ();
 FILLCELL_X32 FILLER_112_1592 ();
 FILLCELL_X32 FILLER_112_1624 ();
 FILLCELL_X32 FILLER_112_1656 ();
 FILLCELL_X32 FILLER_112_1688 ();
 FILLCELL_X16 FILLER_112_1720 ();
 FILLCELL_X2 FILLER_112_1736 ();
 FILLCELL_X1 FILLER_112_1738 ();
 FILLCELL_X8 FILLER_112_1742 ();
 FILLCELL_X4 FILLER_112_1750 ();
 FILLCELL_X16 FILLER_112_1760 ();
 FILLCELL_X8 FILLER_112_1776 ();
 FILLCELL_X4 FILLER_112_1784 ();
 FILLCELL_X2 FILLER_112_1788 ();
 FILLCELL_X1 FILLER_112_1790 ();
 FILLCELL_X1 FILLER_113_4 ();
 FILLCELL_X32 FILLER_113_23 ();
 FILLCELL_X32 FILLER_113_55 ();
 FILLCELL_X32 FILLER_113_87 ();
 FILLCELL_X32 FILLER_113_119 ();
 FILLCELL_X32 FILLER_113_151 ();
 FILLCELL_X32 FILLER_113_183 ();
 FILLCELL_X32 FILLER_113_215 ();
 FILLCELL_X32 FILLER_113_247 ();
 FILLCELL_X32 FILLER_113_279 ();
 FILLCELL_X32 FILLER_113_311 ();
 FILLCELL_X32 FILLER_113_343 ();
 FILLCELL_X32 FILLER_113_375 ();
 FILLCELL_X32 FILLER_113_407 ();
 FILLCELL_X32 FILLER_113_439 ();
 FILLCELL_X32 FILLER_113_471 ();
 FILLCELL_X32 FILLER_113_503 ();
 FILLCELL_X32 FILLER_113_535 ();
 FILLCELL_X32 FILLER_113_567 ();
 FILLCELL_X32 FILLER_113_599 ();
 FILLCELL_X32 FILLER_113_631 ();
 FILLCELL_X32 FILLER_113_663 ();
 FILLCELL_X32 FILLER_113_695 ();
 FILLCELL_X32 FILLER_113_727 ();
 FILLCELL_X32 FILLER_113_759 ();
 FILLCELL_X32 FILLER_113_791 ();
 FILLCELL_X32 FILLER_113_823 ();
 FILLCELL_X32 FILLER_113_855 ();
 FILLCELL_X32 FILLER_113_887 ();
 FILLCELL_X32 FILLER_113_919 ();
 FILLCELL_X32 FILLER_113_951 ();
 FILLCELL_X32 FILLER_113_983 ();
 FILLCELL_X32 FILLER_113_1015 ();
 FILLCELL_X32 FILLER_113_1047 ();
 FILLCELL_X32 FILLER_113_1079 ();
 FILLCELL_X32 FILLER_113_1111 ();
 FILLCELL_X32 FILLER_113_1143 ();
 FILLCELL_X32 FILLER_113_1175 ();
 FILLCELL_X32 FILLER_113_1207 ();
 FILLCELL_X16 FILLER_113_1239 ();
 FILLCELL_X8 FILLER_113_1255 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X32 FILLER_113_1552 ();
 FILLCELL_X32 FILLER_113_1584 ();
 FILLCELL_X32 FILLER_113_1616 ();
 FILLCELL_X32 FILLER_113_1648 ();
 FILLCELL_X32 FILLER_113_1680 ();
 FILLCELL_X16 FILLER_113_1712 ();
 FILLCELL_X4 FILLER_113_1728 ();
 FILLCELL_X4 FILLER_113_1750 ();
 FILLCELL_X1 FILLER_113_1754 ();
 FILLCELL_X4 FILLER_113_1766 ();
 FILLCELL_X2 FILLER_113_1770 ();
 FILLCELL_X1 FILLER_113_1772 ();
 FILLCELL_X1 FILLER_113_1793 ();
 FILLCELL_X8 FILLER_114_1 ();
 FILLCELL_X4 FILLER_114_9 ();
 FILLCELL_X2 FILLER_114_13 ();
 FILLCELL_X1 FILLER_114_15 ();
 FILLCELL_X2 FILLER_114_19 ();
 FILLCELL_X1 FILLER_114_21 ();
 FILLCELL_X2 FILLER_114_28 ();
 FILLCELL_X1 FILLER_114_30 ();
 FILLCELL_X1 FILLER_114_50 ();
 FILLCELL_X32 FILLER_114_53 ();
 FILLCELL_X32 FILLER_114_85 ();
 FILLCELL_X32 FILLER_114_117 ();
 FILLCELL_X32 FILLER_114_149 ();
 FILLCELL_X32 FILLER_114_181 ();
 FILLCELL_X32 FILLER_114_213 ();
 FILLCELL_X32 FILLER_114_245 ();
 FILLCELL_X32 FILLER_114_277 ();
 FILLCELL_X32 FILLER_114_309 ();
 FILLCELL_X32 FILLER_114_341 ();
 FILLCELL_X32 FILLER_114_373 ();
 FILLCELL_X32 FILLER_114_405 ();
 FILLCELL_X32 FILLER_114_437 ();
 FILLCELL_X32 FILLER_114_469 ();
 FILLCELL_X32 FILLER_114_501 ();
 FILLCELL_X32 FILLER_114_533 ();
 FILLCELL_X32 FILLER_114_565 ();
 FILLCELL_X32 FILLER_114_597 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X32 FILLER_114_952 ();
 FILLCELL_X32 FILLER_114_984 ();
 FILLCELL_X32 FILLER_114_1016 ();
 FILLCELL_X32 FILLER_114_1048 ();
 FILLCELL_X32 FILLER_114_1080 ();
 FILLCELL_X32 FILLER_114_1112 ();
 FILLCELL_X32 FILLER_114_1144 ();
 FILLCELL_X32 FILLER_114_1176 ();
 FILLCELL_X32 FILLER_114_1208 ();
 FILLCELL_X32 FILLER_114_1240 ();
 FILLCELL_X32 FILLER_114_1272 ();
 FILLCELL_X32 FILLER_114_1304 ();
 FILLCELL_X32 FILLER_114_1336 ();
 FILLCELL_X32 FILLER_114_1368 ();
 FILLCELL_X32 FILLER_114_1400 ();
 FILLCELL_X32 FILLER_114_1432 ();
 FILLCELL_X32 FILLER_114_1464 ();
 FILLCELL_X32 FILLER_114_1496 ();
 FILLCELL_X32 FILLER_114_1528 ();
 FILLCELL_X32 FILLER_114_1560 ();
 FILLCELL_X32 FILLER_114_1592 ();
 FILLCELL_X32 FILLER_114_1624 ();
 FILLCELL_X32 FILLER_114_1656 ();
 FILLCELL_X32 FILLER_114_1688 ();
 FILLCELL_X4 FILLER_114_1720 ();
 FILLCELL_X2 FILLER_114_1724 ();
 FILLCELL_X1 FILLER_114_1726 ();
 FILLCELL_X32 FILLER_114_1731 ();
 FILLCELL_X4 FILLER_114_1766 ();
 FILLCELL_X2 FILLER_114_1770 ();
 FILLCELL_X1 FILLER_114_1772 ();
 FILLCELL_X2 FILLER_114_1776 ();
 FILLCELL_X4 FILLER_115_1 ();
 FILLCELL_X8 FILLER_115_26 ();
 FILLCELL_X4 FILLER_115_34 ();
 FILLCELL_X2 FILLER_115_38 ();
 FILLCELL_X1 FILLER_115_40 ();
 FILLCELL_X32 FILLER_115_58 ();
 FILLCELL_X32 FILLER_115_90 ();
 FILLCELL_X32 FILLER_115_122 ();
 FILLCELL_X32 FILLER_115_154 ();
 FILLCELL_X32 FILLER_115_186 ();
 FILLCELL_X32 FILLER_115_218 ();
 FILLCELL_X32 FILLER_115_250 ();
 FILLCELL_X32 FILLER_115_282 ();
 FILLCELL_X32 FILLER_115_314 ();
 FILLCELL_X32 FILLER_115_346 ();
 FILLCELL_X32 FILLER_115_378 ();
 FILLCELL_X32 FILLER_115_410 ();
 FILLCELL_X32 FILLER_115_442 ();
 FILLCELL_X32 FILLER_115_474 ();
 FILLCELL_X32 FILLER_115_506 ();
 FILLCELL_X32 FILLER_115_538 ();
 FILLCELL_X32 FILLER_115_570 ();
 FILLCELL_X32 FILLER_115_602 ();
 FILLCELL_X32 FILLER_115_634 ();
 FILLCELL_X32 FILLER_115_666 ();
 FILLCELL_X32 FILLER_115_698 ();
 FILLCELL_X32 FILLER_115_730 ();
 FILLCELL_X32 FILLER_115_762 ();
 FILLCELL_X32 FILLER_115_794 ();
 FILLCELL_X32 FILLER_115_826 ();
 FILLCELL_X32 FILLER_115_858 ();
 FILLCELL_X32 FILLER_115_890 ();
 FILLCELL_X32 FILLER_115_922 ();
 FILLCELL_X32 FILLER_115_954 ();
 FILLCELL_X32 FILLER_115_986 ();
 FILLCELL_X32 FILLER_115_1018 ();
 FILLCELL_X32 FILLER_115_1050 ();
 FILLCELL_X32 FILLER_115_1082 ();
 FILLCELL_X32 FILLER_115_1114 ();
 FILLCELL_X32 FILLER_115_1146 ();
 FILLCELL_X32 FILLER_115_1178 ();
 FILLCELL_X32 FILLER_115_1210 ();
 FILLCELL_X16 FILLER_115_1242 ();
 FILLCELL_X4 FILLER_115_1258 ();
 FILLCELL_X1 FILLER_115_1262 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X32 FILLER_115_1552 ();
 FILLCELL_X32 FILLER_115_1584 ();
 FILLCELL_X32 FILLER_115_1616 ();
 FILLCELL_X32 FILLER_115_1648 ();
 FILLCELL_X32 FILLER_115_1680 ();
 FILLCELL_X32 FILLER_115_1712 ();
 FILLCELL_X8 FILLER_115_1744 ();
 FILLCELL_X4 FILLER_115_1752 ();
 FILLCELL_X1 FILLER_115_1756 ();
 FILLCELL_X8 FILLER_115_1772 ();
 FILLCELL_X4 FILLER_115_1780 ();
 FILLCELL_X4 FILLER_115_1787 ();
 FILLCELL_X2 FILLER_115_1791 ();
 FILLCELL_X1 FILLER_115_1793 ();
 FILLCELL_X8 FILLER_116_28 ();
 FILLCELL_X4 FILLER_116_36 ();
 FILLCELL_X32 FILLER_116_53 ();
 FILLCELL_X32 FILLER_116_85 ();
 FILLCELL_X32 FILLER_116_117 ();
 FILLCELL_X32 FILLER_116_149 ();
 FILLCELL_X32 FILLER_116_181 ();
 FILLCELL_X32 FILLER_116_213 ();
 FILLCELL_X32 FILLER_116_245 ();
 FILLCELL_X32 FILLER_116_277 ();
 FILLCELL_X32 FILLER_116_309 ();
 FILLCELL_X32 FILLER_116_341 ();
 FILLCELL_X32 FILLER_116_373 ();
 FILLCELL_X32 FILLER_116_405 ();
 FILLCELL_X32 FILLER_116_437 ();
 FILLCELL_X32 FILLER_116_469 ();
 FILLCELL_X32 FILLER_116_501 ();
 FILLCELL_X32 FILLER_116_533 ();
 FILLCELL_X32 FILLER_116_565 ();
 FILLCELL_X32 FILLER_116_597 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X2 FILLER_116_824 ();
 FILLCELL_X1 FILLER_116_826 ();
 FILLCELL_X32 FILLER_116_834 ();
 FILLCELL_X32 FILLER_116_866 ();
 FILLCELL_X32 FILLER_116_898 ();
 FILLCELL_X32 FILLER_116_930 ();
 FILLCELL_X32 FILLER_116_962 ();
 FILLCELL_X32 FILLER_116_994 ();
 FILLCELL_X32 FILLER_116_1026 ();
 FILLCELL_X32 FILLER_116_1058 ();
 FILLCELL_X32 FILLER_116_1090 ();
 FILLCELL_X32 FILLER_116_1122 ();
 FILLCELL_X32 FILLER_116_1154 ();
 FILLCELL_X32 FILLER_116_1186 ();
 FILLCELL_X32 FILLER_116_1218 ();
 FILLCELL_X32 FILLER_116_1250 ();
 FILLCELL_X32 FILLER_116_1282 ();
 FILLCELL_X32 FILLER_116_1314 ();
 FILLCELL_X32 FILLER_116_1346 ();
 FILLCELL_X32 FILLER_116_1378 ();
 FILLCELL_X32 FILLER_116_1410 ();
 FILLCELL_X32 FILLER_116_1442 ();
 FILLCELL_X32 FILLER_116_1474 ();
 FILLCELL_X32 FILLER_116_1506 ();
 FILLCELL_X32 FILLER_116_1538 ();
 FILLCELL_X32 FILLER_116_1570 ();
 FILLCELL_X32 FILLER_116_1602 ();
 FILLCELL_X32 FILLER_116_1634 ();
 FILLCELL_X32 FILLER_116_1666 ();
 FILLCELL_X32 FILLER_116_1698 ();
 FILLCELL_X16 FILLER_116_1730 ();
 FILLCELL_X4 FILLER_116_1746 ();
 FILLCELL_X1 FILLER_116_1750 ();
 FILLCELL_X2 FILLER_116_1773 ();
 FILLCELL_X1 FILLER_116_1775 ();
 FILLCELL_X2 FILLER_116_1792 ();
 FILLCELL_X2 FILLER_117_1 ();
 FILLCELL_X1 FILLER_117_10 ();
 FILLCELL_X2 FILLER_117_21 ();
 FILLCELL_X1 FILLER_117_23 ();
 FILLCELL_X2 FILLER_117_34 ();
 FILLCELL_X2 FILLER_117_43 ();
 FILLCELL_X32 FILLER_117_48 ();
 FILLCELL_X32 FILLER_117_80 ();
 FILLCELL_X32 FILLER_117_112 ();
 FILLCELL_X32 FILLER_117_144 ();
 FILLCELL_X32 FILLER_117_176 ();
 FILLCELL_X32 FILLER_117_208 ();
 FILLCELL_X32 FILLER_117_240 ();
 FILLCELL_X32 FILLER_117_272 ();
 FILLCELL_X32 FILLER_117_304 ();
 FILLCELL_X32 FILLER_117_336 ();
 FILLCELL_X32 FILLER_117_368 ();
 FILLCELL_X32 FILLER_117_400 ();
 FILLCELL_X32 FILLER_117_432 ();
 FILLCELL_X32 FILLER_117_464 ();
 FILLCELL_X32 FILLER_117_496 ();
 FILLCELL_X32 FILLER_117_528 ();
 FILLCELL_X32 FILLER_117_560 ();
 FILLCELL_X32 FILLER_117_592 ();
 FILLCELL_X32 FILLER_117_624 ();
 FILLCELL_X32 FILLER_117_656 ();
 FILLCELL_X32 FILLER_117_688 ();
 FILLCELL_X32 FILLER_117_720 ();
 FILLCELL_X32 FILLER_117_752 ();
 FILLCELL_X32 FILLER_117_784 ();
 FILLCELL_X4 FILLER_117_816 ();
 FILLCELL_X2 FILLER_117_820 ();
 FILLCELL_X1 FILLER_117_822 ();
 FILLCELL_X4 FILLER_117_828 ();
 FILLCELL_X32 FILLER_117_836 ();
 FILLCELL_X32 FILLER_117_868 ();
 FILLCELL_X32 FILLER_117_900 ();
 FILLCELL_X32 FILLER_117_932 ();
 FILLCELL_X32 FILLER_117_964 ();
 FILLCELL_X32 FILLER_117_996 ();
 FILLCELL_X32 FILLER_117_1028 ();
 FILLCELL_X32 FILLER_117_1060 ();
 FILLCELL_X32 FILLER_117_1092 ();
 FILLCELL_X32 FILLER_117_1124 ();
 FILLCELL_X32 FILLER_117_1156 ();
 FILLCELL_X32 FILLER_117_1188 ();
 FILLCELL_X32 FILLER_117_1220 ();
 FILLCELL_X8 FILLER_117_1252 ();
 FILLCELL_X2 FILLER_117_1260 ();
 FILLCELL_X1 FILLER_117_1262 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X32 FILLER_117_1552 ();
 FILLCELL_X32 FILLER_117_1584 ();
 FILLCELL_X32 FILLER_117_1616 ();
 FILLCELL_X32 FILLER_117_1648 ();
 FILLCELL_X32 FILLER_117_1680 ();
 FILLCELL_X32 FILLER_117_1712 ();
 FILLCELL_X1 FILLER_117_1744 ();
 FILLCELL_X4 FILLER_117_1752 ();
 FILLCELL_X8 FILLER_117_1774 ();
 FILLCELL_X4 FILLER_117_1782 ();
 FILLCELL_X2 FILLER_117_1786 ();
 FILLCELL_X1 FILLER_117_1788 ();
 FILLCELL_X2 FILLER_117_1791 ();
 FILLCELL_X1 FILLER_117_1793 ();
 FILLCELL_X16 FILLER_118_1 ();
 FILLCELL_X4 FILLER_118_17 ();
 FILLCELL_X2 FILLER_118_21 ();
 FILLCELL_X4 FILLER_118_27 ();
 FILLCELL_X2 FILLER_118_31 ();
 FILLCELL_X1 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_42 ();
 FILLCELL_X32 FILLER_118_74 ();
 FILLCELL_X32 FILLER_118_106 ();
 FILLCELL_X32 FILLER_118_138 ();
 FILLCELL_X32 FILLER_118_170 ();
 FILLCELL_X32 FILLER_118_202 ();
 FILLCELL_X32 FILLER_118_234 ();
 FILLCELL_X32 FILLER_118_266 ();
 FILLCELL_X32 FILLER_118_298 ();
 FILLCELL_X32 FILLER_118_330 ();
 FILLCELL_X32 FILLER_118_362 ();
 FILLCELL_X32 FILLER_118_394 ();
 FILLCELL_X32 FILLER_118_426 ();
 FILLCELL_X32 FILLER_118_458 ();
 FILLCELL_X32 FILLER_118_490 ();
 FILLCELL_X32 FILLER_118_522 ();
 FILLCELL_X32 FILLER_118_554 ();
 FILLCELL_X32 FILLER_118_586 ();
 FILLCELL_X8 FILLER_118_618 ();
 FILLCELL_X4 FILLER_118_626 ();
 FILLCELL_X1 FILLER_118_630 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X16 FILLER_118_792 ();
 FILLCELL_X8 FILLER_118_808 ();
 FILLCELL_X4 FILLER_118_816 ();
 FILLCELL_X1 FILLER_118_820 ();
 FILLCELL_X32 FILLER_118_838 ();
 FILLCELL_X32 FILLER_118_870 ();
 FILLCELL_X32 FILLER_118_902 ();
 FILLCELL_X32 FILLER_118_934 ();
 FILLCELL_X32 FILLER_118_966 ();
 FILLCELL_X32 FILLER_118_998 ();
 FILLCELL_X32 FILLER_118_1030 ();
 FILLCELL_X32 FILLER_118_1062 ();
 FILLCELL_X32 FILLER_118_1094 ();
 FILLCELL_X32 FILLER_118_1126 ();
 FILLCELL_X32 FILLER_118_1158 ();
 FILLCELL_X32 FILLER_118_1190 ();
 FILLCELL_X32 FILLER_118_1222 ();
 FILLCELL_X32 FILLER_118_1254 ();
 FILLCELL_X32 FILLER_118_1286 ();
 FILLCELL_X32 FILLER_118_1318 ();
 FILLCELL_X32 FILLER_118_1350 ();
 FILLCELL_X32 FILLER_118_1382 ();
 FILLCELL_X32 FILLER_118_1414 ();
 FILLCELL_X32 FILLER_118_1446 ();
 FILLCELL_X32 FILLER_118_1478 ();
 FILLCELL_X32 FILLER_118_1510 ();
 FILLCELL_X32 FILLER_118_1542 ();
 FILLCELL_X32 FILLER_118_1574 ();
 FILLCELL_X32 FILLER_118_1606 ();
 FILLCELL_X32 FILLER_118_1638 ();
 FILLCELL_X32 FILLER_118_1670 ();
 FILLCELL_X16 FILLER_118_1702 ();
 FILLCELL_X1 FILLER_118_1718 ();
 FILLCELL_X16 FILLER_118_1731 ();
 FILLCELL_X4 FILLER_118_1747 ();
 FILLCELL_X2 FILLER_118_1751 ();
 FILLCELL_X16 FILLER_118_1762 ();
 FILLCELL_X8 FILLER_118_1778 ();
 FILLCELL_X4 FILLER_118_1786 ();
 FILLCELL_X1 FILLER_118_1790 ();
 FILLCELL_X1 FILLER_119_7 ();
 FILLCELL_X4 FILLER_119_18 ();
 FILLCELL_X1 FILLER_119_26 ();
 FILLCELL_X8 FILLER_119_36 ();
 FILLCELL_X4 FILLER_119_44 ();
 FILLCELL_X32 FILLER_119_61 ();
 FILLCELL_X32 FILLER_119_93 ();
 FILLCELL_X32 FILLER_119_125 ();
 FILLCELL_X32 FILLER_119_157 ();
 FILLCELL_X32 FILLER_119_189 ();
 FILLCELL_X32 FILLER_119_221 ();
 FILLCELL_X32 FILLER_119_253 ();
 FILLCELL_X32 FILLER_119_285 ();
 FILLCELL_X32 FILLER_119_317 ();
 FILLCELL_X32 FILLER_119_349 ();
 FILLCELL_X32 FILLER_119_381 ();
 FILLCELL_X32 FILLER_119_413 ();
 FILLCELL_X32 FILLER_119_445 ();
 FILLCELL_X32 FILLER_119_477 ();
 FILLCELL_X32 FILLER_119_509 ();
 FILLCELL_X32 FILLER_119_541 ();
 FILLCELL_X32 FILLER_119_573 ();
 FILLCELL_X32 FILLER_119_605 ();
 FILLCELL_X32 FILLER_119_637 ();
 FILLCELL_X32 FILLER_119_669 ();
 FILLCELL_X32 FILLER_119_701 ();
 FILLCELL_X32 FILLER_119_733 ();
 FILLCELL_X32 FILLER_119_765 ();
 FILLCELL_X16 FILLER_119_797 ();
 FILLCELL_X2 FILLER_119_813 ();
 FILLCELL_X1 FILLER_119_815 ();
 FILLCELL_X32 FILLER_119_834 ();
 FILLCELL_X4 FILLER_119_866 ();
 FILLCELL_X2 FILLER_119_870 ();
 FILLCELL_X32 FILLER_119_885 ();
 FILLCELL_X32 FILLER_119_917 ();
 FILLCELL_X32 FILLER_119_949 ();
 FILLCELL_X32 FILLER_119_981 ();
 FILLCELL_X32 FILLER_119_1013 ();
 FILLCELL_X32 FILLER_119_1045 ();
 FILLCELL_X32 FILLER_119_1077 ();
 FILLCELL_X32 FILLER_119_1109 ();
 FILLCELL_X32 FILLER_119_1141 ();
 FILLCELL_X32 FILLER_119_1173 ();
 FILLCELL_X32 FILLER_119_1205 ();
 FILLCELL_X16 FILLER_119_1237 ();
 FILLCELL_X8 FILLER_119_1253 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X32 FILLER_119_1552 ();
 FILLCELL_X32 FILLER_119_1584 ();
 FILLCELL_X32 FILLER_119_1616 ();
 FILLCELL_X32 FILLER_119_1648 ();
 FILLCELL_X32 FILLER_119_1680 ();
 FILLCELL_X1 FILLER_119_1712 ();
 FILLCELL_X16 FILLER_119_1732 ();
 FILLCELL_X8 FILLER_119_1748 ();
 FILLCELL_X1 FILLER_119_1756 ();
 FILLCELL_X2 FILLER_119_1763 ();
 FILLCELL_X1 FILLER_119_1765 ();
 FILLCELL_X4 FILLER_119_1769 ();
 FILLCELL_X1 FILLER_119_1773 ();
 FILLCELL_X2 FILLER_119_1777 ();
 FILLCELL_X1 FILLER_119_1779 ();
 FILLCELL_X2 FILLER_120_4 ();
 FILLCELL_X1 FILLER_120_6 ();
 FILLCELL_X16 FILLER_120_13 ();
 FILLCELL_X4 FILLER_120_29 ();
 FILLCELL_X1 FILLER_120_33 ();
 FILLCELL_X4 FILLER_120_38 ();
 FILLCELL_X2 FILLER_120_42 ();
 FILLCELL_X2 FILLER_120_49 ();
 FILLCELL_X1 FILLER_120_51 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X8 FILLER_120_792 ();
 FILLCELL_X4 FILLER_120_800 ();
 FILLCELL_X2 FILLER_120_804 ();
 FILLCELL_X1 FILLER_120_806 ();
 FILLCELL_X2 FILLER_120_812 ();
 FILLCELL_X2 FILLER_120_821 ();
 FILLCELL_X1 FILLER_120_827 ();
 FILLCELL_X4 FILLER_120_832 ();
 FILLCELL_X16 FILLER_120_849 ();
 FILLCELL_X2 FILLER_120_865 ();
 FILLCELL_X2 FILLER_120_878 ();
 FILLCELL_X32 FILLER_120_887 ();
 FILLCELL_X2 FILLER_120_919 ();
 FILLCELL_X1 FILLER_120_921 ();
 FILLCELL_X32 FILLER_120_936 ();
 FILLCELL_X32 FILLER_120_968 ();
 FILLCELL_X32 FILLER_120_1000 ();
 FILLCELL_X32 FILLER_120_1032 ();
 FILLCELL_X32 FILLER_120_1064 ();
 FILLCELL_X32 FILLER_120_1096 ();
 FILLCELL_X32 FILLER_120_1128 ();
 FILLCELL_X32 FILLER_120_1160 ();
 FILLCELL_X32 FILLER_120_1192 ();
 FILLCELL_X32 FILLER_120_1224 ();
 FILLCELL_X32 FILLER_120_1256 ();
 FILLCELL_X32 FILLER_120_1288 ();
 FILLCELL_X32 FILLER_120_1320 ();
 FILLCELL_X32 FILLER_120_1352 ();
 FILLCELL_X32 FILLER_120_1384 ();
 FILLCELL_X32 FILLER_120_1416 ();
 FILLCELL_X32 FILLER_120_1448 ();
 FILLCELL_X32 FILLER_120_1480 ();
 FILLCELL_X32 FILLER_120_1512 ();
 FILLCELL_X32 FILLER_120_1544 ();
 FILLCELL_X32 FILLER_120_1576 ();
 FILLCELL_X32 FILLER_120_1608 ();
 FILLCELL_X32 FILLER_120_1640 ();
 FILLCELL_X32 FILLER_120_1672 ();
 FILLCELL_X4 FILLER_120_1704 ();
 FILLCELL_X2 FILLER_120_1708 ();
 FILLCELL_X4 FILLER_120_1719 ();
 FILLCELL_X1 FILLER_120_1723 ();
 FILLCELL_X16 FILLER_120_1729 ();
 FILLCELL_X1 FILLER_120_1745 ();
 FILLCELL_X8 FILLER_120_1764 ();
 FILLCELL_X4 FILLER_120_1772 ();
 FILLCELL_X2 FILLER_120_1792 ();
 FILLCELL_X4 FILLER_121_1 ();
 FILLCELL_X2 FILLER_121_5 ();
 FILLCELL_X1 FILLER_121_15 ();
 FILLCELL_X8 FILLER_121_26 ();
 FILLCELL_X2 FILLER_121_47 ();
 FILLCELL_X1 FILLER_121_49 ();
 FILLCELL_X2 FILLER_121_53 ();
 FILLCELL_X1 FILLER_121_55 ();
 FILLCELL_X1 FILLER_121_63 ();
 FILLCELL_X16 FILLER_121_70 ();
 FILLCELL_X8 FILLER_121_86 ();
 FILLCELL_X4 FILLER_121_94 ();
 FILLCELL_X2 FILLER_121_98 ();
 FILLCELL_X1 FILLER_121_100 ();
 FILLCELL_X32 FILLER_121_105 ();
 FILLCELL_X32 FILLER_121_137 ();
 FILLCELL_X32 FILLER_121_169 ();
 FILLCELL_X32 FILLER_121_201 ();
 FILLCELL_X32 FILLER_121_233 ();
 FILLCELL_X32 FILLER_121_265 ();
 FILLCELL_X32 FILLER_121_297 ();
 FILLCELL_X32 FILLER_121_329 ();
 FILLCELL_X32 FILLER_121_361 ();
 FILLCELL_X32 FILLER_121_393 ();
 FILLCELL_X32 FILLER_121_425 ();
 FILLCELL_X32 FILLER_121_457 ();
 FILLCELL_X32 FILLER_121_489 ();
 FILLCELL_X32 FILLER_121_521 ();
 FILLCELL_X32 FILLER_121_553 ();
 FILLCELL_X32 FILLER_121_585 ();
 FILLCELL_X32 FILLER_121_617 ();
 FILLCELL_X32 FILLER_121_649 ();
 FILLCELL_X32 FILLER_121_681 ();
 FILLCELL_X32 FILLER_121_713 ();
 FILLCELL_X32 FILLER_121_745 ();
 FILLCELL_X32 FILLER_121_777 ();
 FILLCELL_X4 FILLER_121_809 ();
 FILLCELL_X16 FILLER_121_839 ();
 FILLCELL_X4 FILLER_121_855 ();
 FILLCELL_X2 FILLER_121_859 ();
 FILLCELL_X1 FILLER_121_861 ();
 FILLCELL_X16 FILLER_121_867 ();
 FILLCELL_X4 FILLER_121_883 ();
 FILLCELL_X16 FILLER_121_900 ();
 FILLCELL_X4 FILLER_121_916 ();
 FILLCELL_X2 FILLER_121_920 ();
 FILLCELL_X1 FILLER_121_922 ();
 FILLCELL_X32 FILLER_121_934 ();
 FILLCELL_X32 FILLER_121_966 ();
 FILLCELL_X32 FILLER_121_998 ();
 FILLCELL_X32 FILLER_121_1030 ();
 FILLCELL_X32 FILLER_121_1062 ();
 FILLCELL_X32 FILLER_121_1094 ();
 FILLCELL_X32 FILLER_121_1126 ();
 FILLCELL_X32 FILLER_121_1158 ();
 FILLCELL_X32 FILLER_121_1190 ();
 FILLCELL_X32 FILLER_121_1222 ();
 FILLCELL_X8 FILLER_121_1254 ();
 FILLCELL_X1 FILLER_121_1262 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X32 FILLER_121_1552 ();
 FILLCELL_X32 FILLER_121_1584 ();
 FILLCELL_X32 FILLER_121_1616 ();
 FILLCELL_X32 FILLER_121_1648 ();
 FILLCELL_X32 FILLER_121_1680 ();
 FILLCELL_X32 FILLER_121_1712 ();
 FILLCELL_X2 FILLER_121_1744 ();
 FILLCELL_X1 FILLER_121_1748 ();
 FILLCELL_X8 FILLER_121_1765 ();
 FILLCELL_X2 FILLER_121_1776 ();
 FILLCELL_X1 FILLER_121_1778 ();
 FILLCELL_X2 FILLER_121_1783 ();
 FILLCELL_X2 FILLER_121_1791 ();
 FILLCELL_X1 FILLER_121_1793 ();
 FILLCELL_X2 FILLER_122_4 ();
 FILLCELL_X1 FILLER_122_9 ();
 FILLCELL_X2 FILLER_122_13 ();
 FILLCELL_X16 FILLER_122_21 ();
 FILLCELL_X1 FILLER_122_40 ();
 FILLCELL_X1 FILLER_122_44 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X16 FILLER_122_792 ();
 FILLCELL_X4 FILLER_122_808 ();
 FILLCELL_X2 FILLER_122_812 ();
 FILLCELL_X1 FILLER_122_814 ();
 FILLCELL_X16 FILLER_122_834 ();
 FILLCELL_X8 FILLER_122_850 ();
 FILLCELL_X32 FILLER_122_867 ();
 FILLCELL_X16 FILLER_122_899 ();
 FILLCELL_X1 FILLER_122_915 ();
 FILLCELL_X32 FILLER_122_934 ();
 FILLCELL_X32 FILLER_122_966 ();
 FILLCELL_X32 FILLER_122_998 ();
 FILLCELL_X32 FILLER_122_1030 ();
 FILLCELL_X32 FILLER_122_1062 ();
 FILLCELL_X32 FILLER_122_1094 ();
 FILLCELL_X32 FILLER_122_1126 ();
 FILLCELL_X32 FILLER_122_1158 ();
 FILLCELL_X32 FILLER_122_1190 ();
 FILLCELL_X32 FILLER_122_1222 ();
 FILLCELL_X32 FILLER_122_1254 ();
 FILLCELL_X32 FILLER_122_1286 ();
 FILLCELL_X32 FILLER_122_1318 ();
 FILLCELL_X32 FILLER_122_1350 ();
 FILLCELL_X32 FILLER_122_1382 ();
 FILLCELL_X32 FILLER_122_1414 ();
 FILLCELL_X32 FILLER_122_1446 ();
 FILLCELL_X32 FILLER_122_1478 ();
 FILLCELL_X32 FILLER_122_1510 ();
 FILLCELL_X32 FILLER_122_1542 ();
 FILLCELL_X32 FILLER_122_1574 ();
 FILLCELL_X32 FILLER_122_1606 ();
 FILLCELL_X32 FILLER_122_1638 ();
 FILLCELL_X32 FILLER_122_1670 ();
 FILLCELL_X32 FILLER_122_1702 ();
 FILLCELL_X4 FILLER_122_1734 ();
 FILLCELL_X2 FILLER_122_1738 ();
 FILLCELL_X4 FILLER_122_1752 ();
 FILLCELL_X1 FILLER_122_1756 ();
 FILLCELL_X8 FILLER_122_1767 ();
 FILLCELL_X4 FILLER_122_1775 ();
 FILLCELL_X4 FILLER_122_1782 ();
 FILLCELL_X2 FILLER_122_1786 ();
 FILLCELL_X1 FILLER_122_1788 ();
 FILLCELL_X2 FILLER_122_1795 ();
 FILLCELL_X8 FILLER_123_1 ();
 FILLCELL_X4 FILLER_123_9 ();
 FILLCELL_X2 FILLER_123_13 ();
 FILLCELL_X4 FILLER_123_23 ();
 FILLCELL_X2 FILLER_123_33 ();
 FILLCELL_X8 FILLER_123_48 ();
 FILLCELL_X4 FILLER_123_56 ();
 FILLCELL_X1 FILLER_123_60 ();
 FILLCELL_X32 FILLER_123_71 ();
 FILLCELL_X32 FILLER_123_103 ();
 FILLCELL_X32 FILLER_123_135 ();
 FILLCELL_X32 FILLER_123_167 ();
 FILLCELL_X32 FILLER_123_199 ();
 FILLCELL_X32 FILLER_123_231 ();
 FILLCELL_X32 FILLER_123_263 ();
 FILLCELL_X32 FILLER_123_295 ();
 FILLCELL_X32 FILLER_123_327 ();
 FILLCELL_X32 FILLER_123_359 ();
 FILLCELL_X32 FILLER_123_391 ();
 FILLCELL_X32 FILLER_123_423 ();
 FILLCELL_X32 FILLER_123_455 ();
 FILLCELL_X32 FILLER_123_487 ();
 FILLCELL_X32 FILLER_123_519 ();
 FILLCELL_X32 FILLER_123_551 ();
 FILLCELL_X32 FILLER_123_583 ();
 FILLCELL_X32 FILLER_123_615 ();
 FILLCELL_X32 FILLER_123_647 ();
 FILLCELL_X32 FILLER_123_679 ();
 FILLCELL_X32 FILLER_123_711 ();
 FILLCELL_X32 FILLER_123_743 ();
 FILLCELL_X32 FILLER_123_775 ();
 FILLCELL_X8 FILLER_123_807 ();
 FILLCELL_X4 FILLER_123_815 ();
 FILLCELL_X2 FILLER_123_819 ();
 FILLCELL_X8 FILLER_123_830 ();
 FILLCELL_X4 FILLER_123_838 ();
 FILLCELL_X2 FILLER_123_842 ();
 FILLCELL_X1 FILLER_123_844 ();
 FILLCELL_X32 FILLER_123_869 ();
 FILLCELL_X32 FILLER_123_901 ();
 FILLCELL_X32 FILLER_123_933 ();
 FILLCELL_X32 FILLER_123_965 ();
 FILLCELL_X32 FILLER_123_997 ();
 FILLCELL_X32 FILLER_123_1029 ();
 FILLCELL_X32 FILLER_123_1061 ();
 FILLCELL_X32 FILLER_123_1093 ();
 FILLCELL_X32 FILLER_123_1125 ();
 FILLCELL_X32 FILLER_123_1157 ();
 FILLCELL_X32 FILLER_123_1189 ();
 FILLCELL_X32 FILLER_123_1221 ();
 FILLCELL_X8 FILLER_123_1253 ();
 FILLCELL_X2 FILLER_123_1261 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X32 FILLER_123_1552 ();
 FILLCELL_X32 FILLER_123_1584 ();
 FILLCELL_X32 FILLER_123_1616 ();
 FILLCELL_X32 FILLER_123_1648 ();
 FILLCELL_X32 FILLER_123_1680 ();
 FILLCELL_X32 FILLER_123_1712 ();
 FILLCELL_X16 FILLER_123_1744 ();
 FILLCELL_X2 FILLER_123_1760 ();
 FILLCELL_X1 FILLER_123_1762 ();
 FILLCELL_X4 FILLER_123_1765 ();
 FILLCELL_X1 FILLER_123_1769 ();
 FILLCELL_X16 FILLER_123_1773 ();
 FILLCELL_X8 FILLER_123_1789 ();
 FILLCELL_X4 FILLER_124_1 ();
 FILLCELL_X4 FILLER_124_16 ();
 FILLCELL_X2 FILLER_124_20 ();
 FILLCELL_X16 FILLER_124_25 ();
 FILLCELL_X8 FILLER_124_41 ();
 FILLCELL_X32 FILLER_124_61 ();
 FILLCELL_X32 FILLER_124_93 ();
 FILLCELL_X32 FILLER_124_125 ();
 FILLCELL_X32 FILLER_124_157 ();
 FILLCELL_X32 FILLER_124_189 ();
 FILLCELL_X32 FILLER_124_221 ();
 FILLCELL_X32 FILLER_124_253 ();
 FILLCELL_X32 FILLER_124_285 ();
 FILLCELL_X32 FILLER_124_317 ();
 FILLCELL_X32 FILLER_124_349 ();
 FILLCELL_X32 FILLER_124_381 ();
 FILLCELL_X32 FILLER_124_413 ();
 FILLCELL_X32 FILLER_124_445 ();
 FILLCELL_X32 FILLER_124_477 ();
 FILLCELL_X32 FILLER_124_509 ();
 FILLCELL_X32 FILLER_124_541 ();
 FILLCELL_X32 FILLER_124_573 ();
 FILLCELL_X16 FILLER_124_605 ();
 FILLCELL_X8 FILLER_124_621 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X32 FILLER_124_1144 ();
 FILLCELL_X32 FILLER_124_1176 ();
 FILLCELL_X32 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_124_1240 ();
 FILLCELL_X32 FILLER_124_1272 ();
 FILLCELL_X32 FILLER_124_1304 ();
 FILLCELL_X32 FILLER_124_1336 ();
 FILLCELL_X32 FILLER_124_1368 ();
 FILLCELL_X32 FILLER_124_1400 ();
 FILLCELL_X32 FILLER_124_1432 ();
 FILLCELL_X32 FILLER_124_1464 ();
 FILLCELL_X32 FILLER_124_1496 ();
 FILLCELL_X32 FILLER_124_1528 ();
 FILLCELL_X32 FILLER_124_1560 ();
 FILLCELL_X32 FILLER_124_1592 ();
 FILLCELL_X32 FILLER_124_1624 ();
 FILLCELL_X32 FILLER_124_1656 ();
 FILLCELL_X32 FILLER_124_1688 ();
 FILLCELL_X32 FILLER_124_1720 ();
 FILLCELL_X4 FILLER_124_1752 ();
 FILLCELL_X2 FILLER_124_1756 ();
 FILLCELL_X1 FILLER_124_1758 ();
 FILLCELL_X2 FILLER_124_1762 ();
 FILLCELL_X1 FILLER_124_1764 ();
 FILLCELL_X2 FILLER_124_1768 ();
 FILLCELL_X2 FILLER_124_1789 ();
 FILLCELL_X4 FILLER_125_4 ();
 FILLCELL_X1 FILLER_125_12 ();
 FILLCELL_X16 FILLER_125_23 ();
 FILLCELL_X8 FILLER_125_42 ();
 FILLCELL_X4 FILLER_125_50 ();
 FILLCELL_X2 FILLER_125_54 ();
 FILLCELL_X32 FILLER_125_58 ();
 FILLCELL_X32 FILLER_125_90 ();
 FILLCELL_X32 FILLER_125_122 ();
 FILLCELL_X32 FILLER_125_154 ();
 FILLCELL_X32 FILLER_125_186 ();
 FILLCELL_X32 FILLER_125_218 ();
 FILLCELL_X32 FILLER_125_250 ();
 FILLCELL_X32 FILLER_125_282 ();
 FILLCELL_X32 FILLER_125_314 ();
 FILLCELL_X32 FILLER_125_346 ();
 FILLCELL_X32 FILLER_125_378 ();
 FILLCELL_X32 FILLER_125_410 ();
 FILLCELL_X32 FILLER_125_442 ();
 FILLCELL_X32 FILLER_125_474 ();
 FILLCELL_X32 FILLER_125_506 ();
 FILLCELL_X32 FILLER_125_538 ();
 FILLCELL_X32 FILLER_125_570 ();
 FILLCELL_X32 FILLER_125_602 ();
 FILLCELL_X32 FILLER_125_634 ();
 FILLCELL_X32 FILLER_125_666 ();
 FILLCELL_X32 FILLER_125_698 ();
 FILLCELL_X32 FILLER_125_730 ();
 FILLCELL_X32 FILLER_125_762 ();
 FILLCELL_X32 FILLER_125_794 ();
 FILLCELL_X32 FILLER_125_826 ();
 FILLCELL_X32 FILLER_125_858 ();
 FILLCELL_X32 FILLER_125_890 ();
 FILLCELL_X32 FILLER_125_922 ();
 FILLCELL_X32 FILLER_125_954 ();
 FILLCELL_X32 FILLER_125_986 ();
 FILLCELL_X32 FILLER_125_1018 ();
 FILLCELL_X32 FILLER_125_1050 ();
 FILLCELL_X32 FILLER_125_1082 ();
 FILLCELL_X32 FILLER_125_1114 ();
 FILLCELL_X32 FILLER_125_1146 ();
 FILLCELL_X32 FILLER_125_1178 ();
 FILLCELL_X32 FILLER_125_1210 ();
 FILLCELL_X16 FILLER_125_1242 ();
 FILLCELL_X4 FILLER_125_1258 ();
 FILLCELL_X1 FILLER_125_1262 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X32 FILLER_125_1648 ();
 FILLCELL_X32 FILLER_125_1680 ();
 FILLCELL_X8 FILLER_125_1712 ();
 FILLCELL_X2 FILLER_125_1720 ();
 FILLCELL_X4 FILLER_125_1724 ();
 FILLCELL_X2 FILLER_125_1728 ();
 FILLCELL_X1 FILLER_125_1730 ();
 FILLCELL_X16 FILLER_125_1745 ();
 FILLCELL_X4 FILLER_125_1761 ();
 FILLCELL_X2 FILLER_125_1765 ();
 FILLCELL_X1 FILLER_125_1781 ();
 FILLCELL_X4 FILLER_125_1789 ();
 FILLCELL_X1 FILLER_125_1796 ();
 FILLCELL_X1 FILLER_126_1 ();
 FILLCELL_X2 FILLER_126_5 ();
 FILLCELL_X4 FILLER_126_17 ();
 FILLCELL_X2 FILLER_126_21 ();
 FILLCELL_X1 FILLER_126_35 ();
 FILLCELL_X32 FILLER_126_38 ();
 FILLCELL_X32 FILLER_126_70 ();
 FILLCELL_X32 FILLER_126_102 ();
 FILLCELL_X32 FILLER_126_134 ();
 FILLCELL_X32 FILLER_126_166 ();
 FILLCELL_X32 FILLER_126_198 ();
 FILLCELL_X32 FILLER_126_230 ();
 FILLCELL_X32 FILLER_126_262 ();
 FILLCELL_X32 FILLER_126_294 ();
 FILLCELL_X32 FILLER_126_326 ();
 FILLCELL_X32 FILLER_126_358 ();
 FILLCELL_X32 FILLER_126_390 ();
 FILLCELL_X32 FILLER_126_422 ();
 FILLCELL_X32 FILLER_126_454 ();
 FILLCELL_X32 FILLER_126_486 ();
 FILLCELL_X32 FILLER_126_518 ();
 FILLCELL_X32 FILLER_126_550 ();
 FILLCELL_X32 FILLER_126_582 ();
 FILLCELL_X16 FILLER_126_614 ();
 FILLCELL_X1 FILLER_126_630 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X1 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_994 ();
 FILLCELL_X32 FILLER_126_1026 ();
 FILLCELL_X32 FILLER_126_1058 ();
 FILLCELL_X32 FILLER_126_1090 ();
 FILLCELL_X32 FILLER_126_1122 ();
 FILLCELL_X32 FILLER_126_1154 ();
 FILLCELL_X32 FILLER_126_1186 ();
 FILLCELL_X32 FILLER_126_1218 ();
 FILLCELL_X32 FILLER_126_1250 ();
 FILLCELL_X32 FILLER_126_1282 ();
 FILLCELL_X32 FILLER_126_1314 ();
 FILLCELL_X32 FILLER_126_1346 ();
 FILLCELL_X32 FILLER_126_1378 ();
 FILLCELL_X32 FILLER_126_1410 ();
 FILLCELL_X32 FILLER_126_1442 ();
 FILLCELL_X32 FILLER_126_1474 ();
 FILLCELL_X32 FILLER_126_1506 ();
 FILLCELL_X32 FILLER_126_1538 ();
 FILLCELL_X32 FILLER_126_1570 ();
 FILLCELL_X32 FILLER_126_1602 ();
 FILLCELL_X32 FILLER_126_1634 ();
 FILLCELL_X32 FILLER_126_1666 ();
 FILLCELL_X16 FILLER_126_1698 ();
 FILLCELL_X1 FILLER_126_1714 ();
 FILLCELL_X8 FILLER_126_1726 ();
 FILLCELL_X1 FILLER_126_1734 ();
 FILLCELL_X16 FILLER_126_1741 ();
 FILLCELL_X1 FILLER_126_1757 ();
 FILLCELL_X8 FILLER_126_1761 ();
 FILLCELL_X4 FILLER_126_1769 ();
 FILLCELL_X2 FILLER_126_1773 ();
 FILLCELL_X1 FILLER_126_1779 ();
 FILLCELL_X1 FILLER_126_1796 ();
 FILLCELL_X16 FILLER_127_4 ();
 FILLCELL_X4 FILLER_127_20 ();
 FILLCELL_X2 FILLER_127_24 ();
 FILLCELL_X32 FILLER_127_32 ();
 FILLCELL_X32 FILLER_127_64 ();
 FILLCELL_X32 FILLER_127_96 ();
 FILLCELL_X32 FILLER_127_128 ();
 FILLCELL_X32 FILLER_127_160 ();
 FILLCELL_X32 FILLER_127_192 ();
 FILLCELL_X32 FILLER_127_224 ();
 FILLCELL_X32 FILLER_127_256 ();
 FILLCELL_X32 FILLER_127_288 ();
 FILLCELL_X32 FILLER_127_320 ();
 FILLCELL_X32 FILLER_127_352 ();
 FILLCELL_X32 FILLER_127_384 ();
 FILLCELL_X32 FILLER_127_416 ();
 FILLCELL_X32 FILLER_127_448 ();
 FILLCELL_X32 FILLER_127_480 ();
 FILLCELL_X32 FILLER_127_512 ();
 FILLCELL_X32 FILLER_127_544 ();
 FILLCELL_X32 FILLER_127_576 ();
 FILLCELL_X32 FILLER_127_608 ();
 FILLCELL_X32 FILLER_127_640 ();
 FILLCELL_X32 FILLER_127_672 ();
 FILLCELL_X32 FILLER_127_704 ();
 FILLCELL_X32 FILLER_127_736 ();
 FILLCELL_X32 FILLER_127_768 ();
 FILLCELL_X32 FILLER_127_800 ();
 FILLCELL_X32 FILLER_127_832 ();
 FILLCELL_X32 FILLER_127_864 ();
 FILLCELL_X32 FILLER_127_896 ();
 FILLCELL_X16 FILLER_127_928 ();
 FILLCELL_X4 FILLER_127_944 ();
 FILLCELL_X16 FILLER_127_961 ();
 FILLCELL_X2 FILLER_127_977 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X32 FILLER_127_1089 ();
 FILLCELL_X32 FILLER_127_1121 ();
 FILLCELL_X32 FILLER_127_1153 ();
 FILLCELL_X32 FILLER_127_1185 ();
 FILLCELL_X32 FILLER_127_1217 ();
 FILLCELL_X8 FILLER_127_1249 ();
 FILLCELL_X4 FILLER_127_1257 ();
 FILLCELL_X2 FILLER_127_1261 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X32 FILLER_127_1584 ();
 FILLCELL_X32 FILLER_127_1616 ();
 FILLCELL_X32 FILLER_127_1648 ();
 FILLCELL_X32 FILLER_127_1680 ();
 FILLCELL_X8 FILLER_127_1712 ();
 FILLCELL_X2 FILLER_127_1720 ();
 FILLCELL_X16 FILLER_127_1732 ();
 FILLCELL_X4 FILLER_127_1748 ();
 FILLCELL_X2 FILLER_127_1752 ();
 FILLCELL_X1 FILLER_127_1764 ();
 FILLCELL_X4 FILLER_127_1774 ();
 FILLCELL_X4 FILLER_127_1781 ();
 FILLCELL_X2 FILLER_127_1785 ();
 FILLCELL_X1 FILLER_127_1787 ();
 FILLCELL_X2 FILLER_127_1791 ();
 FILLCELL_X1 FILLER_127_1793 ();
 FILLCELL_X4 FILLER_128_1 ();
 FILLCELL_X1 FILLER_128_5 ();
 FILLCELL_X4 FILLER_128_24 ();
 FILLCELL_X2 FILLER_128_28 ();
 FILLCELL_X1 FILLER_128_30 ();
 FILLCELL_X4 FILLER_128_45 ();
 FILLCELL_X32 FILLER_128_59 ();
 FILLCELL_X32 FILLER_128_91 ();
 FILLCELL_X32 FILLER_128_123 ();
 FILLCELL_X32 FILLER_128_155 ();
 FILLCELL_X32 FILLER_128_187 ();
 FILLCELL_X32 FILLER_128_219 ();
 FILLCELL_X32 FILLER_128_251 ();
 FILLCELL_X32 FILLER_128_283 ();
 FILLCELL_X32 FILLER_128_315 ();
 FILLCELL_X32 FILLER_128_347 ();
 FILLCELL_X32 FILLER_128_379 ();
 FILLCELL_X32 FILLER_128_411 ();
 FILLCELL_X32 FILLER_128_443 ();
 FILLCELL_X32 FILLER_128_475 ();
 FILLCELL_X32 FILLER_128_507 ();
 FILLCELL_X32 FILLER_128_539 ();
 FILLCELL_X32 FILLER_128_571 ();
 FILLCELL_X16 FILLER_128_603 ();
 FILLCELL_X8 FILLER_128_619 ();
 FILLCELL_X4 FILLER_128_627 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X2 FILLER_128_824 ();
 FILLCELL_X1 FILLER_128_826 ();
 FILLCELL_X32 FILLER_128_832 ();
 FILLCELL_X32 FILLER_128_864 ();
 FILLCELL_X32 FILLER_128_896 ();
 FILLCELL_X16 FILLER_128_928 ();
 FILLCELL_X4 FILLER_128_944 ();
 FILLCELL_X1 FILLER_128_948 ();
 FILLCELL_X32 FILLER_128_956 ();
 FILLCELL_X32 FILLER_128_988 ();
 FILLCELL_X32 FILLER_128_1020 ();
 FILLCELL_X32 FILLER_128_1052 ();
 FILLCELL_X32 FILLER_128_1084 ();
 FILLCELL_X32 FILLER_128_1116 ();
 FILLCELL_X32 FILLER_128_1148 ();
 FILLCELL_X32 FILLER_128_1180 ();
 FILLCELL_X32 FILLER_128_1212 ();
 FILLCELL_X32 FILLER_128_1244 ();
 FILLCELL_X32 FILLER_128_1276 ();
 FILLCELL_X32 FILLER_128_1308 ();
 FILLCELL_X32 FILLER_128_1340 ();
 FILLCELL_X32 FILLER_128_1372 ();
 FILLCELL_X32 FILLER_128_1404 ();
 FILLCELL_X32 FILLER_128_1436 ();
 FILLCELL_X32 FILLER_128_1468 ();
 FILLCELL_X32 FILLER_128_1500 ();
 FILLCELL_X32 FILLER_128_1532 ();
 FILLCELL_X32 FILLER_128_1564 ();
 FILLCELL_X32 FILLER_128_1596 ();
 FILLCELL_X32 FILLER_128_1628 ();
 FILLCELL_X32 FILLER_128_1660 ();
 FILLCELL_X32 FILLER_128_1692 ();
 FILLCELL_X16 FILLER_128_1724 ();
 FILLCELL_X8 FILLER_128_1740 ();
 FILLCELL_X4 FILLER_128_1748 ();
 FILLCELL_X16 FILLER_128_1757 ();
 FILLCELL_X8 FILLER_128_1773 ();
 FILLCELL_X4 FILLER_128_1781 ();
 FILLCELL_X8 FILLER_128_1788 ();
 FILLCELL_X1 FILLER_128_1796 ();
 FILLCELL_X1 FILLER_129_1 ();
 FILLCELL_X1 FILLER_129_14 ();
 FILLCELL_X1 FILLER_129_28 ();
 FILLCELL_X8 FILLER_129_32 ();
 FILLCELL_X2 FILLER_129_46 ();
 FILLCELL_X1 FILLER_129_48 ();
 FILLCELL_X2 FILLER_129_51 ();
 FILLCELL_X32 FILLER_129_56 ();
 FILLCELL_X32 FILLER_129_88 ();
 FILLCELL_X32 FILLER_129_120 ();
 FILLCELL_X32 FILLER_129_152 ();
 FILLCELL_X32 FILLER_129_184 ();
 FILLCELL_X32 FILLER_129_216 ();
 FILLCELL_X32 FILLER_129_248 ();
 FILLCELL_X32 FILLER_129_280 ();
 FILLCELL_X32 FILLER_129_312 ();
 FILLCELL_X32 FILLER_129_344 ();
 FILLCELL_X32 FILLER_129_376 ();
 FILLCELL_X32 FILLER_129_408 ();
 FILLCELL_X32 FILLER_129_440 ();
 FILLCELL_X32 FILLER_129_472 ();
 FILLCELL_X32 FILLER_129_504 ();
 FILLCELL_X32 FILLER_129_536 ();
 FILLCELL_X32 FILLER_129_568 ();
 FILLCELL_X32 FILLER_129_600 ();
 FILLCELL_X32 FILLER_129_632 ();
 FILLCELL_X32 FILLER_129_664 ();
 FILLCELL_X32 FILLER_129_696 ();
 FILLCELL_X32 FILLER_129_728 ();
 FILLCELL_X32 FILLER_129_760 ();
 FILLCELL_X32 FILLER_129_792 ();
 FILLCELL_X32 FILLER_129_824 ();
 FILLCELL_X32 FILLER_129_856 ();
 FILLCELL_X32 FILLER_129_888 ();
 FILLCELL_X2 FILLER_129_920 ();
 FILLCELL_X16 FILLER_129_931 ();
 FILLCELL_X1 FILLER_129_947 ();
 FILLCELL_X1 FILLER_129_953 ();
 FILLCELL_X2 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_966 ();
 FILLCELL_X32 FILLER_129_998 ();
 FILLCELL_X32 FILLER_129_1030 ();
 FILLCELL_X32 FILLER_129_1062 ();
 FILLCELL_X32 FILLER_129_1094 ();
 FILLCELL_X32 FILLER_129_1126 ();
 FILLCELL_X32 FILLER_129_1158 ();
 FILLCELL_X32 FILLER_129_1190 ();
 FILLCELL_X32 FILLER_129_1222 ();
 FILLCELL_X8 FILLER_129_1254 ();
 FILLCELL_X1 FILLER_129_1262 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X32 FILLER_129_1584 ();
 FILLCELL_X32 FILLER_129_1616 ();
 FILLCELL_X32 FILLER_129_1648 ();
 FILLCELL_X16 FILLER_129_1680 ();
 FILLCELL_X8 FILLER_129_1696 ();
 FILLCELL_X4 FILLER_129_1704 ();
 FILLCELL_X2 FILLER_129_1708 ();
 FILLCELL_X1 FILLER_129_1735 ();
 FILLCELL_X1 FILLER_129_1741 ();
 FILLCELL_X1 FILLER_129_1745 ();
 FILLCELL_X2 FILLER_129_1749 ();
 FILLCELL_X1 FILLER_129_1751 ();
 FILLCELL_X2 FILLER_129_1759 ();
 FILLCELL_X1 FILLER_129_1761 ();
 FILLCELL_X4 FILLER_129_1769 ();
 FILLCELL_X2 FILLER_129_1773 ();
 FILLCELL_X1 FILLER_129_1778 ();
 FILLCELL_X4 FILLER_129_1783 ();
 FILLCELL_X4 FILLER_129_1790 ();
 FILLCELL_X2 FILLER_129_1794 ();
 FILLCELL_X1 FILLER_129_1796 ();
 FILLCELL_X8 FILLER_130_1 ();
 FILLCELL_X16 FILLER_130_14 ();
 FILLCELL_X8 FILLER_130_30 ();
 FILLCELL_X4 FILLER_130_38 ();
 FILLCELL_X1 FILLER_130_46 ();
 FILLCELL_X32 FILLER_130_58 ();
 FILLCELL_X32 FILLER_130_90 ();
 FILLCELL_X32 FILLER_130_122 ();
 FILLCELL_X32 FILLER_130_154 ();
 FILLCELL_X32 FILLER_130_186 ();
 FILLCELL_X32 FILLER_130_218 ();
 FILLCELL_X32 FILLER_130_250 ();
 FILLCELL_X32 FILLER_130_282 ();
 FILLCELL_X32 FILLER_130_314 ();
 FILLCELL_X32 FILLER_130_346 ();
 FILLCELL_X32 FILLER_130_378 ();
 FILLCELL_X32 FILLER_130_410 ();
 FILLCELL_X32 FILLER_130_442 ();
 FILLCELL_X32 FILLER_130_474 ();
 FILLCELL_X32 FILLER_130_506 ();
 FILLCELL_X32 FILLER_130_538 ();
 FILLCELL_X32 FILLER_130_570 ();
 FILLCELL_X16 FILLER_130_602 ();
 FILLCELL_X8 FILLER_130_618 ();
 FILLCELL_X4 FILLER_130_626 ();
 FILLCELL_X1 FILLER_130_630 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X16 FILLER_130_792 ();
 FILLCELL_X8 FILLER_130_808 ();
 FILLCELL_X1 FILLER_130_816 ();
 FILLCELL_X32 FILLER_130_834 ();
 FILLCELL_X32 FILLER_130_866 ();
 FILLCELL_X16 FILLER_130_898 ();
 FILLCELL_X8 FILLER_130_914 ();
 FILLCELL_X4 FILLER_130_922 ();
 FILLCELL_X2 FILLER_130_926 ();
 FILLCELL_X1 FILLER_130_928 ();
 FILLCELL_X4 FILLER_130_936 ();
 FILLCELL_X2 FILLER_130_940 ();
 FILLCELL_X1 FILLER_130_942 ();
 FILLCELL_X4 FILLER_130_951 ();
 FILLCELL_X2 FILLER_130_955 ();
 FILLCELL_X32 FILLER_130_970 ();
 FILLCELL_X32 FILLER_130_1002 ();
 FILLCELL_X32 FILLER_130_1034 ();
 FILLCELL_X32 FILLER_130_1066 ();
 FILLCELL_X32 FILLER_130_1098 ();
 FILLCELL_X32 FILLER_130_1130 ();
 FILLCELL_X32 FILLER_130_1162 ();
 FILLCELL_X32 FILLER_130_1194 ();
 FILLCELL_X32 FILLER_130_1226 ();
 FILLCELL_X32 FILLER_130_1258 ();
 FILLCELL_X32 FILLER_130_1290 ();
 FILLCELL_X32 FILLER_130_1322 ();
 FILLCELL_X32 FILLER_130_1354 ();
 FILLCELL_X32 FILLER_130_1386 ();
 FILLCELL_X32 FILLER_130_1418 ();
 FILLCELL_X32 FILLER_130_1450 ();
 FILLCELL_X32 FILLER_130_1482 ();
 FILLCELL_X32 FILLER_130_1514 ();
 FILLCELL_X32 FILLER_130_1546 ();
 FILLCELL_X32 FILLER_130_1578 ();
 FILLCELL_X32 FILLER_130_1610 ();
 FILLCELL_X32 FILLER_130_1642 ();
 FILLCELL_X32 FILLER_130_1674 ();
 FILLCELL_X8 FILLER_130_1706 ();
 FILLCELL_X1 FILLER_130_1714 ();
 FILLCELL_X1 FILLER_130_1719 ();
 FILLCELL_X8 FILLER_130_1723 ();
 FILLCELL_X4 FILLER_130_1731 ();
 FILLCELL_X2 FILLER_130_1735 ();
 FILLCELL_X16 FILLER_130_1748 ();
 FILLCELL_X1 FILLER_130_1778 ();
 FILLCELL_X2 FILLER_130_1792 ();
 FILLCELL_X1 FILLER_131_1 ();
 FILLCELL_X1 FILLER_131_20 ();
 FILLCELL_X8 FILLER_131_30 ();
 FILLCELL_X4 FILLER_131_51 ();
 FILLCELL_X1 FILLER_131_55 ();
 FILLCELL_X32 FILLER_131_80 ();
 FILLCELL_X32 FILLER_131_112 ();
 FILLCELL_X32 FILLER_131_144 ();
 FILLCELL_X32 FILLER_131_176 ();
 FILLCELL_X32 FILLER_131_208 ();
 FILLCELL_X32 FILLER_131_240 ();
 FILLCELL_X32 FILLER_131_272 ();
 FILLCELL_X32 FILLER_131_304 ();
 FILLCELL_X32 FILLER_131_336 ();
 FILLCELL_X32 FILLER_131_368 ();
 FILLCELL_X32 FILLER_131_400 ();
 FILLCELL_X32 FILLER_131_432 ();
 FILLCELL_X32 FILLER_131_464 ();
 FILLCELL_X32 FILLER_131_496 ();
 FILLCELL_X32 FILLER_131_528 ();
 FILLCELL_X32 FILLER_131_560 ();
 FILLCELL_X32 FILLER_131_592 ();
 FILLCELL_X32 FILLER_131_624 ();
 FILLCELL_X32 FILLER_131_656 ();
 FILLCELL_X32 FILLER_131_688 ();
 FILLCELL_X32 FILLER_131_720 ();
 FILLCELL_X32 FILLER_131_752 ();
 FILLCELL_X4 FILLER_131_784 ();
 FILLCELL_X2 FILLER_131_788 ();
 FILLCELL_X2 FILLER_131_793 ();
 FILLCELL_X1 FILLER_131_795 ();
 FILLCELL_X1 FILLER_131_816 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X16 FILLER_131_897 ();
 FILLCELL_X4 FILLER_131_913 ();
 FILLCELL_X32 FILLER_131_930 ();
 FILLCELL_X32 FILLER_131_962 ();
 FILLCELL_X32 FILLER_131_994 ();
 FILLCELL_X32 FILLER_131_1026 ();
 FILLCELL_X32 FILLER_131_1058 ();
 FILLCELL_X32 FILLER_131_1090 ();
 FILLCELL_X32 FILLER_131_1122 ();
 FILLCELL_X32 FILLER_131_1154 ();
 FILLCELL_X32 FILLER_131_1186 ();
 FILLCELL_X32 FILLER_131_1218 ();
 FILLCELL_X8 FILLER_131_1250 ();
 FILLCELL_X4 FILLER_131_1258 ();
 FILLCELL_X1 FILLER_131_1262 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X32 FILLER_131_1584 ();
 FILLCELL_X32 FILLER_131_1616 ();
 FILLCELL_X32 FILLER_131_1648 ();
 FILLCELL_X32 FILLER_131_1680 ();
 FILLCELL_X32 FILLER_131_1712 ();
 FILLCELL_X16 FILLER_131_1744 ();
 FILLCELL_X4 FILLER_131_1760 ();
 FILLCELL_X2 FILLER_131_1771 ();
 FILLCELL_X1 FILLER_131_1773 ();
 FILLCELL_X2 FILLER_131_1780 ();
 FILLCELL_X2 FILLER_131_1791 ();
 FILLCELL_X1 FILLER_131_1796 ();
 FILLCELL_X2 FILLER_132_1 ();
 FILLCELL_X1 FILLER_132_6 ();
 FILLCELL_X4 FILLER_132_16 ();
 FILLCELL_X1 FILLER_132_20 ();
 FILLCELL_X1 FILLER_132_25 ();
 FILLCELL_X2 FILLER_132_30 ();
 FILLCELL_X32 FILLER_132_59 ();
 FILLCELL_X32 FILLER_132_91 ();
 FILLCELL_X32 FILLER_132_123 ();
 FILLCELL_X32 FILLER_132_155 ();
 FILLCELL_X32 FILLER_132_187 ();
 FILLCELL_X32 FILLER_132_219 ();
 FILLCELL_X32 FILLER_132_251 ();
 FILLCELL_X32 FILLER_132_283 ();
 FILLCELL_X32 FILLER_132_315 ();
 FILLCELL_X32 FILLER_132_347 ();
 FILLCELL_X32 FILLER_132_379 ();
 FILLCELL_X32 FILLER_132_411 ();
 FILLCELL_X32 FILLER_132_443 ();
 FILLCELL_X32 FILLER_132_475 ();
 FILLCELL_X32 FILLER_132_507 ();
 FILLCELL_X32 FILLER_132_539 ();
 FILLCELL_X32 FILLER_132_571 ();
 FILLCELL_X16 FILLER_132_603 ();
 FILLCELL_X8 FILLER_132_619 ();
 FILLCELL_X4 FILLER_132_627 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X16 FILLER_132_792 ();
 FILLCELL_X8 FILLER_132_808 ();
 FILLCELL_X1 FILLER_132_816 ();
 FILLCELL_X8 FILLER_132_820 ();
 FILLCELL_X2 FILLER_132_828 ();
 FILLCELL_X32 FILLER_132_855 ();
 FILLCELL_X32 FILLER_132_887 ();
 FILLCELL_X32 FILLER_132_919 ();
 FILLCELL_X32 FILLER_132_951 ();
 FILLCELL_X32 FILLER_132_983 ();
 FILLCELL_X32 FILLER_132_1015 ();
 FILLCELL_X32 FILLER_132_1047 ();
 FILLCELL_X32 FILLER_132_1079 ();
 FILLCELL_X32 FILLER_132_1111 ();
 FILLCELL_X32 FILLER_132_1143 ();
 FILLCELL_X32 FILLER_132_1175 ();
 FILLCELL_X32 FILLER_132_1207 ();
 FILLCELL_X32 FILLER_132_1239 ();
 FILLCELL_X32 FILLER_132_1271 ();
 FILLCELL_X32 FILLER_132_1303 ();
 FILLCELL_X32 FILLER_132_1335 ();
 FILLCELL_X32 FILLER_132_1367 ();
 FILLCELL_X32 FILLER_132_1399 ();
 FILLCELL_X32 FILLER_132_1431 ();
 FILLCELL_X32 FILLER_132_1463 ();
 FILLCELL_X32 FILLER_132_1495 ();
 FILLCELL_X32 FILLER_132_1527 ();
 FILLCELL_X32 FILLER_132_1559 ();
 FILLCELL_X32 FILLER_132_1591 ();
 FILLCELL_X32 FILLER_132_1623 ();
 FILLCELL_X32 FILLER_132_1655 ();
 FILLCELL_X32 FILLER_132_1687 ();
 FILLCELL_X16 FILLER_132_1719 ();
 FILLCELL_X2 FILLER_132_1735 ();
 FILLCELL_X4 FILLER_132_1739 ();
 FILLCELL_X2 FILLER_132_1743 ();
 FILLCELL_X32 FILLER_132_1755 ();
 FILLCELL_X2 FILLER_132_1787 ();
 FILLCELL_X4 FILLER_132_1792 ();
 FILLCELL_X1 FILLER_132_1796 ();
 FILLCELL_X16 FILLER_133_4 ();
 FILLCELL_X4 FILLER_133_20 ();
 FILLCELL_X2 FILLER_133_24 ();
 FILLCELL_X32 FILLER_133_32 ();
 FILLCELL_X32 FILLER_133_64 ();
 FILLCELL_X32 FILLER_133_96 ();
 FILLCELL_X32 FILLER_133_128 ();
 FILLCELL_X32 FILLER_133_160 ();
 FILLCELL_X32 FILLER_133_192 ();
 FILLCELL_X32 FILLER_133_224 ();
 FILLCELL_X32 FILLER_133_256 ();
 FILLCELL_X32 FILLER_133_288 ();
 FILLCELL_X32 FILLER_133_320 ();
 FILLCELL_X32 FILLER_133_352 ();
 FILLCELL_X32 FILLER_133_384 ();
 FILLCELL_X32 FILLER_133_416 ();
 FILLCELL_X32 FILLER_133_448 ();
 FILLCELL_X32 FILLER_133_480 ();
 FILLCELL_X32 FILLER_133_512 ();
 FILLCELL_X32 FILLER_133_544 ();
 FILLCELL_X32 FILLER_133_576 ();
 FILLCELL_X32 FILLER_133_608 ();
 FILLCELL_X32 FILLER_133_640 ();
 FILLCELL_X32 FILLER_133_672 ();
 FILLCELL_X32 FILLER_133_704 ();
 FILLCELL_X32 FILLER_133_736 ();
 FILLCELL_X32 FILLER_133_768 ();
 FILLCELL_X32 FILLER_133_800 ();
 FILLCELL_X32 FILLER_133_832 ();
 FILLCELL_X32 FILLER_133_864 ();
 FILLCELL_X32 FILLER_133_896 ();
 FILLCELL_X32 FILLER_133_928 ();
 FILLCELL_X32 FILLER_133_960 ();
 FILLCELL_X32 FILLER_133_992 ();
 FILLCELL_X32 FILLER_133_1024 ();
 FILLCELL_X32 FILLER_133_1056 ();
 FILLCELL_X32 FILLER_133_1088 ();
 FILLCELL_X32 FILLER_133_1120 ();
 FILLCELL_X32 FILLER_133_1152 ();
 FILLCELL_X32 FILLER_133_1184 ();
 FILLCELL_X32 FILLER_133_1216 ();
 FILLCELL_X8 FILLER_133_1248 ();
 FILLCELL_X4 FILLER_133_1256 ();
 FILLCELL_X2 FILLER_133_1260 ();
 FILLCELL_X1 FILLER_133_1262 ();
 FILLCELL_X32 FILLER_133_1264 ();
 FILLCELL_X32 FILLER_133_1296 ();
 FILLCELL_X32 FILLER_133_1328 ();
 FILLCELL_X32 FILLER_133_1360 ();
 FILLCELL_X32 FILLER_133_1392 ();
 FILLCELL_X32 FILLER_133_1424 ();
 FILLCELL_X32 FILLER_133_1456 ();
 FILLCELL_X32 FILLER_133_1488 ();
 FILLCELL_X32 FILLER_133_1520 ();
 FILLCELL_X32 FILLER_133_1552 ();
 FILLCELL_X32 FILLER_133_1584 ();
 FILLCELL_X32 FILLER_133_1616 ();
 FILLCELL_X32 FILLER_133_1648 ();
 FILLCELL_X32 FILLER_133_1680 ();
 FILLCELL_X16 FILLER_133_1712 ();
 FILLCELL_X1 FILLER_133_1728 ();
 FILLCELL_X8 FILLER_133_1739 ();
 FILLCELL_X2 FILLER_133_1747 ();
 FILLCELL_X8 FILLER_133_1751 ();
 FILLCELL_X4 FILLER_133_1759 ();
 FILLCELL_X1 FILLER_133_1763 ();
 FILLCELL_X4 FILLER_133_1793 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X32 FILLER_134_1016 ();
 FILLCELL_X32 FILLER_134_1048 ();
 FILLCELL_X32 FILLER_134_1080 ();
 FILLCELL_X32 FILLER_134_1112 ();
 FILLCELL_X32 FILLER_134_1144 ();
 FILLCELL_X32 FILLER_134_1176 ();
 FILLCELL_X32 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_134_1240 ();
 FILLCELL_X32 FILLER_134_1272 ();
 FILLCELL_X32 FILLER_134_1304 ();
 FILLCELL_X32 FILLER_134_1336 ();
 FILLCELL_X32 FILLER_134_1368 ();
 FILLCELL_X32 FILLER_134_1400 ();
 FILLCELL_X32 FILLER_134_1432 ();
 FILLCELL_X32 FILLER_134_1464 ();
 FILLCELL_X32 FILLER_134_1496 ();
 FILLCELL_X32 FILLER_134_1528 ();
 FILLCELL_X32 FILLER_134_1560 ();
 FILLCELL_X32 FILLER_134_1592 ();
 FILLCELL_X32 FILLER_134_1624 ();
 FILLCELL_X16 FILLER_134_1656 ();
 FILLCELL_X4 FILLER_134_1672 ();
 FILLCELL_X2 FILLER_134_1676 ();
 FILLCELL_X32 FILLER_134_1688 ();
 FILLCELL_X16 FILLER_134_1720 ();
 FILLCELL_X2 FILLER_134_1736 ();
 FILLCELL_X1 FILLER_134_1738 ();
 FILLCELL_X16 FILLER_134_1748 ();
 FILLCELL_X2 FILLER_134_1764 ();
 FILLCELL_X1 FILLER_134_1766 ();
 FILLCELL_X8 FILLER_134_1771 ();
 FILLCELL_X2 FILLER_134_1779 ();
 FILLCELL_X1 FILLER_134_1781 ();
 FILLCELL_X4 FILLER_134_1788 ();
 FILLCELL_X2 FILLER_134_1792 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X32 FILLER_135_993 ();
 FILLCELL_X32 FILLER_135_1025 ();
 FILLCELL_X32 FILLER_135_1057 ();
 FILLCELL_X32 FILLER_135_1089 ();
 FILLCELL_X32 FILLER_135_1121 ();
 FILLCELL_X32 FILLER_135_1153 ();
 FILLCELL_X32 FILLER_135_1185 ();
 FILLCELL_X32 FILLER_135_1217 ();
 FILLCELL_X8 FILLER_135_1249 ();
 FILLCELL_X4 FILLER_135_1257 ();
 FILLCELL_X2 FILLER_135_1261 ();
 FILLCELL_X32 FILLER_135_1264 ();
 FILLCELL_X32 FILLER_135_1296 ();
 FILLCELL_X32 FILLER_135_1328 ();
 FILLCELL_X32 FILLER_135_1360 ();
 FILLCELL_X32 FILLER_135_1392 ();
 FILLCELL_X32 FILLER_135_1424 ();
 FILLCELL_X32 FILLER_135_1456 ();
 FILLCELL_X32 FILLER_135_1488 ();
 FILLCELL_X32 FILLER_135_1520 ();
 FILLCELL_X32 FILLER_135_1552 ();
 FILLCELL_X32 FILLER_135_1584 ();
 FILLCELL_X32 FILLER_135_1616 ();
 FILLCELL_X32 FILLER_135_1648 ();
 FILLCELL_X32 FILLER_135_1680 ();
 FILLCELL_X32 FILLER_135_1712 ();
 FILLCELL_X16 FILLER_135_1744 ();
 FILLCELL_X8 FILLER_135_1760 ();
 FILLCELL_X2 FILLER_135_1768 ();
 FILLCELL_X2 FILLER_135_1772 ();
 FILLCELL_X1 FILLER_135_1774 ();
 FILLCELL_X2 FILLER_135_1794 ();
 FILLCELL_X1 FILLER_135_1796 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X32 FILLER_136_1016 ();
 FILLCELL_X32 FILLER_136_1048 ();
 FILLCELL_X32 FILLER_136_1080 ();
 FILLCELL_X32 FILLER_136_1112 ();
 FILLCELL_X32 FILLER_136_1144 ();
 FILLCELL_X32 FILLER_136_1176 ();
 FILLCELL_X32 FILLER_136_1208 ();
 FILLCELL_X32 FILLER_136_1240 ();
 FILLCELL_X32 FILLER_136_1272 ();
 FILLCELL_X32 FILLER_136_1304 ();
 FILLCELL_X32 FILLER_136_1336 ();
 FILLCELL_X32 FILLER_136_1368 ();
 FILLCELL_X32 FILLER_136_1400 ();
 FILLCELL_X32 FILLER_136_1432 ();
 FILLCELL_X32 FILLER_136_1464 ();
 FILLCELL_X32 FILLER_136_1496 ();
 FILLCELL_X32 FILLER_136_1528 ();
 FILLCELL_X32 FILLER_136_1560 ();
 FILLCELL_X32 FILLER_136_1592 ();
 FILLCELL_X32 FILLER_136_1624 ();
 FILLCELL_X32 FILLER_136_1656 ();
 FILLCELL_X32 FILLER_136_1688 ();
 FILLCELL_X2 FILLER_136_1720 ();
 FILLCELL_X1 FILLER_136_1722 ();
 FILLCELL_X1 FILLER_136_1750 ();
 FILLCELL_X2 FILLER_136_1760 ();
 FILLCELL_X1 FILLER_136_1766 ();
 FILLCELL_X2 FILLER_136_1771 ();
 FILLCELL_X2 FILLER_136_1783 ();
 FILLCELL_X1 FILLER_136_1785 ();
 FILLCELL_X8 FILLER_136_1789 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X32 FILLER_137_801 ();
 FILLCELL_X32 FILLER_137_833 ();
 FILLCELL_X32 FILLER_137_865 ();
 FILLCELL_X32 FILLER_137_897 ();
 FILLCELL_X32 FILLER_137_929 ();
 FILLCELL_X32 FILLER_137_961 ();
 FILLCELL_X32 FILLER_137_993 ();
 FILLCELL_X32 FILLER_137_1025 ();
 FILLCELL_X32 FILLER_137_1057 ();
 FILLCELL_X32 FILLER_137_1089 ();
 FILLCELL_X32 FILLER_137_1121 ();
 FILLCELL_X32 FILLER_137_1153 ();
 FILLCELL_X32 FILLER_137_1185 ();
 FILLCELL_X32 FILLER_137_1217 ();
 FILLCELL_X8 FILLER_137_1249 ();
 FILLCELL_X4 FILLER_137_1257 ();
 FILLCELL_X2 FILLER_137_1261 ();
 FILLCELL_X32 FILLER_137_1264 ();
 FILLCELL_X32 FILLER_137_1296 ();
 FILLCELL_X32 FILLER_137_1328 ();
 FILLCELL_X32 FILLER_137_1360 ();
 FILLCELL_X32 FILLER_137_1392 ();
 FILLCELL_X32 FILLER_137_1424 ();
 FILLCELL_X32 FILLER_137_1456 ();
 FILLCELL_X32 FILLER_137_1488 ();
 FILLCELL_X32 FILLER_137_1520 ();
 FILLCELL_X32 FILLER_137_1552 ();
 FILLCELL_X32 FILLER_137_1584 ();
 FILLCELL_X32 FILLER_137_1616 ();
 FILLCELL_X32 FILLER_137_1648 ();
 FILLCELL_X32 FILLER_137_1680 ();
 FILLCELL_X16 FILLER_137_1712 ();
 FILLCELL_X8 FILLER_137_1728 ();
 FILLCELL_X4 FILLER_137_1736 ();
 FILLCELL_X2 FILLER_137_1740 ();
 FILLCELL_X1 FILLER_137_1742 ();
 FILLCELL_X32 FILLER_137_1747 ();
 FILLCELL_X16 FILLER_137_1779 ();
 FILLCELL_X2 FILLER_137_1795 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X16 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X32 FILLER_138_824 ();
 FILLCELL_X32 FILLER_138_856 ();
 FILLCELL_X32 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_920 ();
 FILLCELL_X32 FILLER_138_952 ();
 FILLCELL_X32 FILLER_138_984 ();
 FILLCELL_X32 FILLER_138_1016 ();
 FILLCELL_X32 FILLER_138_1048 ();
 FILLCELL_X32 FILLER_138_1080 ();
 FILLCELL_X32 FILLER_138_1112 ();
 FILLCELL_X32 FILLER_138_1144 ();
 FILLCELL_X32 FILLER_138_1176 ();
 FILLCELL_X32 FILLER_138_1208 ();
 FILLCELL_X32 FILLER_138_1240 ();
 FILLCELL_X32 FILLER_138_1272 ();
 FILLCELL_X32 FILLER_138_1304 ();
 FILLCELL_X32 FILLER_138_1336 ();
 FILLCELL_X32 FILLER_138_1368 ();
 FILLCELL_X32 FILLER_138_1400 ();
 FILLCELL_X32 FILLER_138_1432 ();
 FILLCELL_X32 FILLER_138_1464 ();
 FILLCELL_X32 FILLER_138_1496 ();
 FILLCELL_X32 FILLER_138_1528 ();
 FILLCELL_X32 FILLER_138_1560 ();
 FILLCELL_X32 FILLER_138_1592 ();
 FILLCELL_X32 FILLER_138_1624 ();
 FILLCELL_X32 FILLER_138_1656 ();
 FILLCELL_X32 FILLER_138_1688 ();
 FILLCELL_X32 FILLER_138_1720 ();
 FILLCELL_X32 FILLER_138_1752 ();
 FILLCELL_X8 FILLER_138_1784 ();
 FILLCELL_X4 FILLER_138_1792 ();
 FILLCELL_X1 FILLER_138_1796 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X32 FILLER_139_577 ();
 FILLCELL_X32 FILLER_139_609 ();
 FILLCELL_X32 FILLER_139_641 ();
 FILLCELL_X32 FILLER_139_673 ();
 FILLCELL_X32 FILLER_139_705 ();
 FILLCELL_X32 FILLER_139_737 ();
 FILLCELL_X32 FILLER_139_769 ();
 FILLCELL_X32 FILLER_139_801 ();
 FILLCELL_X32 FILLER_139_833 ();
 FILLCELL_X32 FILLER_139_865 ();
 FILLCELL_X32 FILLER_139_897 ();
 FILLCELL_X32 FILLER_139_929 ();
 FILLCELL_X32 FILLER_139_961 ();
 FILLCELL_X32 FILLER_139_993 ();
 FILLCELL_X32 FILLER_139_1025 ();
 FILLCELL_X32 FILLER_139_1057 ();
 FILLCELL_X32 FILLER_139_1089 ();
 FILLCELL_X32 FILLER_139_1121 ();
 FILLCELL_X32 FILLER_139_1153 ();
 FILLCELL_X32 FILLER_139_1185 ();
 FILLCELL_X32 FILLER_139_1217 ();
 FILLCELL_X8 FILLER_139_1249 ();
 FILLCELL_X4 FILLER_139_1257 ();
 FILLCELL_X2 FILLER_139_1261 ();
 FILLCELL_X32 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1296 ();
 FILLCELL_X32 FILLER_139_1328 ();
 FILLCELL_X32 FILLER_139_1360 ();
 FILLCELL_X32 FILLER_139_1392 ();
 FILLCELL_X32 FILLER_139_1424 ();
 FILLCELL_X32 FILLER_139_1456 ();
 FILLCELL_X32 FILLER_139_1488 ();
 FILLCELL_X32 FILLER_139_1520 ();
 FILLCELL_X32 FILLER_139_1552 ();
 FILLCELL_X32 FILLER_139_1584 ();
 FILLCELL_X32 FILLER_139_1616 ();
 FILLCELL_X32 FILLER_139_1648 ();
 FILLCELL_X32 FILLER_139_1680 ();
 FILLCELL_X32 FILLER_139_1712 ();
 FILLCELL_X32 FILLER_139_1744 ();
 FILLCELL_X16 FILLER_139_1776 ();
 FILLCELL_X4 FILLER_139_1792 ();
 FILLCELL_X1 FILLER_139_1796 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X32 FILLER_140_1048 ();
 FILLCELL_X32 FILLER_140_1080 ();
 FILLCELL_X32 FILLER_140_1112 ();
 FILLCELL_X32 FILLER_140_1144 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X32 FILLER_140_1240 ();
 FILLCELL_X32 FILLER_140_1272 ();
 FILLCELL_X32 FILLER_140_1304 ();
 FILLCELL_X32 FILLER_140_1336 ();
 FILLCELL_X32 FILLER_140_1368 ();
 FILLCELL_X32 FILLER_140_1400 ();
 FILLCELL_X32 FILLER_140_1432 ();
 FILLCELL_X32 FILLER_140_1464 ();
 FILLCELL_X32 FILLER_140_1496 ();
 FILLCELL_X32 FILLER_140_1528 ();
 FILLCELL_X32 FILLER_140_1560 ();
 FILLCELL_X32 FILLER_140_1592 ();
 FILLCELL_X32 FILLER_140_1624 ();
 FILLCELL_X32 FILLER_140_1656 ();
 FILLCELL_X32 FILLER_140_1688 ();
 FILLCELL_X32 FILLER_140_1720 ();
 FILLCELL_X32 FILLER_140_1752 ();
 FILLCELL_X8 FILLER_140_1784 ();
 FILLCELL_X4 FILLER_140_1792 ();
 FILLCELL_X1 FILLER_140_1796 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X32 FILLER_141_993 ();
 FILLCELL_X32 FILLER_141_1025 ();
 FILLCELL_X32 FILLER_141_1057 ();
 FILLCELL_X32 FILLER_141_1089 ();
 FILLCELL_X32 FILLER_141_1121 ();
 FILLCELL_X32 FILLER_141_1153 ();
 FILLCELL_X32 FILLER_141_1185 ();
 FILLCELL_X32 FILLER_141_1217 ();
 FILLCELL_X8 FILLER_141_1249 ();
 FILLCELL_X4 FILLER_141_1257 ();
 FILLCELL_X2 FILLER_141_1261 ();
 FILLCELL_X32 FILLER_141_1264 ();
 FILLCELL_X32 FILLER_141_1296 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X32 FILLER_141_1360 ();
 FILLCELL_X32 FILLER_141_1392 ();
 FILLCELL_X32 FILLER_141_1424 ();
 FILLCELL_X32 FILLER_141_1456 ();
 FILLCELL_X32 FILLER_141_1488 ();
 FILLCELL_X32 FILLER_141_1520 ();
 FILLCELL_X32 FILLER_141_1552 ();
 FILLCELL_X32 FILLER_141_1584 ();
 FILLCELL_X32 FILLER_141_1616 ();
 FILLCELL_X32 FILLER_141_1648 ();
 FILLCELL_X32 FILLER_141_1680 ();
 FILLCELL_X32 FILLER_141_1712 ();
 FILLCELL_X32 FILLER_141_1744 ();
 FILLCELL_X16 FILLER_141_1776 ();
 FILLCELL_X4 FILLER_141_1792 ();
 FILLCELL_X1 FILLER_141_1796 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X32 FILLER_142_1112 ();
 FILLCELL_X32 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_142_1176 ();
 FILLCELL_X32 FILLER_142_1208 ();
 FILLCELL_X32 FILLER_142_1240 ();
 FILLCELL_X32 FILLER_142_1272 ();
 FILLCELL_X32 FILLER_142_1304 ();
 FILLCELL_X32 FILLER_142_1336 ();
 FILLCELL_X32 FILLER_142_1368 ();
 FILLCELL_X32 FILLER_142_1400 ();
 FILLCELL_X32 FILLER_142_1432 ();
 FILLCELL_X32 FILLER_142_1464 ();
 FILLCELL_X32 FILLER_142_1496 ();
 FILLCELL_X32 FILLER_142_1528 ();
 FILLCELL_X32 FILLER_142_1560 ();
 FILLCELL_X32 FILLER_142_1592 ();
 FILLCELL_X32 FILLER_142_1624 ();
 FILLCELL_X32 FILLER_142_1656 ();
 FILLCELL_X32 FILLER_142_1688 ();
 FILLCELL_X32 FILLER_142_1720 ();
 FILLCELL_X32 FILLER_142_1752 ();
 FILLCELL_X8 FILLER_142_1784 ();
 FILLCELL_X4 FILLER_142_1792 ();
 FILLCELL_X1 FILLER_142_1796 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X32 FILLER_143_1089 ();
 FILLCELL_X32 FILLER_143_1121 ();
 FILLCELL_X32 FILLER_143_1153 ();
 FILLCELL_X32 FILLER_143_1185 ();
 FILLCELL_X32 FILLER_143_1217 ();
 FILLCELL_X8 FILLER_143_1249 ();
 FILLCELL_X4 FILLER_143_1257 ();
 FILLCELL_X2 FILLER_143_1261 ();
 FILLCELL_X32 FILLER_143_1264 ();
 FILLCELL_X32 FILLER_143_1296 ();
 FILLCELL_X32 FILLER_143_1328 ();
 FILLCELL_X32 FILLER_143_1360 ();
 FILLCELL_X32 FILLER_143_1392 ();
 FILLCELL_X32 FILLER_143_1424 ();
 FILLCELL_X32 FILLER_143_1456 ();
 FILLCELL_X32 FILLER_143_1488 ();
 FILLCELL_X32 FILLER_143_1520 ();
 FILLCELL_X32 FILLER_143_1552 ();
 FILLCELL_X32 FILLER_143_1584 ();
 FILLCELL_X32 FILLER_143_1616 ();
 FILLCELL_X32 FILLER_143_1648 ();
 FILLCELL_X32 FILLER_143_1680 ();
 FILLCELL_X32 FILLER_143_1712 ();
 FILLCELL_X32 FILLER_143_1744 ();
 FILLCELL_X16 FILLER_143_1776 ();
 FILLCELL_X4 FILLER_143_1792 ();
 FILLCELL_X1 FILLER_143_1796 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X32 FILLER_144_1144 ();
 FILLCELL_X32 FILLER_144_1176 ();
 FILLCELL_X32 FILLER_144_1208 ();
 FILLCELL_X32 FILLER_144_1240 ();
 FILLCELL_X32 FILLER_144_1272 ();
 FILLCELL_X32 FILLER_144_1304 ();
 FILLCELL_X32 FILLER_144_1336 ();
 FILLCELL_X32 FILLER_144_1368 ();
 FILLCELL_X32 FILLER_144_1400 ();
 FILLCELL_X32 FILLER_144_1432 ();
 FILLCELL_X32 FILLER_144_1464 ();
 FILLCELL_X32 FILLER_144_1496 ();
 FILLCELL_X32 FILLER_144_1528 ();
 FILLCELL_X32 FILLER_144_1560 ();
 FILLCELL_X32 FILLER_144_1592 ();
 FILLCELL_X32 FILLER_144_1624 ();
 FILLCELL_X32 FILLER_144_1656 ();
 FILLCELL_X32 FILLER_144_1688 ();
 FILLCELL_X32 FILLER_144_1720 ();
 FILLCELL_X32 FILLER_144_1752 ();
 FILLCELL_X8 FILLER_144_1784 ();
 FILLCELL_X4 FILLER_144_1792 ();
 FILLCELL_X1 FILLER_144_1796 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X32 FILLER_145_1153 ();
 FILLCELL_X32 FILLER_145_1185 ();
 FILLCELL_X32 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1249 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X32 FILLER_145_1584 ();
 FILLCELL_X32 FILLER_145_1616 ();
 FILLCELL_X32 FILLER_145_1648 ();
 FILLCELL_X32 FILLER_145_1680 ();
 FILLCELL_X32 FILLER_145_1712 ();
 FILLCELL_X32 FILLER_145_1744 ();
 FILLCELL_X16 FILLER_145_1776 ();
 FILLCELL_X4 FILLER_145_1792 ();
 FILLCELL_X1 FILLER_145_1796 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X32 FILLER_146_1144 ();
 FILLCELL_X32 FILLER_146_1176 ();
 FILLCELL_X32 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_146_1240 ();
 FILLCELL_X32 FILLER_146_1272 ();
 FILLCELL_X32 FILLER_146_1304 ();
 FILLCELL_X32 FILLER_146_1336 ();
 FILLCELL_X32 FILLER_146_1368 ();
 FILLCELL_X32 FILLER_146_1400 ();
 FILLCELL_X32 FILLER_146_1432 ();
 FILLCELL_X32 FILLER_146_1464 ();
 FILLCELL_X32 FILLER_146_1496 ();
 FILLCELL_X32 FILLER_146_1528 ();
 FILLCELL_X32 FILLER_146_1560 ();
 FILLCELL_X32 FILLER_146_1592 ();
 FILLCELL_X32 FILLER_146_1624 ();
 FILLCELL_X32 FILLER_146_1656 ();
 FILLCELL_X32 FILLER_146_1688 ();
 FILLCELL_X32 FILLER_146_1720 ();
 FILLCELL_X32 FILLER_146_1752 ();
 FILLCELL_X8 FILLER_146_1784 ();
 FILLCELL_X4 FILLER_146_1792 ();
 FILLCELL_X1 FILLER_146_1796 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X32 FILLER_147_1185 ();
 FILLCELL_X32 FILLER_147_1217 ();
 FILLCELL_X8 FILLER_147_1249 ();
 FILLCELL_X4 FILLER_147_1257 ();
 FILLCELL_X2 FILLER_147_1261 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X32 FILLER_147_1584 ();
 FILLCELL_X32 FILLER_147_1616 ();
 FILLCELL_X32 FILLER_147_1648 ();
 FILLCELL_X32 FILLER_147_1680 ();
 FILLCELL_X32 FILLER_147_1712 ();
 FILLCELL_X32 FILLER_147_1744 ();
 FILLCELL_X16 FILLER_147_1776 ();
 FILLCELL_X4 FILLER_147_1792 ();
 FILLCELL_X1 FILLER_147_1796 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X32 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_148_1240 ();
 FILLCELL_X32 FILLER_148_1272 ();
 FILLCELL_X32 FILLER_148_1304 ();
 FILLCELL_X32 FILLER_148_1336 ();
 FILLCELL_X32 FILLER_148_1368 ();
 FILLCELL_X32 FILLER_148_1400 ();
 FILLCELL_X32 FILLER_148_1432 ();
 FILLCELL_X32 FILLER_148_1464 ();
 FILLCELL_X32 FILLER_148_1496 ();
 FILLCELL_X32 FILLER_148_1528 ();
 FILLCELL_X32 FILLER_148_1560 ();
 FILLCELL_X32 FILLER_148_1592 ();
 FILLCELL_X32 FILLER_148_1624 ();
 FILLCELL_X32 FILLER_148_1656 ();
 FILLCELL_X32 FILLER_148_1688 ();
 FILLCELL_X32 FILLER_148_1720 ();
 FILLCELL_X32 FILLER_148_1752 ();
 FILLCELL_X8 FILLER_148_1784 ();
 FILLCELL_X4 FILLER_148_1792 ();
 FILLCELL_X1 FILLER_148_1796 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X32 FILLER_149_1584 ();
 FILLCELL_X32 FILLER_149_1616 ();
 FILLCELL_X32 FILLER_149_1648 ();
 FILLCELL_X32 FILLER_149_1680 ();
 FILLCELL_X32 FILLER_149_1712 ();
 FILLCELL_X32 FILLER_149_1744 ();
 FILLCELL_X16 FILLER_149_1776 ();
 FILLCELL_X4 FILLER_149_1792 ();
 FILLCELL_X1 FILLER_149_1796 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X32 FILLER_150_1304 ();
 FILLCELL_X32 FILLER_150_1336 ();
 FILLCELL_X32 FILLER_150_1368 ();
 FILLCELL_X32 FILLER_150_1400 ();
 FILLCELL_X32 FILLER_150_1432 ();
 FILLCELL_X32 FILLER_150_1464 ();
 FILLCELL_X32 FILLER_150_1496 ();
 FILLCELL_X32 FILLER_150_1528 ();
 FILLCELL_X32 FILLER_150_1560 ();
 FILLCELL_X32 FILLER_150_1592 ();
 FILLCELL_X32 FILLER_150_1624 ();
 FILLCELL_X32 FILLER_150_1656 ();
 FILLCELL_X32 FILLER_150_1688 ();
 FILLCELL_X32 FILLER_150_1720 ();
 FILLCELL_X32 FILLER_150_1752 ();
 FILLCELL_X8 FILLER_150_1784 ();
 FILLCELL_X4 FILLER_150_1792 ();
 FILLCELL_X1 FILLER_150_1796 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X32 FILLER_151_1025 ();
 FILLCELL_X32 FILLER_151_1057 ();
 FILLCELL_X32 FILLER_151_1089 ();
 FILLCELL_X32 FILLER_151_1121 ();
 FILLCELL_X32 FILLER_151_1153 ();
 FILLCELL_X32 FILLER_151_1185 ();
 FILLCELL_X32 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1249 ();
 FILLCELL_X4 FILLER_151_1257 ();
 FILLCELL_X2 FILLER_151_1261 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X32 FILLER_151_1648 ();
 FILLCELL_X32 FILLER_151_1680 ();
 FILLCELL_X32 FILLER_151_1712 ();
 FILLCELL_X32 FILLER_151_1744 ();
 FILLCELL_X16 FILLER_151_1776 ();
 FILLCELL_X4 FILLER_151_1792 ();
 FILLCELL_X1 FILLER_151_1796 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X32 FILLER_152_1304 ();
 FILLCELL_X32 FILLER_152_1336 ();
 FILLCELL_X32 FILLER_152_1368 ();
 FILLCELL_X32 FILLER_152_1400 ();
 FILLCELL_X32 FILLER_152_1432 ();
 FILLCELL_X32 FILLER_152_1464 ();
 FILLCELL_X32 FILLER_152_1496 ();
 FILLCELL_X32 FILLER_152_1528 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X32 FILLER_152_1592 ();
 FILLCELL_X32 FILLER_152_1624 ();
 FILLCELL_X32 FILLER_152_1656 ();
 FILLCELL_X32 FILLER_152_1688 ();
 FILLCELL_X32 FILLER_152_1720 ();
 FILLCELL_X32 FILLER_152_1752 ();
 FILLCELL_X8 FILLER_152_1784 ();
 FILLCELL_X4 FILLER_152_1792 ();
 FILLCELL_X1 FILLER_152_1796 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X32 FILLER_153_961 ();
 FILLCELL_X32 FILLER_153_993 ();
 FILLCELL_X32 FILLER_153_1025 ();
 FILLCELL_X32 FILLER_153_1057 ();
 FILLCELL_X32 FILLER_153_1089 ();
 FILLCELL_X32 FILLER_153_1121 ();
 FILLCELL_X32 FILLER_153_1153 ();
 FILLCELL_X32 FILLER_153_1185 ();
 FILLCELL_X32 FILLER_153_1217 ();
 FILLCELL_X8 FILLER_153_1249 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X32 FILLER_153_1584 ();
 FILLCELL_X32 FILLER_153_1616 ();
 FILLCELL_X32 FILLER_153_1648 ();
 FILLCELL_X32 FILLER_153_1680 ();
 FILLCELL_X32 FILLER_153_1712 ();
 FILLCELL_X32 FILLER_153_1744 ();
 FILLCELL_X16 FILLER_153_1776 ();
 FILLCELL_X4 FILLER_153_1792 ();
 FILLCELL_X1 FILLER_153_1796 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X32 FILLER_154_1304 ();
 FILLCELL_X32 FILLER_154_1336 ();
 FILLCELL_X32 FILLER_154_1368 ();
 FILLCELL_X32 FILLER_154_1400 ();
 FILLCELL_X32 FILLER_154_1432 ();
 FILLCELL_X32 FILLER_154_1464 ();
 FILLCELL_X32 FILLER_154_1496 ();
 FILLCELL_X32 FILLER_154_1528 ();
 FILLCELL_X32 FILLER_154_1560 ();
 FILLCELL_X32 FILLER_154_1592 ();
 FILLCELL_X32 FILLER_154_1624 ();
 FILLCELL_X32 FILLER_154_1656 ();
 FILLCELL_X32 FILLER_154_1688 ();
 FILLCELL_X32 FILLER_154_1720 ();
 FILLCELL_X32 FILLER_154_1752 ();
 FILLCELL_X8 FILLER_154_1784 ();
 FILLCELL_X4 FILLER_154_1792 ();
 FILLCELL_X1 FILLER_154_1796 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X32 FILLER_155_929 ();
 FILLCELL_X32 FILLER_155_961 ();
 FILLCELL_X32 FILLER_155_993 ();
 FILLCELL_X32 FILLER_155_1025 ();
 FILLCELL_X32 FILLER_155_1057 ();
 FILLCELL_X32 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1121 ();
 FILLCELL_X32 FILLER_155_1153 ();
 FILLCELL_X32 FILLER_155_1185 ();
 FILLCELL_X32 FILLER_155_1217 ();
 FILLCELL_X8 FILLER_155_1249 ();
 FILLCELL_X4 FILLER_155_1257 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X32 FILLER_155_1584 ();
 FILLCELL_X32 FILLER_155_1616 ();
 FILLCELL_X32 FILLER_155_1648 ();
 FILLCELL_X32 FILLER_155_1680 ();
 FILLCELL_X32 FILLER_155_1712 ();
 FILLCELL_X32 FILLER_155_1744 ();
 FILLCELL_X16 FILLER_155_1776 ();
 FILLCELL_X4 FILLER_155_1792 ();
 FILLCELL_X1 FILLER_155_1796 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X32 FILLER_156_1080 ();
 FILLCELL_X32 FILLER_156_1112 ();
 FILLCELL_X32 FILLER_156_1144 ();
 FILLCELL_X32 FILLER_156_1176 ();
 FILLCELL_X32 FILLER_156_1208 ();
 FILLCELL_X32 FILLER_156_1240 ();
 FILLCELL_X32 FILLER_156_1272 ();
 FILLCELL_X32 FILLER_156_1304 ();
 FILLCELL_X32 FILLER_156_1336 ();
 FILLCELL_X32 FILLER_156_1368 ();
 FILLCELL_X32 FILLER_156_1400 ();
 FILLCELL_X32 FILLER_156_1432 ();
 FILLCELL_X32 FILLER_156_1464 ();
 FILLCELL_X32 FILLER_156_1496 ();
 FILLCELL_X32 FILLER_156_1528 ();
 FILLCELL_X32 FILLER_156_1560 ();
 FILLCELL_X32 FILLER_156_1592 ();
 FILLCELL_X32 FILLER_156_1624 ();
 FILLCELL_X32 FILLER_156_1656 ();
 FILLCELL_X32 FILLER_156_1688 ();
 FILLCELL_X32 FILLER_156_1720 ();
 FILLCELL_X32 FILLER_156_1752 ();
 FILLCELL_X8 FILLER_156_1784 ();
 FILLCELL_X4 FILLER_156_1792 ();
 FILLCELL_X1 FILLER_156_1796 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X32 FILLER_157_929 ();
 FILLCELL_X32 FILLER_157_961 ();
 FILLCELL_X32 FILLER_157_993 ();
 FILLCELL_X32 FILLER_157_1025 ();
 FILLCELL_X32 FILLER_157_1057 ();
 FILLCELL_X32 FILLER_157_1089 ();
 FILLCELL_X32 FILLER_157_1121 ();
 FILLCELL_X32 FILLER_157_1153 ();
 FILLCELL_X32 FILLER_157_1185 ();
 FILLCELL_X32 FILLER_157_1217 ();
 FILLCELL_X8 FILLER_157_1249 ();
 FILLCELL_X4 FILLER_157_1257 ();
 FILLCELL_X2 FILLER_157_1261 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X32 FILLER_157_1584 ();
 FILLCELL_X32 FILLER_157_1616 ();
 FILLCELL_X32 FILLER_157_1648 ();
 FILLCELL_X32 FILLER_157_1680 ();
 FILLCELL_X32 FILLER_157_1712 ();
 FILLCELL_X32 FILLER_157_1744 ();
 FILLCELL_X16 FILLER_157_1776 ();
 FILLCELL_X4 FILLER_157_1792 ();
 FILLCELL_X1 FILLER_157_1796 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X32 FILLER_158_1304 ();
 FILLCELL_X32 FILLER_158_1336 ();
 FILLCELL_X32 FILLER_158_1368 ();
 FILLCELL_X32 FILLER_158_1400 ();
 FILLCELL_X32 FILLER_158_1432 ();
 FILLCELL_X32 FILLER_158_1464 ();
 FILLCELL_X32 FILLER_158_1496 ();
 FILLCELL_X32 FILLER_158_1528 ();
 FILLCELL_X32 FILLER_158_1560 ();
 FILLCELL_X32 FILLER_158_1592 ();
 FILLCELL_X32 FILLER_158_1624 ();
 FILLCELL_X32 FILLER_158_1656 ();
 FILLCELL_X32 FILLER_158_1688 ();
 FILLCELL_X32 FILLER_158_1720 ();
 FILLCELL_X32 FILLER_158_1752 ();
 FILLCELL_X8 FILLER_158_1784 ();
 FILLCELL_X4 FILLER_158_1792 ();
 FILLCELL_X1 FILLER_158_1796 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X32 FILLER_159_929 ();
 FILLCELL_X32 FILLER_159_961 ();
 FILLCELL_X32 FILLER_159_993 ();
 FILLCELL_X32 FILLER_159_1025 ();
 FILLCELL_X32 FILLER_159_1057 ();
 FILLCELL_X32 FILLER_159_1089 ();
 FILLCELL_X32 FILLER_159_1121 ();
 FILLCELL_X32 FILLER_159_1153 ();
 FILLCELL_X32 FILLER_159_1185 ();
 FILLCELL_X32 FILLER_159_1217 ();
 FILLCELL_X8 FILLER_159_1249 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X32 FILLER_159_1584 ();
 FILLCELL_X32 FILLER_159_1616 ();
 FILLCELL_X32 FILLER_159_1648 ();
 FILLCELL_X32 FILLER_159_1680 ();
 FILLCELL_X32 FILLER_159_1712 ();
 FILLCELL_X32 FILLER_159_1744 ();
 FILLCELL_X16 FILLER_159_1776 ();
 FILLCELL_X4 FILLER_159_1792 ();
 FILLCELL_X1 FILLER_159_1796 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X32 FILLER_160_1304 ();
 FILLCELL_X32 FILLER_160_1336 ();
 FILLCELL_X32 FILLER_160_1368 ();
 FILLCELL_X32 FILLER_160_1400 ();
 FILLCELL_X32 FILLER_160_1432 ();
 FILLCELL_X32 FILLER_160_1464 ();
 FILLCELL_X32 FILLER_160_1496 ();
 FILLCELL_X32 FILLER_160_1528 ();
 FILLCELL_X32 FILLER_160_1560 ();
 FILLCELL_X32 FILLER_160_1592 ();
 FILLCELL_X32 FILLER_160_1624 ();
 FILLCELL_X32 FILLER_160_1656 ();
 FILLCELL_X32 FILLER_160_1688 ();
 FILLCELL_X32 FILLER_160_1720 ();
 FILLCELL_X32 FILLER_160_1752 ();
 FILLCELL_X8 FILLER_160_1784 ();
 FILLCELL_X4 FILLER_160_1792 ();
 FILLCELL_X1 FILLER_160_1796 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X32 FILLER_161_993 ();
 FILLCELL_X32 FILLER_161_1025 ();
 FILLCELL_X32 FILLER_161_1057 ();
 FILLCELL_X32 FILLER_161_1089 ();
 FILLCELL_X32 FILLER_161_1121 ();
 FILLCELL_X32 FILLER_161_1153 ();
 FILLCELL_X32 FILLER_161_1185 ();
 FILLCELL_X32 FILLER_161_1217 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X32 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1520 ();
 FILLCELL_X32 FILLER_161_1552 ();
 FILLCELL_X32 FILLER_161_1584 ();
 FILLCELL_X32 FILLER_161_1616 ();
 FILLCELL_X32 FILLER_161_1648 ();
 FILLCELL_X32 FILLER_161_1680 ();
 FILLCELL_X32 FILLER_161_1712 ();
 FILLCELL_X32 FILLER_161_1744 ();
 FILLCELL_X16 FILLER_161_1776 ();
 FILLCELL_X4 FILLER_161_1792 ();
 FILLCELL_X1 FILLER_161_1796 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X32 FILLER_162_1304 ();
 FILLCELL_X32 FILLER_162_1336 ();
 FILLCELL_X32 FILLER_162_1368 ();
 FILLCELL_X32 FILLER_162_1400 ();
 FILLCELL_X32 FILLER_162_1432 ();
 FILLCELL_X32 FILLER_162_1464 ();
 FILLCELL_X32 FILLER_162_1496 ();
 FILLCELL_X32 FILLER_162_1528 ();
 FILLCELL_X32 FILLER_162_1560 ();
 FILLCELL_X32 FILLER_162_1592 ();
 FILLCELL_X32 FILLER_162_1624 ();
 FILLCELL_X32 FILLER_162_1656 ();
 FILLCELL_X32 FILLER_162_1688 ();
 FILLCELL_X32 FILLER_162_1720 ();
 FILLCELL_X32 FILLER_162_1752 ();
 FILLCELL_X8 FILLER_162_1784 ();
 FILLCELL_X4 FILLER_162_1792 ();
 FILLCELL_X1 FILLER_162_1796 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X32 FILLER_163_961 ();
 FILLCELL_X32 FILLER_163_993 ();
 FILLCELL_X32 FILLER_163_1025 ();
 FILLCELL_X32 FILLER_163_1057 ();
 FILLCELL_X32 FILLER_163_1089 ();
 FILLCELL_X32 FILLER_163_1121 ();
 FILLCELL_X32 FILLER_163_1153 ();
 FILLCELL_X32 FILLER_163_1185 ();
 FILLCELL_X32 FILLER_163_1217 ();
 FILLCELL_X8 FILLER_163_1249 ();
 FILLCELL_X4 FILLER_163_1257 ();
 FILLCELL_X2 FILLER_163_1261 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X32 FILLER_163_1584 ();
 FILLCELL_X32 FILLER_163_1616 ();
 FILLCELL_X32 FILLER_163_1648 ();
 FILLCELL_X32 FILLER_163_1680 ();
 FILLCELL_X32 FILLER_163_1712 ();
 FILLCELL_X32 FILLER_163_1744 ();
 FILLCELL_X16 FILLER_163_1776 ();
 FILLCELL_X4 FILLER_163_1792 ();
 FILLCELL_X1 FILLER_163_1796 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X32 FILLER_164_1304 ();
 FILLCELL_X32 FILLER_164_1336 ();
 FILLCELL_X32 FILLER_164_1368 ();
 FILLCELL_X32 FILLER_164_1400 ();
 FILLCELL_X32 FILLER_164_1432 ();
 FILLCELL_X32 FILLER_164_1464 ();
 FILLCELL_X32 FILLER_164_1496 ();
 FILLCELL_X32 FILLER_164_1528 ();
 FILLCELL_X32 FILLER_164_1560 ();
 FILLCELL_X32 FILLER_164_1592 ();
 FILLCELL_X32 FILLER_164_1624 ();
 FILLCELL_X32 FILLER_164_1656 ();
 FILLCELL_X32 FILLER_164_1688 ();
 FILLCELL_X32 FILLER_164_1720 ();
 FILLCELL_X32 FILLER_164_1752 ();
 FILLCELL_X8 FILLER_164_1784 ();
 FILLCELL_X4 FILLER_164_1792 ();
 FILLCELL_X1 FILLER_164_1796 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X32 FILLER_165_993 ();
 FILLCELL_X32 FILLER_165_1025 ();
 FILLCELL_X32 FILLER_165_1057 ();
 FILLCELL_X32 FILLER_165_1089 ();
 FILLCELL_X32 FILLER_165_1121 ();
 FILLCELL_X32 FILLER_165_1153 ();
 FILLCELL_X32 FILLER_165_1185 ();
 FILLCELL_X32 FILLER_165_1217 ();
 FILLCELL_X8 FILLER_165_1249 ();
 FILLCELL_X4 FILLER_165_1257 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X32 FILLER_165_1584 ();
 FILLCELL_X32 FILLER_165_1616 ();
 FILLCELL_X32 FILLER_165_1648 ();
 FILLCELL_X32 FILLER_165_1680 ();
 FILLCELL_X32 FILLER_165_1712 ();
 FILLCELL_X32 FILLER_165_1744 ();
 FILLCELL_X16 FILLER_165_1776 ();
 FILLCELL_X4 FILLER_165_1792 ();
 FILLCELL_X1 FILLER_165_1796 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X32 FILLER_166_1048 ();
 FILLCELL_X32 FILLER_166_1080 ();
 FILLCELL_X32 FILLER_166_1112 ();
 FILLCELL_X32 FILLER_166_1144 ();
 FILLCELL_X32 FILLER_166_1176 ();
 FILLCELL_X32 FILLER_166_1208 ();
 FILLCELL_X32 FILLER_166_1240 ();
 FILLCELL_X32 FILLER_166_1272 ();
 FILLCELL_X32 FILLER_166_1304 ();
 FILLCELL_X32 FILLER_166_1336 ();
 FILLCELL_X32 FILLER_166_1368 ();
 FILLCELL_X32 FILLER_166_1400 ();
 FILLCELL_X32 FILLER_166_1432 ();
 FILLCELL_X32 FILLER_166_1464 ();
 FILLCELL_X32 FILLER_166_1496 ();
 FILLCELL_X32 FILLER_166_1528 ();
 FILLCELL_X32 FILLER_166_1560 ();
 FILLCELL_X32 FILLER_166_1592 ();
 FILLCELL_X32 FILLER_166_1624 ();
 FILLCELL_X32 FILLER_166_1656 ();
 FILLCELL_X32 FILLER_166_1688 ();
 FILLCELL_X32 FILLER_166_1720 ();
 FILLCELL_X32 FILLER_166_1752 ();
 FILLCELL_X8 FILLER_166_1784 ();
 FILLCELL_X4 FILLER_166_1792 ();
 FILLCELL_X1 FILLER_166_1796 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X32 FILLER_167_801 ();
 FILLCELL_X32 FILLER_167_833 ();
 FILLCELL_X32 FILLER_167_865 ();
 FILLCELL_X32 FILLER_167_897 ();
 FILLCELL_X32 FILLER_167_929 ();
 FILLCELL_X32 FILLER_167_961 ();
 FILLCELL_X32 FILLER_167_993 ();
 FILLCELL_X32 FILLER_167_1025 ();
 FILLCELL_X32 FILLER_167_1057 ();
 FILLCELL_X32 FILLER_167_1089 ();
 FILLCELL_X32 FILLER_167_1121 ();
 FILLCELL_X32 FILLER_167_1153 ();
 FILLCELL_X32 FILLER_167_1185 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X8 FILLER_167_1249 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X32 FILLER_167_1584 ();
 FILLCELL_X32 FILLER_167_1616 ();
 FILLCELL_X32 FILLER_167_1648 ();
 FILLCELL_X32 FILLER_167_1680 ();
 FILLCELL_X32 FILLER_167_1712 ();
 FILLCELL_X32 FILLER_167_1744 ();
 FILLCELL_X16 FILLER_167_1776 ();
 FILLCELL_X4 FILLER_167_1792 ();
 FILLCELL_X1 FILLER_167_1796 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X32 FILLER_168_1176 ();
 FILLCELL_X32 FILLER_168_1208 ();
 FILLCELL_X32 FILLER_168_1240 ();
 FILLCELL_X32 FILLER_168_1272 ();
 FILLCELL_X32 FILLER_168_1304 ();
 FILLCELL_X32 FILLER_168_1336 ();
 FILLCELL_X32 FILLER_168_1368 ();
 FILLCELL_X32 FILLER_168_1400 ();
 FILLCELL_X32 FILLER_168_1432 ();
 FILLCELL_X32 FILLER_168_1464 ();
 FILLCELL_X32 FILLER_168_1496 ();
 FILLCELL_X32 FILLER_168_1528 ();
 FILLCELL_X32 FILLER_168_1560 ();
 FILLCELL_X32 FILLER_168_1592 ();
 FILLCELL_X32 FILLER_168_1624 ();
 FILLCELL_X32 FILLER_168_1656 ();
 FILLCELL_X32 FILLER_168_1688 ();
 FILLCELL_X32 FILLER_168_1720 ();
 FILLCELL_X32 FILLER_168_1752 ();
 FILLCELL_X8 FILLER_168_1784 ();
 FILLCELL_X4 FILLER_168_1792 ();
 FILLCELL_X1 FILLER_168_1796 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X32 FILLER_169_577 ();
 FILLCELL_X32 FILLER_169_609 ();
 FILLCELL_X32 FILLER_169_641 ();
 FILLCELL_X32 FILLER_169_673 ();
 FILLCELL_X32 FILLER_169_705 ();
 FILLCELL_X32 FILLER_169_737 ();
 FILLCELL_X32 FILLER_169_769 ();
 FILLCELL_X32 FILLER_169_801 ();
 FILLCELL_X32 FILLER_169_833 ();
 FILLCELL_X32 FILLER_169_865 ();
 FILLCELL_X32 FILLER_169_897 ();
 FILLCELL_X32 FILLER_169_929 ();
 FILLCELL_X32 FILLER_169_961 ();
 FILLCELL_X32 FILLER_169_993 ();
 FILLCELL_X32 FILLER_169_1025 ();
 FILLCELL_X32 FILLER_169_1057 ();
 FILLCELL_X32 FILLER_169_1089 ();
 FILLCELL_X32 FILLER_169_1121 ();
 FILLCELL_X32 FILLER_169_1153 ();
 FILLCELL_X32 FILLER_169_1185 ();
 FILLCELL_X32 FILLER_169_1217 ();
 FILLCELL_X8 FILLER_169_1249 ();
 FILLCELL_X4 FILLER_169_1257 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X32 FILLER_169_1584 ();
 FILLCELL_X32 FILLER_169_1616 ();
 FILLCELL_X32 FILLER_169_1648 ();
 FILLCELL_X32 FILLER_169_1680 ();
 FILLCELL_X32 FILLER_169_1712 ();
 FILLCELL_X32 FILLER_169_1744 ();
 FILLCELL_X16 FILLER_169_1776 ();
 FILLCELL_X4 FILLER_169_1792 ();
 FILLCELL_X1 FILLER_169_1796 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X32 FILLER_170_1048 ();
 FILLCELL_X32 FILLER_170_1080 ();
 FILLCELL_X32 FILLER_170_1112 ();
 FILLCELL_X32 FILLER_170_1144 ();
 FILLCELL_X32 FILLER_170_1176 ();
 FILLCELL_X32 FILLER_170_1208 ();
 FILLCELL_X32 FILLER_170_1240 ();
 FILLCELL_X32 FILLER_170_1272 ();
 FILLCELL_X32 FILLER_170_1304 ();
 FILLCELL_X32 FILLER_170_1336 ();
 FILLCELL_X32 FILLER_170_1368 ();
 FILLCELL_X32 FILLER_170_1400 ();
 FILLCELL_X32 FILLER_170_1432 ();
 FILLCELL_X32 FILLER_170_1464 ();
 FILLCELL_X32 FILLER_170_1496 ();
 FILLCELL_X32 FILLER_170_1528 ();
 FILLCELL_X32 FILLER_170_1560 ();
 FILLCELL_X32 FILLER_170_1592 ();
 FILLCELL_X32 FILLER_170_1624 ();
 FILLCELL_X32 FILLER_170_1656 ();
 FILLCELL_X32 FILLER_170_1688 ();
 FILLCELL_X32 FILLER_170_1720 ();
 FILLCELL_X32 FILLER_170_1752 ();
 FILLCELL_X8 FILLER_170_1784 ();
 FILLCELL_X4 FILLER_170_1792 ();
 FILLCELL_X1 FILLER_170_1796 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X32 FILLER_171_353 ();
 FILLCELL_X32 FILLER_171_385 ();
 FILLCELL_X32 FILLER_171_417 ();
 FILLCELL_X32 FILLER_171_449 ();
 FILLCELL_X32 FILLER_171_481 ();
 FILLCELL_X32 FILLER_171_513 ();
 FILLCELL_X32 FILLER_171_545 ();
 FILLCELL_X32 FILLER_171_577 ();
 FILLCELL_X32 FILLER_171_609 ();
 FILLCELL_X32 FILLER_171_641 ();
 FILLCELL_X32 FILLER_171_673 ();
 FILLCELL_X32 FILLER_171_705 ();
 FILLCELL_X32 FILLER_171_737 ();
 FILLCELL_X32 FILLER_171_769 ();
 FILLCELL_X32 FILLER_171_801 ();
 FILLCELL_X32 FILLER_171_833 ();
 FILLCELL_X32 FILLER_171_865 ();
 FILLCELL_X32 FILLER_171_897 ();
 FILLCELL_X32 FILLER_171_929 ();
 FILLCELL_X32 FILLER_171_961 ();
 FILLCELL_X32 FILLER_171_993 ();
 FILLCELL_X32 FILLER_171_1025 ();
 FILLCELL_X32 FILLER_171_1057 ();
 FILLCELL_X32 FILLER_171_1089 ();
 FILLCELL_X32 FILLER_171_1121 ();
 FILLCELL_X32 FILLER_171_1153 ();
 FILLCELL_X32 FILLER_171_1185 ();
 FILLCELL_X32 FILLER_171_1217 ();
 FILLCELL_X8 FILLER_171_1249 ();
 FILLCELL_X4 FILLER_171_1257 ();
 FILLCELL_X2 FILLER_171_1261 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X32 FILLER_171_1584 ();
 FILLCELL_X32 FILLER_171_1616 ();
 FILLCELL_X32 FILLER_171_1648 ();
 FILLCELL_X32 FILLER_171_1680 ();
 FILLCELL_X32 FILLER_171_1712 ();
 FILLCELL_X32 FILLER_171_1744 ();
 FILLCELL_X16 FILLER_171_1776 ();
 FILLCELL_X4 FILLER_171_1792 ();
 FILLCELL_X1 FILLER_171_1796 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X32 FILLER_172_1080 ();
 FILLCELL_X32 FILLER_172_1112 ();
 FILLCELL_X32 FILLER_172_1144 ();
 FILLCELL_X32 FILLER_172_1176 ();
 FILLCELL_X32 FILLER_172_1208 ();
 FILLCELL_X32 FILLER_172_1240 ();
 FILLCELL_X32 FILLER_172_1272 ();
 FILLCELL_X32 FILLER_172_1304 ();
 FILLCELL_X32 FILLER_172_1336 ();
 FILLCELL_X32 FILLER_172_1368 ();
 FILLCELL_X32 FILLER_172_1400 ();
 FILLCELL_X32 FILLER_172_1432 ();
 FILLCELL_X32 FILLER_172_1464 ();
 FILLCELL_X32 FILLER_172_1496 ();
 FILLCELL_X32 FILLER_172_1528 ();
 FILLCELL_X32 FILLER_172_1560 ();
 FILLCELL_X32 FILLER_172_1592 ();
 FILLCELL_X32 FILLER_172_1624 ();
 FILLCELL_X32 FILLER_172_1656 ();
 FILLCELL_X32 FILLER_172_1688 ();
 FILLCELL_X32 FILLER_172_1720 ();
 FILLCELL_X32 FILLER_172_1752 ();
 FILLCELL_X8 FILLER_172_1784 ();
 FILLCELL_X4 FILLER_172_1792 ();
 FILLCELL_X1 FILLER_172_1796 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X32 FILLER_173_1089 ();
 FILLCELL_X32 FILLER_173_1121 ();
 FILLCELL_X32 FILLER_173_1153 ();
 FILLCELL_X32 FILLER_173_1185 ();
 FILLCELL_X32 FILLER_173_1217 ();
 FILLCELL_X8 FILLER_173_1249 ();
 FILLCELL_X4 FILLER_173_1257 ();
 FILLCELL_X2 FILLER_173_1261 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X32 FILLER_173_1584 ();
 FILLCELL_X32 FILLER_173_1616 ();
 FILLCELL_X32 FILLER_173_1648 ();
 FILLCELL_X32 FILLER_173_1680 ();
 FILLCELL_X32 FILLER_173_1712 ();
 FILLCELL_X32 FILLER_173_1744 ();
 FILLCELL_X16 FILLER_173_1776 ();
 FILLCELL_X4 FILLER_173_1792 ();
 FILLCELL_X1 FILLER_173_1796 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X32 FILLER_174_1304 ();
 FILLCELL_X32 FILLER_174_1336 ();
 FILLCELL_X32 FILLER_174_1368 ();
 FILLCELL_X32 FILLER_174_1400 ();
 FILLCELL_X32 FILLER_174_1432 ();
 FILLCELL_X32 FILLER_174_1464 ();
 FILLCELL_X32 FILLER_174_1496 ();
 FILLCELL_X32 FILLER_174_1528 ();
 FILLCELL_X32 FILLER_174_1560 ();
 FILLCELL_X32 FILLER_174_1592 ();
 FILLCELL_X32 FILLER_174_1624 ();
 FILLCELL_X32 FILLER_174_1656 ();
 FILLCELL_X32 FILLER_174_1688 ();
 FILLCELL_X32 FILLER_174_1720 ();
 FILLCELL_X32 FILLER_174_1752 ();
 FILLCELL_X8 FILLER_174_1784 ();
 FILLCELL_X4 FILLER_174_1792 ();
 FILLCELL_X1 FILLER_174_1796 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X32 FILLER_175_385 ();
 FILLCELL_X32 FILLER_175_417 ();
 FILLCELL_X32 FILLER_175_449 ();
 FILLCELL_X32 FILLER_175_481 ();
 FILLCELL_X32 FILLER_175_513 ();
 FILLCELL_X32 FILLER_175_545 ();
 FILLCELL_X32 FILLER_175_577 ();
 FILLCELL_X32 FILLER_175_609 ();
 FILLCELL_X32 FILLER_175_641 ();
 FILLCELL_X32 FILLER_175_673 ();
 FILLCELL_X32 FILLER_175_705 ();
 FILLCELL_X32 FILLER_175_737 ();
 FILLCELL_X32 FILLER_175_769 ();
 FILLCELL_X32 FILLER_175_801 ();
 FILLCELL_X32 FILLER_175_833 ();
 FILLCELL_X32 FILLER_175_865 ();
 FILLCELL_X32 FILLER_175_897 ();
 FILLCELL_X32 FILLER_175_929 ();
 FILLCELL_X32 FILLER_175_961 ();
 FILLCELL_X32 FILLER_175_993 ();
 FILLCELL_X32 FILLER_175_1025 ();
 FILLCELL_X32 FILLER_175_1057 ();
 FILLCELL_X32 FILLER_175_1089 ();
 FILLCELL_X32 FILLER_175_1121 ();
 FILLCELL_X32 FILLER_175_1153 ();
 FILLCELL_X32 FILLER_175_1185 ();
 FILLCELL_X32 FILLER_175_1217 ();
 FILLCELL_X8 FILLER_175_1249 ();
 FILLCELL_X4 FILLER_175_1257 ();
 FILLCELL_X2 FILLER_175_1261 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X32 FILLER_175_1584 ();
 FILLCELL_X32 FILLER_175_1616 ();
 FILLCELL_X32 FILLER_175_1648 ();
 FILLCELL_X32 FILLER_175_1680 ();
 FILLCELL_X32 FILLER_175_1712 ();
 FILLCELL_X32 FILLER_175_1744 ();
 FILLCELL_X16 FILLER_175_1776 ();
 FILLCELL_X4 FILLER_175_1792 ();
 FILLCELL_X1 FILLER_175_1796 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X32 FILLER_176_353 ();
 FILLCELL_X32 FILLER_176_385 ();
 FILLCELL_X32 FILLER_176_417 ();
 FILLCELL_X32 FILLER_176_449 ();
 FILLCELL_X32 FILLER_176_481 ();
 FILLCELL_X32 FILLER_176_513 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X32 FILLER_176_577 ();
 FILLCELL_X16 FILLER_176_609 ();
 FILLCELL_X4 FILLER_176_625 ();
 FILLCELL_X2 FILLER_176_629 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X32 FILLER_176_1112 ();
 FILLCELL_X32 FILLER_176_1144 ();
 FILLCELL_X32 FILLER_176_1176 ();
 FILLCELL_X32 FILLER_176_1208 ();
 FILLCELL_X32 FILLER_176_1240 ();
 FILLCELL_X32 FILLER_176_1272 ();
 FILLCELL_X32 FILLER_176_1304 ();
 FILLCELL_X32 FILLER_176_1336 ();
 FILLCELL_X32 FILLER_176_1368 ();
 FILLCELL_X32 FILLER_176_1400 ();
 FILLCELL_X32 FILLER_176_1432 ();
 FILLCELL_X32 FILLER_176_1464 ();
 FILLCELL_X32 FILLER_176_1496 ();
 FILLCELL_X32 FILLER_176_1528 ();
 FILLCELL_X32 FILLER_176_1560 ();
 FILLCELL_X32 FILLER_176_1592 ();
 FILLCELL_X32 FILLER_176_1624 ();
 FILLCELL_X32 FILLER_176_1656 ();
 FILLCELL_X32 FILLER_176_1688 ();
 FILLCELL_X32 FILLER_176_1720 ();
 FILLCELL_X32 FILLER_176_1752 ();
 FILLCELL_X8 FILLER_176_1784 ();
 FILLCELL_X4 FILLER_176_1792 ();
 FILLCELL_X1 FILLER_176_1796 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X32 FILLER_177_1089 ();
 FILLCELL_X32 FILLER_177_1121 ();
 FILLCELL_X32 FILLER_177_1153 ();
 FILLCELL_X32 FILLER_177_1185 ();
 FILLCELL_X32 FILLER_177_1217 ();
 FILLCELL_X8 FILLER_177_1249 ();
 FILLCELL_X4 FILLER_177_1257 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X32 FILLER_177_1584 ();
 FILLCELL_X32 FILLER_177_1616 ();
 FILLCELL_X32 FILLER_177_1648 ();
 FILLCELL_X32 FILLER_177_1680 ();
 FILLCELL_X32 FILLER_177_1712 ();
 FILLCELL_X32 FILLER_177_1744 ();
 FILLCELL_X16 FILLER_177_1776 ();
 FILLCELL_X4 FILLER_177_1792 ();
 FILLCELL_X1 FILLER_177_1796 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X32 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1144 ();
 FILLCELL_X32 FILLER_178_1176 ();
 FILLCELL_X32 FILLER_178_1208 ();
 FILLCELL_X32 FILLER_178_1240 ();
 FILLCELL_X32 FILLER_178_1272 ();
 FILLCELL_X32 FILLER_178_1304 ();
 FILLCELL_X32 FILLER_178_1336 ();
 FILLCELL_X32 FILLER_178_1368 ();
 FILLCELL_X32 FILLER_178_1400 ();
 FILLCELL_X32 FILLER_178_1432 ();
 FILLCELL_X32 FILLER_178_1464 ();
 FILLCELL_X32 FILLER_178_1496 ();
 FILLCELL_X32 FILLER_178_1528 ();
 FILLCELL_X32 FILLER_178_1560 ();
 FILLCELL_X32 FILLER_178_1592 ();
 FILLCELL_X32 FILLER_178_1624 ();
 FILLCELL_X32 FILLER_178_1656 ();
 FILLCELL_X32 FILLER_178_1688 ();
 FILLCELL_X32 FILLER_178_1720 ();
 FILLCELL_X32 FILLER_178_1752 ();
 FILLCELL_X8 FILLER_178_1784 ();
 FILLCELL_X4 FILLER_178_1792 ();
 FILLCELL_X1 FILLER_178_1796 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X32 FILLER_179_1089 ();
 FILLCELL_X32 FILLER_179_1121 ();
 FILLCELL_X32 FILLER_179_1153 ();
 FILLCELL_X32 FILLER_179_1185 ();
 FILLCELL_X32 FILLER_179_1217 ();
 FILLCELL_X8 FILLER_179_1249 ();
 FILLCELL_X4 FILLER_179_1257 ();
 FILLCELL_X2 FILLER_179_1261 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X32 FILLER_179_1584 ();
 FILLCELL_X32 FILLER_179_1616 ();
 FILLCELL_X32 FILLER_179_1648 ();
 FILLCELL_X32 FILLER_179_1680 ();
 FILLCELL_X32 FILLER_179_1712 ();
 FILLCELL_X32 FILLER_179_1744 ();
 FILLCELL_X16 FILLER_179_1776 ();
 FILLCELL_X4 FILLER_179_1792 ();
 FILLCELL_X1 FILLER_179_1796 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X32 FILLER_180_353 ();
 FILLCELL_X32 FILLER_180_385 ();
 FILLCELL_X32 FILLER_180_417 ();
 FILLCELL_X32 FILLER_180_449 ();
 FILLCELL_X32 FILLER_180_481 ();
 FILLCELL_X32 FILLER_180_513 ();
 FILLCELL_X32 FILLER_180_545 ();
 FILLCELL_X32 FILLER_180_577 ();
 FILLCELL_X16 FILLER_180_609 ();
 FILLCELL_X4 FILLER_180_625 ();
 FILLCELL_X2 FILLER_180_629 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X32 FILLER_180_1080 ();
 FILLCELL_X32 FILLER_180_1112 ();
 FILLCELL_X32 FILLER_180_1144 ();
 FILLCELL_X32 FILLER_180_1176 ();
 FILLCELL_X32 FILLER_180_1208 ();
 FILLCELL_X32 FILLER_180_1240 ();
 FILLCELL_X32 FILLER_180_1272 ();
 FILLCELL_X32 FILLER_180_1304 ();
 FILLCELL_X32 FILLER_180_1336 ();
 FILLCELL_X32 FILLER_180_1368 ();
 FILLCELL_X32 FILLER_180_1400 ();
 FILLCELL_X32 FILLER_180_1432 ();
 FILLCELL_X32 FILLER_180_1464 ();
 FILLCELL_X32 FILLER_180_1496 ();
 FILLCELL_X32 FILLER_180_1528 ();
 FILLCELL_X32 FILLER_180_1560 ();
 FILLCELL_X32 FILLER_180_1592 ();
 FILLCELL_X32 FILLER_180_1624 ();
 FILLCELL_X32 FILLER_180_1656 ();
 FILLCELL_X32 FILLER_180_1688 ();
 FILLCELL_X32 FILLER_180_1720 ();
 FILLCELL_X32 FILLER_180_1752 ();
 FILLCELL_X8 FILLER_180_1784 ();
 FILLCELL_X4 FILLER_180_1792 ();
 FILLCELL_X1 FILLER_180_1796 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X32 FILLER_181_1089 ();
 FILLCELL_X32 FILLER_181_1121 ();
 FILLCELL_X32 FILLER_181_1153 ();
 FILLCELL_X32 FILLER_181_1185 ();
 FILLCELL_X32 FILLER_181_1217 ();
 FILLCELL_X8 FILLER_181_1249 ();
 FILLCELL_X4 FILLER_181_1257 ();
 FILLCELL_X2 FILLER_181_1261 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X32 FILLER_181_1584 ();
 FILLCELL_X32 FILLER_181_1616 ();
 FILLCELL_X32 FILLER_181_1648 ();
 FILLCELL_X32 FILLER_181_1680 ();
 FILLCELL_X32 FILLER_181_1712 ();
 FILLCELL_X32 FILLER_181_1744 ();
 FILLCELL_X16 FILLER_181_1776 ();
 FILLCELL_X4 FILLER_181_1792 ();
 FILLCELL_X1 FILLER_181_1796 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X32 FILLER_182_1080 ();
 FILLCELL_X32 FILLER_182_1112 ();
 FILLCELL_X32 FILLER_182_1144 ();
 FILLCELL_X32 FILLER_182_1176 ();
 FILLCELL_X32 FILLER_182_1208 ();
 FILLCELL_X32 FILLER_182_1240 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X32 FILLER_182_1400 ();
 FILLCELL_X32 FILLER_182_1432 ();
 FILLCELL_X32 FILLER_182_1464 ();
 FILLCELL_X32 FILLER_182_1496 ();
 FILLCELL_X32 FILLER_182_1528 ();
 FILLCELL_X32 FILLER_182_1560 ();
 FILLCELL_X32 FILLER_182_1592 ();
 FILLCELL_X32 FILLER_182_1624 ();
 FILLCELL_X32 FILLER_182_1656 ();
 FILLCELL_X32 FILLER_182_1688 ();
 FILLCELL_X32 FILLER_182_1720 ();
 FILLCELL_X32 FILLER_182_1752 ();
 FILLCELL_X8 FILLER_182_1784 ();
 FILLCELL_X4 FILLER_182_1792 ();
 FILLCELL_X1 FILLER_182_1796 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X32 FILLER_183_1089 ();
 FILLCELL_X32 FILLER_183_1121 ();
 FILLCELL_X32 FILLER_183_1153 ();
 FILLCELL_X32 FILLER_183_1185 ();
 FILLCELL_X32 FILLER_183_1217 ();
 FILLCELL_X8 FILLER_183_1249 ();
 FILLCELL_X4 FILLER_183_1257 ();
 FILLCELL_X2 FILLER_183_1261 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X32 FILLER_183_1584 ();
 FILLCELL_X32 FILLER_183_1616 ();
 FILLCELL_X32 FILLER_183_1648 ();
 FILLCELL_X32 FILLER_183_1680 ();
 FILLCELL_X32 FILLER_183_1712 ();
 FILLCELL_X32 FILLER_183_1744 ();
 FILLCELL_X16 FILLER_183_1776 ();
 FILLCELL_X4 FILLER_183_1792 ();
 FILLCELL_X1 FILLER_183_1796 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X32 FILLER_184_1144 ();
 FILLCELL_X32 FILLER_184_1176 ();
 FILLCELL_X32 FILLER_184_1208 ();
 FILLCELL_X32 FILLER_184_1240 ();
 FILLCELL_X32 FILLER_184_1272 ();
 FILLCELL_X32 FILLER_184_1304 ();
 FILLCELL_X32 FILLER_184_1336 ();
 FILLCELL_X32 FILLER_184_1368 ();
 FILLCELL_X32 FILLER_184_1400 ();
 FILLCELL_X32 FILLER_184_1432 ();
 FILLCELL_X32 FILLER_184_1464 ();
 FILLCELL_X32 FILLER_184_1496 ();
 FILLCELL_X32 FILLER_184_1528 ();
 FILLCELL_X32 FILLER_184_1560 ();
 FILLCELL_X32 FILLER_184_1592 ();
 FILLCELL_X32 FILLER_184_1624 ();
 FILLCELL_X32 FILLER_184_1656 ();
 FILLCELL_X32 FILLER_184_1688 ();
 FILLCELL_X32 FILLER_184_1720 ();
 FILLCELL_X32 FILLER_184_1752 ();
 FILLCELL_X8 FILLER_184_1784 ();
 FILLCELL_X4 FILLER_184_1792 ();
 FILLCELL_X1 FILLER_184_1796 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X32 FILLER_185_1185 ();
 FILLCELL_X32 FILLER_185_1217 ();
 FILLCELL_X8 FILLER_185_1249 ();
 FILLCELL_X4 FILLER_185_1257 ();
 FILLCELL_X2 FILLER_185_1261 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X32 FILLER_185_1584 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X32 FILLER_185_1648 ();
 FILLCELL_X32 FILLER_185_1680 ();
 FILLCELL_X32 FILLER_185_1712 ();
 FILLCELL_X32 FILLER_185_1744 ();
 FILLCELL_X16 FILLER_185_1776 ();
 FILLCELL_X4 FILLER_185_1792 ();
 FILLCELL_X1 FILLER_185_1796 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X32 FILLER_186_1240 ();
 FILLCELL_X32 FILLER_186_1272 ();
 FILLCELL_X32 FILLER_186_1304 ();
 FILLCELL_X32 FILLER_186_1336 ();
 FILLCELL_X32 FILLER_186_1368 ();
 FILLCELL_X32 FILLER_186_1400 ();
 FILLCELL_X32 FILLER_186_1432 ();
 FILLCELL_X32 FILLER_186_1464 ();
 FILLCELL_X32 FILLER_186_1496 ();
 FILLCELL_X32 FILLER_186_1528 ();
 FILLCELL_X32 FILLER_186_1560 ();
 FILLCELL_X32 FILLER_186_1592 ();
 FILLCELL_X32 FILLER_186_1624 ();
 FILLCELL_X32 FILLER_186_1656 ();
 FILLCELL_X32 FILLER_186_1688 ();
 FILLCELL_X32 FILLER_186_1720 ();
 FILLCELL_X32 FILLER_186_1752 ();
 FILLCELL_X8 FILLER_186_1784 ();
 FILLCELL_X4 FILLER_186_1792 ();
 FILLCELL_X1 FILLER_186_1796 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X32 FILLER_187_1217 ();
 FILLCELL_X8 FILLER_187_1249 ();
 FILLCELL_X4 FILLER_187_1257 ();
 FILLCELL_X2 FILLER_187_1261 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X32 FILLER_187_1584 ();
 FILLCELL_X32 FILLER_187_1616 ();
 FILLCELL_X32 FILLER_187_1648 ();
 FILLCELL_X32 FILLER_187_1680 ();
 FILLCELL_X32 FILLER_187_1712 ();
 FILLCELL_X32 FILLER_187_1744 ();
 FILLCELL_X16 FILLER_187_1776 ();
 FILLCELL_X4 FILLER_187_1792 ();
 FILLCELL_X1 FILLER_187_1796 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X32 FILLER_188_1240 ();
 FILLCELL_X32 FILLER_188_1272 ();
 FILLCELL_X32 FILLER_188_1304 ();
 FILLCELL_X32 FILLER_188_1336 ();
 FILLCELL_X32 FILLER_188_1368 ();
 FILLCELL_X32 FILLER_188_1400 ();
 FILLCELL_X32 FILLER_188_1432 ();
 FILLCELL_X32 FILLER_188_1464 ();
 FILLCELL_X32 FILLER_188_1496 ();
 FILLCELL_X32 FILLER_188_1528 ();
 FILLCELL_X32 FILLER_188_1560 ();
 FILLCELL_X32 FILLER_188_1592 ();
 FILLCELL_X32 FILLER_188_1624 ();
 FILLCELL_X32 FILLER_188_1656 ();
 FILLCELL_X32 FILLER_188_1688 ();
 FILLCELL_X32 FILLER_188_1720 ();
 FILLCELL_X32 FILLER_188_1752 ();
 FILLCELL_X8 FILLER_188_1784 ();
 FILLCELL_X4 FILLER_188_1792 ();
 FILLCELL_X1 FILLER_188_1796 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X8 FILLER_189_1249 ();
 FILLCELL_X4 FILLER_189_1257 ();
 FILLCELL_X2 FILLER_189_1261 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X32 FILLER_189_1584 ();
 FILLCELL_X32 FILLER_189_1616 ();
 FILLCELL_X32 FILLER_189_1648 ();
 FILLCELL_X32 FILLER_189_1680 ();
 FILLCELL_X32 FILLER_189_1712 ();
 FILLCELL_X32 FILLER_189_1744 ();
 FILLCELL_X16 FILLER_189_1776 ();
 FILLCELL_X4 FILLER_189_1792 ();
 FILLCELL_X1 FILLER_189_1796 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X32 FILLER_190_1240 ();
 FILLCELL_X32 FILLER_190_1272 ();
 FILLCELL_X32 FILLER_190_1304 ();
 FILLCELL_X32 FILLER_190_1336 ();
 FILLCELL_X32 FILLER_190_1368 ();
 FILLCELL_X32 FILLER_190_1400 ();
 FILLCELL_X32 FILLER_190_1432 ();
 FILLCELL_X32 FILLER_190_1464 ();
 FILLCELL_X32 FILLER_190_1496 ();
 FILLCELL_X32 FILLER_190_1528 ();
 FILLCELL_X32 FILLER_190_1560 ();
 FILLCELL_X32 FILLER_190_1592 ();
 FILLCELL_X32 FILLER_190_1624 ();
 FILLCELL_X32 FILLER_190_1656 ();
 FILLCELL_X32 FILLER_190_1688 ();
 FILLCELL_X32 FILLER_190_1720 ();
 FILLCELL_X32 FILLER_190_1752 ();
 FILLCELL_X8 FILLER_190_1784 ();
 FILLCELL_X4 FILLER_190_1792 ();
 FILLCELL_X1 FILLER_190_1796 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X32 FILLER_191_1217 ();
 FILLCELL_X8 FILLER_191_1249 ();
 FILLCELL_X4 FILLER_191_1257 ();
 FILLCELL_X2 FILLER_191_1261 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X32 FILLER_191_1584 ();
 FILLCELL_X32 FILLER_191_1616 ();
 FILLCELL_X32 FILLER_191_1648 ();
 FILLCELL_X32 FILLER_191_1680 ();
 FILLCELL_X32 FILLER_191_1712 ();
 FILLCELL_X32 FILLER_191_1744 ();
 FILLCELL_X16 FILLER_191_1776 ();
 FILLCELL_X4 FILLER_191_1792 ();
 FILLCELL_X1 FILLER_191_1796 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X32 FILLER_192_1208 ();
 FILLCELL_X32 FILLER_192_1240 ();
 FILLCELL_X32 FILLER_192_1272 ();
 FILLCELL_X32 FILLER_192_1304 ();
 FILLCELL_X32 FILLER_192_1336 ();
 FILLCELL_X32 FILLER_192_1368 ();
 FILLCELL_X32 FILLER_192_1400 ();
 FILLCELL_X32 FILLER_192_1432 ();
 FILLCELL_X32 FILLER_192_1464 ();
 FILLCELL_X32 FILLER_192_1496 ();
 FILLCELL_X32 FILLER_192_1528 ();
 FILLCELL_X32 FILLER_192_1560 ();
 FILLCELL_X32 FILLER_192_1592 ();
 FILLCELL_X32 FILLER_192_1624 ();
 FILLCELL_X32 FILLER_192_1656 ();
 FILLCELL_X32 FILLER_192_1688 ();
 FILLCELL_X32 FILLER_192_1720 ();
 FILLCELL_X32 FILLER_192_1752 ();
 FILLCELL_X8 FILLER_192_1784 ();
 FILLCELL_X4 FILLER_192_1792 ();
 FILLCELL_X1 FILLER_192_1796 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X32 FILLER_193_1584 ();
 FILLCELL_X32 FILLER_193_1616 ();
 FILLCELL_X32 FILLER_193_1648 ();
 FILLCELL_X32 FILLER_193_1680 ();
 FILLCELL_X32 FILLER_193_1712 ();
 FILLCELL_X32 FILLER_193_1744 ();
 FILLCELL_X16 FILLER_193_1776 ();
 FILLCELL_X4 FILLER_193_1792 ();
 FILLCELL_X1 FILLER_193_1796 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X32 FILLER_194_1208 ();
 FILLCELL_X32 FILLER_194_1240 ();
 FILLCELL_X32 FILLER_194_1272 ();
 FILLCELL_X32 FILLER_194_1304 ();
 FILLCELL_X32 FILLER_194_1336 ();
 FILLCELL_X32 FILLER_194_1368 ();
 FILLCELL_X32 FILLER_194_1400 ();
 FILLCELL_X32 FILLER_194_1432 ();
 FILLCELL_X32 FILLER_194_1464 ();
 FILLCELL_X32 FILLER_194_1496 ();
 FILLCELL_X32 FILLER_194_1528 ();
 FILLCELL_X32 FILLER_194_1560 ();
 FILLCELL_X32 FILLER_194_1592 ();
 FILLCELL_X32 FILLER_194_1624 ();
 FILLCELL_X32 FILLER_194_1656 ();
 FILLCELL_X32 FILLER_194_1688 ();
 FILLCELL_X32 FILLER_194_1720 ();
 FILLCELL_X32 FILLER_194_1752 ();
 FILLCELL_X8 FILLER_194_1784 ();
 FILLCELL_X4 FILLER_194_1792 ();
 FILLCELL_X1 FILLER_194_1796 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X32 FILLER_195_1217 ();
 FILLCELL_X8 FILLER_195_1249 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X32 FILLER_195_1584 ();
 FILLCELL_X32 FILLER_195_1616 ();
 FILLCELL_X32 FILLER_195_1648 ();
 FILLCELL_X32 FILLER_195_1680 ();
 FILLCELL_X32 FILLER_195_1712 ();
 FILLCELL_X32 FILLER_195_1744 ();
 FILLCELL_X16 FILLER_195_1776 ();
 FILLCELL_X4 FILLER_195_1792 ();
 FILLCELL_X1 FILLER_195_1796 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X32 FILLER_196_1272 ();
 FILLCELL_X32 FILLER_196_1304 ();
 FILLCELL_X32 FILLER_196_1336 ();
 FILLCELL_X32 FILLER_196_1368 ();
 FILLCELL_X32 FILLER_196_1400 ();
 FILLCELL_X32 FILLER_196_1432 ();
 FILLCELL_X32 FILLER_196_1464 ();
 FILLCELL_X32 FILLER_196_1496 ();
 FILLCELL_X32 FILLER_196_1528 ();
 FILLCELL_X32 FILLER_196_1560 ();
 FILLCELL_X32 FILLER_196_1592 ();
 FILLCELL_X32 FILLER_196_1624 ();
 FILLCELL_X32 FILLER_196_1656 ();
 FILLCELL_X32 FILLER_196_1688 ();
 FILLCELL_X32 FILLER_196_1720 ();
 FILLCELL_X32 FILLER_196_1752 ();
 FILLCELL_X8 FILLER_196_1784 ();
 FILLCELL_X4 FILLER_196_1792 ();
 FILLCELL_X1 FILLER_196_1796 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X32 FILLER_197_1584 ();
 FILLCELL_X32 FILLER_197_1616 ();
 FILLCELL_X32 FILLER_197_1648 ();
 FILLCELL_X32 FILLER_197_1680 ();
 FILLCELL_X32 FILLER_197_1712 ();
 FILLCELL_X32 FILLER_197_1744 ();
 FILLCELL_X16 FILLER_197_1776 ();
 FILLCELL_X4 FILLER_197_1792 ();
 FILLCELL_X1 FILLER_197_1796 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X32 FILLER_198_1208 ();
 FILLCELL_X32 FILLER_198_1240 ();
 FILLCELL_X32 FILLER_198_1272 ();
 FILLCELL_X32 FILLER_198_1304 ();
 FILLCELL_X32 FILLER_198_1336 ();
 FILLCELL_X32 FILLER_198_1368 ();
 FILLCELL_X32 FILLER_198_1400 ();
 FILLCELL_X32 FILLER_198_1432 ();
 FILLCELL_X32 FILLER_198_1464 ();
 FILLCELL_X32 FILLER_198_1496 ();
 FILLCELL_X32 FILLER_198_1528 ();
 FILLCELL_X32 FILLER_198_1560 ();
 FILLCELL_X32 FILLER_198_1592 ();
 FILLCELL_X32 FILLER_198_1624 ();
 FILLCELL_X32 FILLER_198_1656 ();
 FILLCELL_X32 FILLER_198_1688 ();
 FILLCELL_X32 FILLER_198_1720 ();
 FILLCELL_X32 FILLER_198_1752 ();
 FILLCELL_X8 FILLER_198_1784 ();
 FILLCELL_X4 FILLER_198_1792 ();
 FILLCELL_X1 FILLER_198_1796 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X32 FILLER_199_1584 ();
 FILLCELL_X32 FILLER_199_1616 ();
 FILLCELL_X32 FILLER_199_1648 ();
 FILLCELL_X32 FILLER_199_1680 ();
 FILLCELL_X32 FILLER_199_1712 ();
 FILLCELL_X32 FILLER_199_1744 ();
 FILLCELL_X16 FILLER_199_1776 ();
 FILLCELL_X4 FILLER_199_1792 ();
 FILLCELL_X1 FILLER_199_1796 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X32 FILLER_200_1304 ();
 FILLCELL_X32 FILLER_200_1336 ();
 FILLCELL_X32 FILLER_200_1368 ();
 FILLCELL_X32 FILLER_200_1400 ();
 FILLCELL_X32 FILLER_200_1432 ();
 FILLCELL_X32 FILLER_200_1464 ();
 FILLCELL_X32 FILLER_200_1496 ();
 FILLCELL_X32 FILLER_200_1528 ();
 FILLCELL_X32 FILLER_200_1560 ();
 FILLCELL_X32 FILLER_200_1592 ();
 FILLCELL_X32 FILLER_200_1624 ();
 FILLCELL_X32 FILLER_200_1656 ();
 FILLCELL_X32 FILLER_200_1688 ();
 FILLCELL_X32 FILLER_200_1720 ();
 FILLCELL_X32 FILLER_200_1752 ();
 FILLCELL_X8 FILLER_200_1784 ();
 FILLCELL_X4 FILLER_200_1792 ();
 FILLCELL_X1 FILLER_200_1796 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X32 FILLER_201_1648 ();
 FILLCELL_X32 FILLER_201_1680 ();
 FILLCELL_X32 FILLER_201_1712 ();
 FILLCELL_X32 FILLER_201_1744 ();
 FILLCELL_X16 FILLER_201_1776 ();
 FILLCELL_X4 FILLER_201_1792 ();
 FILLCELL_X1 FILLER_201_1796 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X32 FILLER_202_1592 ();
 FILLCELL_X32 FILLER_202_1624 ();
 FILLCELL_X32 FILLER_202_1656 ();
 FILLCELL_X32 FILLER_202_1688 ();
 FILLCELL_X32 FILLER_202_1720 ();
 FILLCELL_X32 FILLER_202_1752 ();
 FILLCELL_X8 FILLER_202_1784 ();
 FILLCELL_X4 FILLER_202_1792 ();
 FILLCELL_X1 FILLER_202_1796 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X32 FILLER_203_1648 ();
 FILLCELL_X32 FILLER_203_1680 ();
 FILLCELL_X32 FILLER_203_1712 ();
 FILLCELL_X32 FILLER_203_1744 ();
 FILLCELL_X16 FILLER_203_1776 ();
 FILLCELL_X4 FILLER_203_1792 ();
 FILLCELL_X1 FILLER_203_1796 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X32 FILLER_204_1592 ();
 FILLCELL_X32 FILLER_204_1624 ();
 FILLCELL_X32 FILLER_204_1656 ();
 FILLCELL_X32 FILLER_204_1688 ();
 FILLCELL_X32 FILLER_204_1720 ();
 FILLCELL_X32 FILLER_204_1752 ();
 FILLCELL_X8 FILLER_204_1784 ();
 FILLCELL_X4 FILLER_204_1792 ();
 FILLCELL_X1 FILLER_204_1796 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X32 FILLER_205_1648 ();
 FILLCELL_X32 FILLER_205_1680 ();
 FILLCELL_X32 FILLER_205_1712 ();
 FILLCELL_X32 FILLER_205_1744 ();
 FILLCELL_X16 FILLER_205_1776 ();
 FILLCELL_X4 FILLER_205_1792 ();
 FILLCELL_X1 FILLER_205_1796 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X32 FILLER_206_1592 ();
 FILLCELL_X32 FILLER_206_1624 ();
 FILLCELL_X32 FILLER_206_1656 ();
 FILLCELL_X32 FILLER_206_1688 ();
 FILLCELL_X32 FILLER_206_1720 ();
 FILLCELL_X32 FILLER_206_1752 ();
 FILLCELL_X8 FILLER_206_1784 ();
 FILLCELL_X4 FILLER_206_1792 ();
 FILLCELL_X1 FILLER_206_1796 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X32 FILLER_207_1648 ();
 FILLCELL_X32 FILLER_207_1680 ();
 FILLCELL_X32 FILLER_207_1712 ();
 FILLCELL_X32 FILLER_207_1744 ();
 FILLCELL_X16 FILLER_207_1776 ();
 FILLCELL_X4 FILLER_207_1792 ();
 FILLCELL_X1 FILLER_207_1796 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X32 FILLER_208_1592 ();
 FILLCELL_X32 FILLER_208_1624 ();
 FILLCELL_X32 FILLER_208_1656 ();
 FILLCELL_X32 FILLER_208_1688 ();
 FILLCELL_X32 FILLER_208_1720 ();
 FILLCELL_X32 FILLER_208_1752 ();
 FILLCELL_X8 FILLER_208_1784 ();
 FILLCELL_X4 FILLER_208_1792 ();
 FILLCELL_X1 FILLER_208_1796 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X32 FILLER_209_1744 ();
 FILLCELL_X16 FILLER_209_1776 ();
 FILLCELL_X4 FILLER_209_1792 ();
 FILLCELL_X1 FILLER_209_1796 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X32 FILLER_210_1752 ();
 FILLCELL_X8 FILLER_210_1784 ();
 FILLCELL_X4 FILLER_210_1792 ();
 FILLCELL_X1 FILLER_210_1796 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X32 FILLER_211_1744 ();
 FILLCELL_X16 FILLER_211_1776 ();
 FILLCELL_X4 FILLER_211_1792 ();
 FILLCELL_X1 FILLER_211_1796 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X32 FILLER_212_1752 ();
 FILLCELL_X8 FILLER_212_1784 ();
 FILLCELL_X4 FILLER_212_1792 ();
 FILLCELL_X1 FILLER_212_1796 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X32 FILLER_213_1744 ();
 FILLCELL_X16 FILLER_213_1776 ();
 FILLCELL_X4 FILLER_213_1792 ();
 FILLCELL_X1 FILLER_213_1796 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X32 FILLER_214_1752 ();
 FILLCELL_X8 FILLER_214_1784 ();
 FILLCELL_X4 FILLER_214_1792 ();
 FILLCELL_X1 FILLER_214_1796 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X32 FILLER_215_1744 ();
 FILLCELL_X16 FILLER_215_1776 ();
 FILLCELL_X4 FILLER_215_1792 ();
 FILLCELL_X1 FILLER_215_1796 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X32 FILLER_216_1752 ();
 FILLCELL_X8 FILLER_216_1784 ();
 FILLCELL_X4 FILLER_216_1792 ();
 FILLCELL_X1 FILLER_216_1796 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X32 FILLER_217_1744 ();
 FILLCELL_X16 FILLER_217_1776 ();
 FILLCELL_X4 FILLER_217_1792 ();
 FILLCELL_X1 FILLER_217_1796 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X32 FILLER_218_1752 ();
 FILLCELL_X8 FILLER_218_1784 ();
 FILLCELL_X4 FILLER_218_1792 ();
 FILLCELL_X1 FILLER_218_1796 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X32 FILLER_219_1744 ();
 FILLCELL_X16 FILLER_219_1776 ();
 FILLCELL_X4 FILLER_219_1792 ();
 FILLCELL_X1 FILLER_219_1796 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X32 FILLER_220_1752 ();
 FILLCELL_X8 FILLER_220_1784 ();
 FILLCELL_X4 FILLER_220_1792 ();
 FILLCELL_X1 FILLER_220_1796 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X32 FILLER_221_1744 ();
 FILLCELL_X16 FILLER_221_1776 ();
 FILLCELL_X4 FILLER_221_1792 ();
 FILLCELL_X1 FILLER_221_1796 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X32 FILLER_222_1720 ();
 FILLCELL_X32 FILLER_222_1752 ();
 FILLCELL_X8 FILLER_222_1784 ();
 FILLCELL_X4 FILLER_222_1792 ();
 FILLCELL_X1 FILLER_222_1796 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X32 FILLER_223_1744 ();
 FILLCELL_X16 FILLER_223_1776 ();
 FILLCELL_X4 FILLER_223_1792 ();
 FILLCELL_X1 FILLER_223_1796 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X32 FILLER_224_1752 ();
 FILLCELL_X8 FILLER_224_1784 ();
 FILLCELL_X4 FILLER_224_1792 ();
 FILLCELL_X1 FILLER_224_1796 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X32 FILLER_225_1744 ();
 FILLCELL_X16 FILLER_225_1776 ();
 FILLCELL_X4 FILLER_225_1792 ();
 FILLCELL_X1 FILLER_225_1796 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X32 FILLER_226_1752 ();
 FILLCELL_X8 FILLER_226_1784 ();
 FILLCELL_X4 FILLER_226_1792 ();
 FILLCELL_X1 FILLER_226_1796 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X32 FILLER_227_1744 ();
 FILLCELL_X16 FILLER_227_1776 ();
 FILLCELL_X4 FILLER_227_1792 ();
 FILLCELL_X1 FILLER_227_1796 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X32 FILLER_228_1752 ();
 FILLCELL_X8 FILLER_228_1784 ();
 FILLCELL_X4 FILLER_228_1792 ();
 FILLCELL_X1 FILLER_228_1796 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X32 FILLER_229_1744 ();
 FILLCELL_X16 FILLER_229_1776 ();
 FILLCELL_X4 FILLER_229_1792 ();
 FILLCELL_X1 FILLER_229_1796 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X32 FILLER_230_1752 ();
 FILLCELL_X8 FILLER_230_1784 ();
 FILLCELL_X4 FILLER_230_1792 ();
 FILLCELL_X1 FILLER_230_1796 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X32 FILLER_231_1744 ();
 FILLCELL_X16 FILLER_231_1776 ();
 FILLCELL_X4 FILLER_231_1792 ();
 FILLCELL_X1 FILLER_231_1796 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X8 FILLER_232_888 ();
 FILLCELL_X4 FILLER_232_896 ();
 FILLCELL_X2 FILLER_232_900 ();
 FILLCELL_X1 FILLER_232_902 ();
 FILLCELL_X32 FILLER_232_905 ();
 FILLCELL_X8 FILLER_232_937 ();
 FILLCELL_X4 FILLER_232_945 ();
 FILLCELL_X2 FILLER_232_949 ();
 FILLCELL_X32 FILLER_232_956 ();
 FILLCELL_X32 FILLER_232_988 ();
 FILLCELL_X32 FILLER_232_1020 ();
 FILLCELL_X32 FILLER_232_1052 ();
 FILLCELL_X32 FILLER_232_1084 ();
 FILLCELL_X32 FILLER_232_1116 ();
 FILLCELL_X32 FILLER_232_1148 ();
 FILLCELL_X32 FILLER_232_1180 ();
 FILLCELL_X32 FILLER_232_1212 ();
 FILLCELL_X32 FILLER_232_1244 ();
 FILLCELL_X32 FILLER_232_1276 ();
 FILLCELL_X32 FILLER_232_1308 ();
 FILLCELL_X32 FILLER_232_1340 ();
 FILLCELL_X32 FILLER_232_1372 ();
 FILLCELL_X32 FILLER_232_1404 ();
 FILLCELL_X32 FILLER_232_1436 ();
 FILLCELL_X32 FILLER_232_1468 ();
 FILLCELL_X32 FILLER_232_1500 ();
 FILLCELL_X32 FILLER_232_1532 ();
 FILLCELL_X32 FILLER_232_1564 ();
 FILLCELL_X32 FILLER_232_1596 ();
 FILLCELL_X32 FILLER_232_1628 ();
 FILLCELL_X32 FILLER_232_1660 ();
 FILLCELL_X32 FILLER_232_1692 ();
 FILLCELL_X32 FILLER_232_1724 ();
 FILLCELL_X32 FILLER_232_1756 ();
 FILLCELL_X8 FILLER_232_1788 ();
 FILLCELL_X1 FILLER_232_1796 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X16 FILLER_233_865 ();
 FILLCELL_X8 FILLER_233_881 ();
 FILLCELL_X4 FILLER_233_889 ();
 FILLCELL_X2 FILLER_233_893 ();
 FILLCELL_X1 FILLER_233_895 ();
 FILLCELL_X16 FILLER_233_925 ();
 FILLCELL_X4 FILLER_233_941 ();
 FILLCELL_X2 FILLER_233_945 ();
 FILLCELL_X1 FILLER_233_947 ();
 FILLCELL_X32 FILLER_233_958 ();
 FILLCELL_X32 FILLER_233_990 ();
 FILLCELL_X32 FILLER_233_1022 ();
 FILLCELL_X32 FILLER_233_1054 ();
 FILLCELL_X32 FILLER_233_1086 ();
 FILLCELL_X32 FILLER_233_1118 ();
 FILLCELL_X32 FILLER_233_1150 ();
 FILLCELL_X32 FILLER_233_1182 ();
 FILLCELL_X32 FILLER_233_1214 ();
 FILLCELL_X16 FILLER_233_1246 ();
 FILLCELL_X1 FILLER_233_1262 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X32 FILLER_233_1744 ();
 FILLCELL_X16 FILLER_233_1776 ();
 FILLCELL_X4 FILLER_233_1792 ();
 FILLCELL_X1 FILLER_233_1796 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X16 FILLER_234_888 ();
 FILLCELL_X8 FILLER_234_904 ();
 FILLCELL_X2 FILLER_234_912 ();
 FILLCELL_X1 FILLER_234_914 ();
 FILLCELL_X16 FILLER_234_921 ();
 FILLCELL_X2 FILLER_234_937 ();
 FILLCELL_X1 FILLER_234_939 ();
 FILLCELL_X32 FILLER_234_953 ();
 FILLCELL_X32 FILLER_234_985 ();
 FILLCELL_X32 FILLER_234_1017 ();
 FILLCELL_X32 FILLER_234_1049 ();
 FILLCELL_X32 FILLER_234_1081 ();
 FILLCELL_X32 FILLER_234_1113 ();
 FILLCELL_X32 FILLER_234_1145 ();
 FILLCELL_X32 FILLER_234_1177 ();
 FILLCELL_X32 FILLER_234_1209 ();
 FILLCELL_X32 FILLER_234_1241 ();
 FILLCELL_X32 FILLER_234_1273 ();
 FILLCELL_X32 FILLER_234_1305 ();
 FILLCELL_X32 FILLER_234_1337 ();
 FILLCELL_X32 FILLER_234_1369 ();
 FILLCELL_X32 FILLER_234_1401 ();
 FILLCELL_X32 FILLER_234_1433 ();
 FILLCELL_X32 FILLER_234_1465 ();
 FILLCELL_X32 FILLER_234_1497 ();
 FILLCELL_X32 FILLER_234_1529 ();
 FILLCELL_X32 FILLER_234_1561 ();
 FILLCELL_X32 FILLER_234_1593 ();
 FILLCELL_X32 FILLER_234_1625 ();
 FILLCELL_X32 FILLER_234_1657 ();
 FILLCELL_X32 FILLER_234_1689 ();
 FILLCELL_X32 FILLER_234_1721 ();
 FILLCELL_X32 FILLER_234_1753 ();
 FILLCELL_X8 FILLER_234_1785 ();
 FILLCELL_X4 FILLER_234_1793 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X8 FILLER_235_897 ();
 FILLCELL_X1 FILLER_235_905 ();
 FILLCELL_X32 FILLER_235_916 ();
 FILLCELL_X32 FILLER_235_948 ();
 FILLCELL_X32 FILLER_235_980 ();
 FILLCELL_X32 FILLER_235_1012 ();
 FILLCELL_X32 FILLER_235_1044 ();
 FILLCELL_X32 FILLER_235_1076 ();
 FILLCELL_X32 FILLER_235_1108 ();
 FILLCELL_X32 FILLER_235_1140 ();
 FILLCELL_X32 FILLER_235_1172 ();
 FILLCELL_X32 FILLER_235_1204 ();
 FILLCELL_X16 FILLER_235_1236 ();
 FILLCELL_X8 FILLER_235_1252 ();
 FILLCELL_X2 FILLER_235_1260 ();
 FILLCELL_X1 FILLER_235_1262 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X32 FILLER_235_1744 ();
 FILLCELL_X16 FILLER_235_1776 ();
 FILLCELL_X4 FILLER_235_1792 ();
 FILLCELL_X1 FILLER_235_1796 ();
 FILLCELL_X32 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_33 ();
 FILLCELL_X32 FILLER_236_65 ();
 FILLCELL_X32 FILLER_236_97 ();
 FILLCELL_X32 FILLER_236_129 ();
 FILLCELL_X32 FILLER_236_161 ();
 FILLCELL_X32 FILLER_236_193 ();
 FILLCELL_X32 FILLER_236_225 ();
 FILLCELL_X32 FILLER_236_257 ();
 FILLCELL_X32 FILLER_236_289 ();
 FILLCELL_X32 FILLER_236_321 ();
 FILLCELL_X32 FILLER_236_353 ();
 FILLCELL_X32 FILLER_236_385 ();
 FILLCELL_X32 FILLER_236_417 ();
 FILLCELL_X32 FILLER_236_449 ();
 FILLCELL_X32 FILLER_236_481 ();
 FILLCELL_X32 FILLER_236_513 ();
 FILLCELL_X32 FILLER_236_545 ();
 FILLCELL_X32 FILLER_236_577 ();
 FILLCELL_X16 FILLER_236_609 ();
 FILLCELL_X4 FILLER_236_625 ();
 FILLCELL_X2 FILLER_236_629 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X16 FILLER_236_888 ();
 FILLCELL_X2 FILLER_236_904 ();
 FILLCELL_X1 FILLER_236_906 ();
 FILLCELL_X16 FILLER_236_924 ();
 FILLCELL_X8 FILLER_236_940 ();
 FILLCELL_X32 FILLER_236_961 ();
 FILLCELL_X32 FILLER_236_993 ();
 FILLCELL_X32 FILLER_236_1025 ();
 FILLCELL_X32 FILLER_236_1057 ();
 FILLCELL_X32 FILLER_236_1089 ();
 FILLCELL_X32 FILLER_236_1121 ();
 FILLCELL_X32 FILLER_236_1153 ();
 FILLCELL_X32 FILLER_236_1185 ();
 FILLCELL_X32 FILLER_236_1217 ();
 FILLCELL_X32 FILLER_236_1249 ();
 FILLCELL_X32 FILLER_236_1281 ();
 FILLCELL_X32 FILLER_236_1313 ();
 FILLCELL_X32 FILLER_236_1345 ();
 FILLCELL_X32 FILLER_236_1377 ();
 FILLCELL_X32 FILLER_236_1409 ();
 FILLCELL_X32 FILLER_236_1441 ();
 FILLCELL_X32 FILLER_236_1473 ();
 FILLCELL_X32 FILLER_236_1505 ();
 FILLCELL_X32 FILLER_236_1537 ();
 FILLCELL_X32 FILLER_236_1569 ();
 FILLCELL_X32 FILLER_236_1601 ();
 FILLCELL_X32 FILLER_236_1633 ();
 FILLCELL_X32 FILLER_236_1665 ();
 FILLCELL_X32 FILLER_236_1697 ();
 FILLCELL_X32 FILLER_236_1729 ();
 FILLCELL_X32 FILLER_236_1761 ();
 FILLCELL_X4 FILLER_236_1793 ();
 FILLCELL_X32 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_33 ();
 FILLCELL_X32 FILLER_237_65 ();
 FILLCELL_X32 FILLER_237_97 ();
 FILLCELL_X32 FILLER_237_129 ();
 FILLCELL_X32 FILLER_237_161 ();
 FILLCELL_X32 FILLER_237_193 ();
 FILLCELL_X32 FILLER_237_225 ();
 FILLCELL_X32 FILLER_237_257 ();
 FILLCELL_X32 FILLER_237_289 ();
 FILLCELL_X32 FILLER_237_321 ();
 FILLCELL_X32 FILLER_237_353 ();
 FILLCELL_X32 FILLER_237_385 ();
 FILLCELL_X32 FILLER_237_417 ();
 FILLCELL_X32 FILLER_237_449 ();
 FILLCELL_X32 FILLER_237_481 ();
 FILLCELL_X32 FILLER_237_513 ();
 FILLCELL_X32 FILLER_237_545 ();
 FILLCELL_X32 FILLER_237_577 ();
 FILLCELL_X32 FILLER_237_609 ();
 FILLCELL_X32 FILLER_237_641 ();
 FILLCELL_X32 FILLER_237_673 ();
 FILLCELL_X32 FILLER_237_705 ();
 FILLCELL_X32 FILLER_237_737 ();
 FILLCELL_X32 FILLER_237_769 ();
 FILLCELL_X32 FILLER_237_801 ();
 FILLCELL_X32 FILLER_237_833 ();
 FILLCELL_X2 FILLER_237_865 ();
 FILLCELL_X1 FILLER_237_867 ();
 FILLCELL_X16 FILLER_237_878 ();
 FILLCELL_X4 FILLER_237_894 ();
 FILLCELL_X2 FILLER_237_898 ();
 FILLCELL_X16 FILLER_237_919 ();
 FILLCELL_X1 FILLER_237_935 ();
 FILLCELL_X32 FILLER_237_961 ();
 FILLCELL_X32 FILLER_237_993 ();
 FILLCELL_X32 FILLER_237_1025 ();
 FILLCELL_X32 FILLER_237_1057 ();
 FILLCELL_X32 FILLER_237_1089 ();
 FILLCELL_X32 FILLER_237_1121 ();
 FILLCELL_X32 FILLER_237_1153 ();
 FILLCELL_X32 FILLER_237_1185 ();
 FILLCELL_X32 FILLER_237_1217 ();
 FILLCELL_X8 FILLER_237_1249 ();
 FILLCELL_X4 FILLER_237_1257 ();
 FILLCELL_X2 FILLER_237_1261 ();
 FILLCELL_X32 FILLER_237_1264 ();
 FILLCELL_X32 FILLER_237_1296 ();
 FILLCELL_X32 FILLER_237_1328 ();
 FILLCELL_X32 FILLER_237_1360 ();
 FILLCELL_X32 FILLER_237_1392 ();
 FILLCELL_X32 FILLER_237_1424 ();
 FILLCELL_X32 FILLER_237_1456 ();
 FILLCELL_X32 FILLER_237_1488 ();
 FILLCELL_X32 FILLER_237_1520 ();
 FILLCELL_X32 FILLER_237_1552 ();
 FILLCELL_X32 FILLER_237_1584 ();
 FILLCELL_X32 FILLER_237_1616 ();
 FILLCELL_X32 FILLER_237_1648 ();
 FILLCELL_X32 FILLER_237_1680 ();
 FILLCELL_X32 FILLER_237_1712 ();
 FILLCELL_X32 FILLER_237_1744 ();
 FILLCELL_X16 FILLER_237_1776 ();
 FILLCELL_X4 FILLER_237_1792 ();
 FILLCELL_X1 FILLER_237_1796 ();
 FILLCELL_X32 FILLER_238_1 ();
 FILLCELL_X32 FILLER_238_33 ();
 FILLCELL_X32 FILLER_238_65 ();
 FILLCELL_X32 FILLER_238_97 ();
 FILLCELL_X32 FILLER_238_129 ();
 FILLCELL_X32 FILLER_238_161 ();
 FILLCELL_X32 FILLER_238_193 ();
 FILLCELL_X32 FILLER_238_225 ();
 FILLCELL_X32 FILLER_238_257 ();
 FILLCELL_X32 FILLER_238_289 ();
 FILLCELL_X32 FILLER_238_321 ();
 FILLCELL_X32 FILLER_238_353 ();
 FILLCELL_X32 FILLER_238_385 ();
 FILLCELL_X32 FILLER_238_417 ();
 FILLCELL_X32 FILLER_238_449 ();
 FILLCELL_X32 FILLER_238_481 ();
 FILLCELL_X32 FILLER_238_513 ();
 FILLCELL_X32 FILLER_238_545 ();
 FILLCELL_X32 FILLER_238_577 ();
 FILLCELL_X16 FILLER_238_609 ();
 FILLCELL_X4 FILLER_238_625 ();
 FILLCELL_X2 FILLER_238_629 ();
 FILLCELL_X32 FILLER_238_632 ();
 FILLCELL_X32 FILLER_238_664 ();
 FILLCELL_X32 FILLER_238_696 ();
 FILLCELL_X32 FILLER_238_728 ();
 FILLCELL_X32 FILLER_238_760 ();
 FILLCELL_X32 FILLER_238_792 ();
 FILLCELL_X32 FILLER_238_824 ();
 FILLCELL_X8 FILLER_238_856 ();
 FILLCELL_X2 FILLER_238_864 ();
 FILLCELL_X1 FILLER_238_866 ();
 FILLCELL_X1 FILLER_238_871 ();
 FILLCELL_X32 FILLER_238_878 ();
 FILLCELL_X4 FILLER_238_910 ();
 FILLCELL_X2 FILLER_238_914 ();
 FILLCELL_X4 FILLER_238_932 ();
 FILLCELL_X1 FILLER_238_938 ();
 FILLCELL_X4 FILLER_238_946 ();
 FILLCELL_X32 FILLER_238_978 ();
 FILLCELL_X32 FILLER_238_1010 ();
 FILLCELL_X32 FILLER_238_1042 ();
 FILLCELL_X32 FILLER_238_1074 ();
 FILLCELL_X32 FILLER_238_1106 ();
 FILLCELL_X32 FILLER_238_1138 ();
 FILLCELL_X32 FILLER_238_1170 ();
 FILLCELL_X32 FILLER_238_1202 ();
 FILLCELL_X32 FILLER_238_1234 ();
 FILLCELL_X32 FILLER_238_1266 ();
 FILLCELL_X32 FILLER_238_1298 ();
 FILLCELL_X32 FILLER_238_1330 ();
 FILLCELL_X32 FILLER_238_1362 ();
 FILLCELL_X32 FILLER_238_1394 ();
 FILLCELL_X32 FILLER_238_1426 ();
 FILLCELL_X32 FILLER_238_1458 ();
 FILLCELL_X32 FILLER_238_1490 ();
 FILLCELL_X32 FILLER_238_1522 ();
 FILLCELL_X32 FILLER_238_1554 ();
 FILLCELL_X32 FILLER_238_1586 ();
 FILLCELL_X32 FILLER_238_1618 ();
 FILLCELL_X32 FILLER_238_1650 ();
 FILLCELL_X32 FILLER_238_1682 ();
 FILLCELL_X32 FILLER_238_1714 ();
 FILLCELL_X32 FILLER_238_1746 ();
 FILLCELL_X16 FILLER_238_1778 ();
 FILLCELL_X2 FILLER_238_1794 ();
 FILLCELL_X1 FILLER_238_1796 ();
 FILLCELL_X32 FILLER_239_1 ();
 FILLCELL_X32 FILLER_239_33 ();
 FILLCELL_X32 FILLER_239_65 ();
 FILLCELL_X32 FILLER_239_97 ();
 FILLCELL_X32 FILLER_239_129 ();
 FILLCELL_X32 FILLER_239_161 ();
 FILLCELL_X32 FILLER_239_193 ();
 FILLCELL_X32 FILLER_239_225 ();
 FILLCELL_X32 FILLER_239_257 ();
 FILLCELL_X32 FILLER_239_289 ();
 FILLCELL_X32 FILLER_239_321 ();
 FILLCELL_X32 FILLER_239_353 ();
 FILLCELL_X32 FILLER_239_385 ();
 FILLCELL_X32 FILLER_239_417 ();
 FILLCELL_X32 FILLER_239_449 ();
 FILLCELL_X32 FILLER_239_481 ();
 FILLCELL_X32 FILLER_239_513 ();
 FILLCELL_X32 FILLER_239_545 ();
 FILLCELL_X32 FILLER_239_577 ();
 FILLCELL_X32 FILLER_239_609 ();
 FILLCELL_X32 FILLER_239_641 ();
 FILLCELL_X32 FILLER_239_673 ();
 FILLCELL_X32 FILLER_239_705 ();
 FILLCELL_X32 FILLER_239_737 ();
 FILLCELL_X32 FILLER_239_769 ();
 FILLCELL_X32 FILLER_239_801 ();
 FILLCELL_X16 FILLER_239_833 ();
 FILLCELL_X8 FILLER_239_849 ();
 FILLCELL_X2 FILLER_239_857 ();
 FILLCELL_X32 FILLER_239_876 ();
 FILLCELL_X16 FILLER_239_908 ();
 FILLCELL_X1 FILLER_239_924 ();
 FILLCELL_X16 FILLER_239_927 ();
 FILLCELL_X4 FILLER_239_943 ();
 FILLCELL_X4 FILLER_239_953 ();
 FILLCELL_X2 FILLER_239_957 ();
 FILLCELL_X1 FILLER_239_959 ();
 FILLCELL_X32 FILLER_239_977 ();
 FILLCELL_X32 FILLER_239_1009 ();
 FILLCELL_X32 FILLER_239_1041 ();
 FILLCELL_X32 FILLER_239_1073 ();
 FILLCELL_X32 FILLER_239_1105 ();
 FILLCELL_X32 FILLER_239_1137 ();
 FILLCELL_X32 FILLER_239_1169 ();
 FILLCELL_X32 FILLER_239_1201 ();
 FILLCELL_X16 FILLER_239_1233 ();
 FILLCELL_X8 FILLER_239_1249 ();
 FILLCELL_X4 FILLER_239_1257 ();
 FILLCELL_X2 FILLER_239_1261 ();
 FILLCELL_X32 FILLER_239_1264 ();
 FILLCELL_X32 FILLER_239_1296 ();
 FILLCELL_X32 FILLER_239_1328 ();
 FILLCELL_X32 FILLER_239_1360 ();
 FILLCELL_X32 FILLER_239_1392 ();
 FILLCELL_X32 FILLER_239_1424 ();
 FILLCELL_X32 FILLER_239_1456 ();
 FILLCELL_X32 FILLER_239_1488 ();
 FILLCELL_X32 FILLER_239_1520 ();
 FILLCELL_X32 FILLER_239_1552 ();
 FILLCELL_X32 FILLER_239_1584 ();
 FILLCELL_X32 FILLER_239_1616 ();
 FILLCELL_X32 FILLER_239_1648 ();
 FILLCELL_X32 FILLER_239_1680 ();
 FILLCELL_X32 FILLER_239_1712 ();
 FILLCELL_X32 FILLER_239_1744 ();
 FILLCELL_X16 FILLER_239_1776 ();
 FILLCELL_X4 FILLER_239_1792 ();
 FILLCELL_X1 FILLER_239_1796 ();
 FILLCELL_X32 FILLER_240_1 ();
 FILLCELL_X32 FILLER_240_33 ();
 FILLCELL_X32 FILLER_240_65 ();
 FILLCELL_X32 FILLER_240_97 ();
 FILLCELL_X32 FILLER_240_129 ();
 FILLCELL_X32 FILLER_240_161 ();
 FILLCELL_X32 FILLER_240_193 ();
 FILLCELL_X32 FILLER_240_225 ();
 FILLCELL_X32 FILLER_240_257 ();
 FILLCELL_X32 FILLER_240_289 ();
 FILLCELL_X32 FILLER_240_321 ();
 FILLCELL_X32 FILLER_240_353 ();
 FILLCELL_X32 FILLER_240_385 ();
 FILLCELL_X32 FILLER_240_417 ();
 FILLCELL_X32 FILLER_240_449 ();
 FILLCELL_X32 FILLER_240_481 ();
 FILLCELL_X32 FILLER_240_513 ();
 FILLCELL_X32 FILLER_240_545 ();
 FILLCELL_X32 FILLER_240_577 ();
 FILLCELL_X16 FILLER_240_609 ();
 FILLCELL_X4 FILLER_240_625 ();
 FILLCELL_X2 FILLER_240_629 ();
 FILLCELL_X32 FILLER_240_632 ();
 FILLCELL_X32 FILLER_240_664 ();
 FILLCELL_X32 FILLER_240_696 ();
 FILLCELL_X32 FILLER_240_728 ();
 FILLCELL_X32 FILLER_240_760 ();
 FILLCELL_X32 FILLER_240_792 ();
 FILLCELL_X8 FILLER_240_824 ();
 FILLCELL_X2 FILLER_240_832 ();
 FILLCELL_X1 FILLER_240_834 ();
 FILLCELL_X32 FILLER_240_855 ();
 FILLCELL_X16 FILLER_240_887 ();
 FILLCELL_X8 FILLER_240_909 ();
 FILLCELL_X1 FILLER_240_917 ();
 FILLCELL_X4 FILLER_240_925 ();
 FILLCELL_X2 FILLER_240_929 ();
 FILLCELL_X8 FILLER_240_941 ();
 FILLCELL_X2 FILLER_240_949 ();
 FILLCELL_X32 FILLER_240_966 ();
 FILLCELL_X32 FILLER_240_998 ();
 FILLCELL_X32 FILLER_240_1030 ();
 FILLCELL_X32 FILLER_240_1062 ();
 FILLCELL_X32 FILLER_240_1094 ();
 FILLCELL_X32 FILLER_240_1126 ();
 FILLCELL_X32 FILLER_240_1158 ();
 FILLCELL_X32 FILLER_240_1190 ();
 FILLCELL_X32 FILLER_240_1222 ();
 FILLCELL_X32 FILLER_240_1254 ();
 FILLCELL_X32 FILLER_240_1286 ();
 FILLCELL_X32 FILLER_240_1318 ();
 FILLCELL_X32 FILLER_240_1350 ();
 FILLCELL_X32 FILLER_240_1382 ();
 FILLCELL_X32 FILLER_240_1414 ();
 FILLCELL_X32 FILLER_240_1446 ();
 FILLCELL_X32 FILLER_240_1478 ();
 FILLCELL_X32 FILLER_240_1510 ();
 FILLCELL_X32 FILLER_240_1542 ();
 FILLCELL_X32 FILLER_240_1574 ();
 FILLCELL_X32 FILLER_240_1606 ();
 FILLCELL_X32 FILLER_240_1638 ();
 FILLCELL_X32 FILLER_240_1670 ();
 FILLCELL_X32 FILLER_240_1702 ();
 FILLCELL_X32 FILLER_240_1734 ();
 FILLCELL_X16 FILLER_240_1766 ();
 FILLCELL_X8 FILLER_240_1782 ();
 FILLCELL_X4 FILLER_240_1790 ();
 FILLCELL_X2 FILLER_240_1794 ();
 FILLCELL_X1 FILLER_240_1796 ();
 FILLCELL_X32 FILLER_241_1 ();
 FILLCELL_X32 FILLER_241_33 ();
 FILLCELL_X32 FILLER_241_65 ();
 FILLCELL_X32 FILLER_241_97 ();
 FILLCELL_X32 FILLER_241_129 ();
 FILLCELL_X32 FILLER_241_161 ();
 FILLCELL_X32 FILLER_241_193 ();
 FILLCELL_X32 FILLER_241_225 ();
 FILLCELL_X32 FILLER_241_257 ();
 FILLCELL_X32 FILLER_241_289 ();
 FILLCELL_X32 FILLER_241_321 ();
 FILLCELL_X32 FILLER_241_353 ();
 FILLCELL_X32 FILLER_241_385 ();
 FILLCELL_X32 FILLER_241_417 ();
 FILLCELL_X32 FILLER_241_449 ();
 FILLCELL_X32 FILLER_241_481 ();
 FILLCELL_X32 FILLER_241_513 ();
 FILLCELL_X32 FILLER_241_545 ();
 FILLCELL_X32 FILLER_241_577 ();
 FILLCELL_X32 FILLER_241_609 ();
 FILLCELL_X32 FILLER_241_641 ();
 FILLCELL_X32 FILLER_241_673 ();
 FILLCELL_X32 FILLER_241_705 ();
 FILLCELL_X32 FILLER_241_737 ();
 FILLCELL_X32 FILLER_241_769 ();
 FILLCELL_X32 FILLER_241_801 ();
 FILLCELL_X4 FILLER_241_833 ();
 FILLCELL_X8 FILLER_241_847 ();
 FILLCELL_X4 FILLER_241_855 ();
 FILLCELL_X2 FILLER_241_859 ();
 FILLCELL_X1 FILLER_241_861 ();
 FILLCELL_X2 FILLER_241_878 ();
 FILLCELL_X1 FILLER_241_880 ();
 FILLCELL_X2 FILLER_241_900 ();
 FILLCELL_X4 FILLER_241_918 ();
 FILLCELL_X2 FILLER_241_932 ();
 FILLCELL_X8 FILLER_241_937 ();
 FILLCELL_X2 FILLER_241_945 ();
 FILLCELL_X1 FILLER_241_947 ();
 FILLCELL_X4 FILLER_241_951 ();
 FILLCELL_X32 FILLER_241_961 ();
 FILLCELL_X16 FILLER_241_993 ();
 FILLCELL_X4 FILLER_241_1009 ();
 FILLCELL_X1 FILLER_241_1013 ();
 FILLCELL_X32 FILLER_241_1021 ();
 FILLCELL_X32 FILLER_241_1053 ();
 FILLCELL_X32 FILLER_241_1085 ();
 FILLCELL_X32 FILLER_241_1117 ();
 FILLCELL_X32 FILLER_241_1149 ();
 FILLCELL_X32 FILLER_241_1181 ();
 FILLCELL_X32 FILLER_241_1213 ();
 FILLCELL_X16 FILLER_241_1245 ();
 FILLCELL_X2 FILLER_241_1261 ();
 FILLCELL_X32 FILLER_241_1264 ();
 FILLCELL_X32 FILLER_241_1296 ();
 FILLCELL_X32 FILLER_241_1328 ();
 FILLCELL_X32 FILLER_241_1360 ();
 FILLCELL_X32 FILLER_241_1392 ();
 FILLCELL_X32 FILLER_241_1424 ();
 FILLCELL_X32 FILLER_241_1456 ();
 FILLCELL_X32 FILLER_241_1488 ();
 FILLCELL_X32 FILLER_241_1520 ();
 FILLCELL_X32 FILLER_241_1552 ();
 FILLCELL_X32 FILLER_241_1584 ();
 FILLCELL_X32 FILLER_241_1616 ();
 FILLCELL_X32 FILLER_241_1648 ();
 FILLCELL_X32 FILLER_241_1680 ();
 FILLCELL_X32 FILLER_241_1712 ();
 FILLCELL_X32 FILLER_241_1744 ();
 FILLCELL_X16 FILLER_241_1776 ();
 FILLCELL_X4 FILLER_241_1792 ();
 FILLCELL_X1 FILLER_241_1796 ();
 FILLCELL_X32 FILLER_242_1 ();
 FILLCELL_X32 FILLER_242_33 ();
 FILLCELL_X32 FILLER_242_65 ();
 FILLCELL_X32 FILLER_242_97 ();
 FILLCELL_X32 FILLER_242_129 ();
 FILLCELL_X32 FILLER_242_161 ();
 FILLCELL_X32 FILLER_242_193 ();
 FILLCELL_X32 FILLER_242_225 ();
 FILLCELL_X32 FILLER_242_257 ();
 FILLCELL_X32 FILLER_242_289 ();
 FILLCELL_X32 FILLER_242_321 ();
 FILLCELL_X32 FILLER_242_353 ();
 FILLCELL_X32 FILLER_242_385 ();
 FILLCELL_X32 FILLER_242_417 ();
 FILLCELL_X32 FILLER_242_449 ();
 FILLCELL_X32 FILLER_242_481 ();
 FILLCELL_X32 FILLER_242_513 ();
 FILLCELL_X32 FILLER_242_545 ();
 FILLCELL_X32 FILLER_242_577 ();
 FILLCELL_X16 FILLER_242_609 ();
 FILLCELL_X4 FILLER_242_625 ();
 FILLCELL_X2 FILLER_242_629 ();
 FILLCELL_X32 FILLER_242_632 ();
 FILLCELL_X32 FILLER_242_664 ();
 FILLCELL_X32 FILLER_242_696 ();
 FILLCELL_X32 FILLER_242_728 ();
 FILLCELL_X32 FILLER_242_760 ();
 FILLCELL_X32 FILLER_242_792 ();
 FILLCELL_X8 FILLER_242_824 ();
 FILLCELL_X4 FILLER_242_832 ();
 FILLCELL_X1 FILLER_242_836 ();
 FILLCELL_X2 FILLER_242_843 ();
 FILLCELL_X1 FILLER_242_845 ();
 FILLCELL_X4 FILLER_242_855 ();
 FILLCELL_X1 FILLER_242_859 ();
 FILLCELL_X1 FILLER_242_863 ();
 FILLCELL_X2 FILLER_242_867 ();
 FILLCELL_X1 FILLER_242_887 ();
 FILLCELL_X1 FILLER_242_891 ();
 FILLCELL_X1 FILLER_242_895 ();
 FILLCELL_X4 FILLER_242_923 ();
 FILLCELL_X2 FILLER_242_927 ();
 FILLCELL_X4 FILLER_242_938 ();
 FILLCELL_X2 FILLER_242_942 ();
 FILLCELL_X1 FILLER_242_947 ();
 FILLCELL_X2 FILLER_242_954 ();
 FILLCELL_X2 FILLER_242_969 ();
 FILLCELL_X16 FILLER_242_975 ();
 FILLCELL_X8 FILLER_242_991 ();
 FILLCELL_X1 FILLER_242_999 ();
 FILLCELL_X16 FILLER_242_1003 ();
 FILLCELL_X4 FILLER_242_1019 ();
 FILLCELL_X1 FILLER_242_1030 ();
 FILLCELL_X32 FILLER_242_1034 ();
 FILLCELL_X32 FILLER_242_1066 ();
 FILLCELL_X32 FILLER_242_1098 ();
 FILLCELL_X32 FILLER_242_1130 ();
 FILLCELL_X32 FILLER_242_1162 ();
 FILLCELL_X32 FILLER_242_1194 ();
 FILLCELL_X32 FILLER_242_1226 ();
 FILLCELL_X4 FILLER_242_1258 ();
 FILLCELL_X32 FILLER_242_1263 ();
 FILLCELL_X32 FILLER_242_1295 ();
 FILLCELL_X32 FILLER_242_1327 ();
 FILLCELL_X32 FILLER_242_1359 ();
 FILLCELL_X32 FILLER_242_1391 ();
 FILLCELL_X32 FILLER_242_1423 ();
 FILLCELL_X32 FILLER_242_1455 ();
 FILLCELL_X32 FILLER_242_1487 ();
 FILLCELL_X32 FILLER_242_1519 ();
 FILLCELL_X32 FILLER_242_1551 ();
 FILLCELL_X32 FILLER_242_1583 ();
 FILLCELL_X32 FILLER_242_1615 ();
 FILLCELL_X32 FILLER_242_1647 ();
 FILLCELL_X32 FILLER_242_1679 ();
 FILLCELL_X32 FILLER_242_1711 ();
 FILLCELL_X32 FILLER_242_1743 ();
 FILLCELL_X16 FILLER_242_1775 ();
 FILLCELL_X4 FILLER_242_1791 ();
 FILLCELL_X2 FILLER_242_1795 ();
endmodule
