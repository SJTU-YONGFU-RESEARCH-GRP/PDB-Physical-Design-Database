module bist_controller (bist_done,
    bist_pass,
    bist_start,
    clk,
    mem_enable,
    mem_write,
    rst_n,
    error_addr,
    error_count,
    mem_addr,
    mem_rdata,
    mem_wdata);
 output bist_done;
 output bist_pass;
 input bist_start;
 input clk;
 output mem_enable;
 output mem_write;
 input rst_n;
 output [4:0] error_addr;
 output [31:0] error_count;
 output [4:0] mem_addr;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire phase_complete;
 wire read_phase;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net113;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _372_ (.I(net77),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _373_ (.I(net76),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _374_ (.I(_363_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _375_ (.A1(_051_),
    .A2(_052_),
    .A3(_053_),
    .Z(_366_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _376_ (.I(_366_),
    .ZN(_369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _377_ (.I(net78),
    .ZN(_365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _378_ (.I(net42),
    .ZN(_353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _379_ (.I(net74),
    .ZN(_359_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _380_ (.I(net53),
    .ZN(_354_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _381_ (.I(net75),
    .ZN(_360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _382_ (.I(\state[3] ),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _383_ (.I(\state[2] ),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _384_ (.I(\state[0] ),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _385_ (.A1(_056_),
    .A2(\state[1] ),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _386_ (.A1(_054_),
    .A2(_055_),
    .A3(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _387_ (.I(_361_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _388_ (.A1(net77),
    .A2(net76),
    .A3(_059_),
    .A4(net78),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _389_ (.A1(_058_),
    .A2(_060_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _390_ (.I(\state[1] ),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _391_ (.A1(_056_),
    .A2(_062_),
    .A3(_055_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _392_ (.I(\state[1] ),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _393_ (.I(\state[2] ),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _394_ (.A1(_064_),
    .A2(_065_),
    .A3(_370_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _395_ (.A1(_063_),
    .A2(_066_),
    .B(_054_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _396_ (.I(_067_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _397_ (.A1(_061_),
    .A2(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _398_ (.A1(\state[0] ),
    .A2(\state[1] ),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _399_ (.A1(_065_),
    .A2(net112),
    .A3(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _400_ (.I(net112),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _401_ (.A1(\state[0] ),
    .A2(\state[1] ),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _402_ (.A1(read_phase),
    .A2(_056_),
    .A3(_062_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _403_ (.A1(_072_),
    .A2(_073_),
    .B(_074_),
    .C(_065_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _404_ (.A1(_071_),
    .A2(_075_),
    .B(phase_complete),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _405_ (.I(net2),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _406_ (.A1(\state[1] ),
    .A2(\state[2] ),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _407_ (.A1(read_phase),
    .A2(_065_),
    .B1(_077_),
    .B2(_078_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _408_ (.I0(_062_),
    .I1(_070_),
    .S(_055_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _409_ (.I(read_phase),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _410_ (.I(\state[3] ),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _411_ (.A1(_056_),
    .A2(_079_),
    .B1(_080_),
    .B2(_081_),
    .C(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _412_ (.I0(net112),
    .I1(read_phase),
    .S(\state[2] ),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _413_ (.A1(_073_),
    .A2(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _414_ (.A1(\state[2] ),
    .A2(net112),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _415_ (.A1(_073_),
    .A2(_086_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _416_ (.A1(_085_),
    .A2(_087_),
    .B(_054_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _417_ (.A1(_076_),
    .A2(_083_),
    .A3(_088_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _418_ (.A1(_054_),
    .A2(_078_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _419_ (.A1(phase_complete),
    .A2(_057_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _420_ (.I(_091_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _421_ (.A1(_089_),
    .A2(_090_),
    .A3(_092_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _422_ (.A1(_082_),
    .A2(\state[2] ),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _423_ (.A1(_370_),
    .A2(_057_),
    .A3(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _424_ (.A1(_091_),
    .A2(_095_),
    .B(_090_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _425_ (.A1(_089_),
    .A2(_096_),
    .B(net74),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _426_ (.A1(net74),
    .A2(_069_),
    .A3(_093_),
    .B(_097_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _427_ (.A1(_095_),
    .A2(_061_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _428_ (.I0(_098_),
    .I1(_068_),
    .S(_362_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _429_ (.A1(\state[3] ),
    .A2(_078_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _430_ (.A1(_100_),
    .A2(_092_),
    .B(_089_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _431_ (.A1(_093_),
    .A2(_099_),
    .B1(_101_),
    .B2(_360_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _432_ (.A1(_063_),
    .A2(_066_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _433_ (.A1(_054_),
    .A2(_053_),
    .A3(_102_),
    .B1(_061_),
    .B2(_059_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _434_ (.A1(net76),
    .A2(_053_),
    .A3(_067_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _435_ (.A1(_370_),
    .A2(_057_),
    .A3(_094_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _436_ (.A1(_052_),
    .A2(_103_),
    .B(_104_),
    .C(_105_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _437_ (.A1(_059_),
    .A2(_058_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _438_ (.A1(_091_),
    .A2(_107_),
    .B(_090_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _439_ (.A1(_089_),
    .A2(_108_),
    .B(net76),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _440_ (.A1(_093_),
    .A2(_106_),
    .B(_109_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _441_ (.A1(net76),
    .A2(net74),
    .A3(net75),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _442_ (.A1(_051_),
    .A2(_110_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _443_ (.A1(net76),
    .A2(net74),
    .A3(net75),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _444_ (.A1(_051_),
    .A2(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _445_ (.A1(_061_),
    .A2(_113_),
    .B(_095_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _446_ (.A1(_067_),
    .A2(_111_),
    .B(_114_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _447_ (.A1(_051_),
    .A2(_101_),
    .B1(_115_),
    .B2(_093_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _448_ (.I(_054_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _449_ (.A1(_062_),
    .A2(_055_),
    .A3(_368_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _450_ (.A1(_367_),
    .A2(_063_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _451_ (.A1(_117_),
    .A2(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _452_ (.A1(net77),
    .A2(net76),
    .A3(_059_),
    .B(_058_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _453_ (.A1(_091_),
    .A2(_120_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _454_ (.A1(_100_),
    .A2(_121_),
    .B(_089_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _455_ (.A1(_116_),
    .A2(_093_),
    .A3(_119_),
    .B1(_122_),
    .B2(_365_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _456_ (.I(net35),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _457_ (.A1(_056_),
    .A2(\state[1] ),
    .A3(\state[2] ),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _458_ (.A1(net2),
    .A2(_124_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _459_ (.A1(_116_),
    .A2(_124_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _460_ (.A1(_123_),
    .A2(_125_),
    .B(_126_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _461_ (.I(_355_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _462_ (.A1(net60),
    .A2(net65),
    .A3(net66),
    .A4(_127_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _463_ (.A1(net51),
    .A2(net61),
    .A3(net62),
    .A4(net63),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _464_ (.A1(net56),
    .A2(net57),
    .A3(net58),
    .A4(net59),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _465_ (.A1(net52),
    .A2(net54),
    .A3(net55),
    .A4(_130_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _466_ (.A1(net70),
    .A2(net71),
    .A3(net72),
    .A4(net73),
    .Z(_132_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _467_ (.A1(net64),
    .A2(net67),
    .A3(net68),
    .A4(net69),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _468_ (.A1(net43),
    .A2(net47),
    .A3(net48),
    .A4(net49),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _469_ (.A1(net44),
    .A2(net45),
    .A3(net46),
    .A4(net50),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _470_ (.A1(_132_),
    .A2(_133_),
    .A3(_134_),
    .A4(_135_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _471_ (.A1(_128_),
    .A2(_129_),
    .A3(_131_),
    .A4(_136_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _472_ (.A1(_116_),
    .A2(net2),
    .B(_124_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _473_ (.A1(net36),
    .A2(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _474_ (.A1(_126_),
    .A2(_137_),
    .B(_139_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _475_ (.A1(_055_),
    .A2(_070_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _476_ (.A1(_054_),
    .A2(_140_),
    .Z(_141_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _477_ (.I(\state[0] ),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _478_ (.A1(_142_),
    .A2(\state[2] ),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _479_ (.A1(_072_),
    .A2(_073_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _480_ (.A1(_064_),
    .A2(net112),
    .B(_055_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _481_ (.I(phase_complete),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _482_ (.A1(_144_),
    .A2(_145_),
    .B(_081_),
    .C(_146_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _483_ (.A1(net11),
    .A2(net15),
    .A3(net18),
    .A4(net17),
    .Z(_148_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _484_ (.A1(net10),
    .A2(net13),
    .A3(net12),
    .A4(net16),
    .Z(_149_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _485_ (.A1(net20),
    .A2(net23),
    .A3(net27),
    .A4(net26),
    .Z(_150_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _486_ (.A1(net19),
    .A2(net22),
    .A3(net21),
    .A4(net24),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _487_ (.A1(_148_),
    .A2(_149_),
    .A3(_150_),
    .A4(_151_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _488_ (.A1(net30),
    .A2(net29),
    .A3(net32),
    .A4(net8),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _489_ (.A1(net14),
    .A2(net3),
    .A3(net28),
    .A4(net25),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _490_ (.A1(net31),
    .A2(net7),
    .A3(net6),
    .A4(net9),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _491_ (.A1(net34),
    .A2(net33),
    .A3(net5),
    .A4(net4),
    .Z(_156_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _492_ (.A1(_153_),
    .A2(_154_),
    .A3(_155_),
    .A4(_156_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _493_ (.A1(_152_),
    .A2(_157_),
    .B(_081_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _494_ (.A1(_143_),
    .A2(_147_),
    .B(\state[3] ),
    .C(_158_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _495_ (.A1(net11),
    .A2(net15),
    .A3(net18),
    .A4(net17),
    .Z(_160_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _496_ (.A1(net10),
    .A2(net13),
    .A3(net12),
    .A4(net16),
    .Z(_161_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _497_ (.A1(net20),
    .A2(net23),
    .A3(net27),
    .A4(net26),
    .Z(_162_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _498_ (.A1(net19),
    .A2(net22),
    .A3(net21),
    .A4(net24),
    .Z(_163_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _499_ (.A1(_160_),
    .A2(_161_),
    .A3(_162_),
    .A4(_163_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _500_ (.A1(net30),
    .A2(net29),
    .A3(net32),
    .A4(net8),
    .Z(_165_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _501_ (.A1(net14),
    .A2(net3),
    .A3(net28),
    .A4(net25),
    .Z(_166_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _502_ (.A1(net31),
    .A2(net7),
    .A3(net6),
    .A4(net9),
    .Z(_167_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _503_ (.A1(net34),
    .A2(net33),
    .A3(net5),
    .A4(net4),
    .Z(_168_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _504_ (.A1(_165_),
    .A2(_166_),
    .A3(_167_),
    .A4(_168_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _505_ (.A1(_164_),
    .A2(_169_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _506_ (.A1(_142_),
    .A2(_094_),
    .B1(_170_),
    .B2(read_phase),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _507_ (.A1(_141_),
    .A2(_159_),
    .A3(_171_),
    .Z(_172_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _508_ (.I(_172_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _509_ (.I(_173_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _510_ (.I0(net74),
    .I1(net37),
    .S(_174_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _511_ (.I0(net75),
    .I1(net38),
    .S(_173_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _512_ (.I0(net76),
    .I1(net39),
    .S(_173_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _513_ (.I0(net77),
    .I1(net40),
    .S(_173_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _514_ (.I0(net78),
    .I1(net41),
    .S(_173_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _515_ (.I(_173_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _516_ (.I(_159_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _517_ (.A1(_056_),
    .A2(_100_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _518_ (.A1(_064_),
    .A2(net2),
    .B(\state[2] ),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _519_ (.A1(_081_),
    .A2(_140_),
    .B1(_178_),
    .B2(_056_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _520_ (.A1(_170_),
    .A2(_177_),
    .B(_179_),
    .C(_082_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _521_ (.I(_180_),
    .Z(_181_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _522_ (.A1(_353_),
    .A2(_176_),
    .A3(_181_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _523_ (.A1(_353_),
    .A2(_175_),
    .B(_182_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _524_ (.A1(net64),
    .A2(net67),
    .A3(net68),
    .Z(_183_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _525_ (.A1(net70),
    .A2(net71),
    .Z(_184_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _526_ (.A1(_357_),
    .A2(net69),
    .A3(_183_),
    .A4(_184_),
    .Z(_185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _527_ (.A1(net72),
    .A2(net73),
    .Z(_186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _528_ (.A1(_185_),
    .A2(_186_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _529_ (.A1(_054_),
    .A2(_140_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _530_ (.I(_188_),
    .Z(_189_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _531_ (.A1(_189_),
    .A2(_187_),
    .Z(_190_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _532_ (.A1(_176_),
    .A2(_181_),
    .A3(_190_),
    .B(net43),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _533_ (.A1(net43),
    .A2(_175_),
    .A3(_187_),
    .B(_191_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _534_ (.A1(net42),
    .A2(net53),
    .Z(_192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _535_ (.A1(net69),
    .A2(net70),
    .Z(_193_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _536_ (.A1(net71),
    .A2(_183_),
    .A3(_192_),
    .A4(_193_),
    .Z(_194_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _537_ (.A1(net43),
    .A2(_186_),
    .A3(_194_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _538_ (.A1(_189_),
    .A2(_195_),
    .Z(_196_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _539_ (.A1(_176_),
    .A2(_181_),
    .A3(_196_),
    .B(net44),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _540_ (.A1(net44),
    .A2(_175_),
    .A3(_195_),
    .B(_197_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _541_ (.A1(net43),
    .A2(net44),
    .Z(_198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _542_ (.A1(_185_),
    .A2(_186_),
    .A3(_198_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _543_ (.A1(_189_),
    .A2(_199_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _544_ (.A1(_176_),
    .A2(_181_),
    .A3(_200_),
    .B(net45),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _545_ (.A1(net45),
    .A2(_175_),
    .A3(_199_),
    .B(_201_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _546_ (.A1(net45),
    .A2(_186_),
    .A3(_198_),
    .Z(_202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _547_ (.A1(_194_),
    .A2(_202_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _548_ (.A1(_189_),
    .A2(_203_),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _549_ (.A1(_176_),
    .A2(_181_),
    .A3(_204_),
    .B(net46),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _550_ (.A1(net46),
    .A2(_175_),
    .A3(_203_),
    .B(_205_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _551_ (.A1(net46),
    .A2(_185_),
    .A3(_202_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _552_ (.A1(_189_),
    .A2(_206_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _553_ (.A1(_176_),
    .A2(_181_),
    .A3(_207_),
    .B(net47),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _554_ (.A1(net47),
    .A2(_175_),
    .A3(_206_),
    .B(_208_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _555_ (.A1(net46),
    .A2(net47),
    .Z(_209_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _556_ (.A1(net45),
    .A2(_186_),
    .A3(_198_),
    .A4(_209_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _557_ (.A1(_194_),
    .A2(_210_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _558_ (.I(_159_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _559_ (.I(_180_),
    .Z(_213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _560_ (.A1(_189_),
    .A2(_211_),
    .Z(_214_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _561_ (.A1(_212_),
    .A2(_213_),
    .A3(_214_),
    .B(net48),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _562_ (.A1(net48),
    .A2(_175_),
    .A3(_211_),
    .B(_215_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _563_ (.A1(net45),
    .A2(net48),
    .A3(_209_),
    .Z(_216_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _564_ (.A1(_185_),
    .A2(_186_),
    .A3(_198_),
    .A4(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _565_ (.A1(_189_),
    .A2(_217_),
    .Z(_218_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _566_ (.A1(_212_),
    .A2(_213_),
    .A3(_218_),
    .B(net49),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _567_ (.A1(net49),
    .A2(_175_),
    .A3(_217_),
    .B(_219_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _568_ (.I(_173_),
    .Z(_220_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _569_ (.A1(net48),
    .A2(net49),
    .Z(_221_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _570_ (.A1(_194_),
    .A2(_210_),
    .A3(_221_),
    .Z(_222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _571_ (.I(_222_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _572_ (.I(_141_),
    .Z(_224_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _573_ (.A1(_224_),
    .A2(_222_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _574_ (.A1(_212_),
    .A2(_213_),
    .A3(_225_),
    .B(net50),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _575_ (.A1(net50),
    .A2(_220_),
    .A3(_223_),
    .B(_226_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _576_ (.A1(_185_),
    .A2(_210_),
    .Z(_227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _577_ (.A1(net50),
    .A2(_221_),
    .A3(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _578_ (.A1(net50),
    .A2(_221_),
    .Z(_229_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _579_ (.A1(_227_),
    .A2(_229_),
    .B(_224_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _580_ (.A1(_212_),
    .A2(_213_),
    .A3(_230_),
    .B(net51),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _581_ (.A1(net51),
    .A2(_220_),
    .A3(_228_),
    .B(_231_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _582_ (.A1(net50),
    .A2(net51),
    .Z(_232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _583_ (.A1(_222_),
    .A2(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _584_ (.A1(_222_),
    .A2(_232_),
    .B(_224_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _585_ (.A1(_212_),
    .A2(_213_),
    .A3(_234_),
    .B(net52),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _586_ (.A1(net52),
    .A2(_220_),
    .A3(_233_),
    .B(_235_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _587_ (.A1(_356_),
    .A2(_189_),
    .Z(_236_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _588_ (.A1(_159_),
    .A2(_180_),
    .Z(_237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _589_ (.I0(_236_),
    .I1(net53),
    .S(_237_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _590_ (.I(net54),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _591_ (.A1(net50),
    .A2(net51),
    .A3(net52),
    .Z(_239_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _592_ (.A1(_185_),
    .A2(_210_),
    .A3(_221_),
    .A4(_239_),
    .Z(_240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _593_ (.A1(_238_),
    .A2(_240_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _594_ (.A1(_224_),
    .A2(_240_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _595_ (.A1(_176_),
    .A2(_181_),
    .A3(_242_),
    .B(net54),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _596_ (.A1(_175_),
    .A2(_241_),
    .B(_243_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _597_ (.A1(_194_),
    .A2(_210_),
    .Z(_244_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _598_ (.A1(net54),
    .A2(_221_),
    .A3(_239_),
    .Z(_245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _599_ (.A1(_244_),
    .A2(_245_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _600_ (.A1(_244_),
    .A2(_245_),
    .B(_224_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _601_ (.A1(_212_),
    .A2(_213_),
    .A3(_247_),
    .B(net55),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _602_ (.A1(net55),
    .A2(_220_),
    .A3(_246_),
    .B(_248_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _603_ (.I(net56),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _604_ (.A1(net55),
    .A2(_185_),
    .A3(_210_),
    .A4(_245_),
    .Z(_250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _605_ (.A1(_249_),
    .A2(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _606_ (.A1(_224_),
    .A2(_250_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _607_ (.A1(_176_),
    .A2(_181_),
    .A3(_252_),
    .B(net56),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _608_ (.A1(_175_),
    .A2(_251_),
    .B(_253_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _609_ (.A1(net55),
    .A2(net56),
    .Z(_254_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _610_ (.A1(net54),
    .A2(_221_),
    .A3(_239_),
    .A4(_254_),
    .Z(_255_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _611_ (.A1(_194_),
    .A2(_210_),
    .A3(_255_),
    .Z(_256_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _612_ (.I(_256_),
    .Z(_257_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _613_ (.I(_257_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _614_ (.A1(_224_),
    .A2(_257_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _615_ (.A1(_212_),
    .A2(_213_),
    .A3(_259_),
    .B(net57),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _616_ (.A1(net57),
    .A2(_220_),
    .A3(_258_),
    .B(_260_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _617_ (.A1(_185_),
    .A2(_210_),
    .A3(_255_),
    .Z(_261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _618_ (.A1(net57),
    .A2(_261_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _619_ (.A1(net57),
    .A2(_261_),
    .B(_224_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _620_ (.A1(_212_),
    .A2(_213_),
    .A3(_263_),
    .B(net58),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _621_ (.A1(net58),
    .A2(_220_),
    .A3(_262_),
    .B(_264_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _622_ (.A1(net57),
    .A2(net58),
    .Z(_265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _623_ (.A1(_257_),
    .A2(_265_),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _624_ (.A1(_257_),
    .A2(_265_),
    .B(_141_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _625_ (.A1(_212_),
    .A2(_213_),
    .A3(_267_),
    .B(net59),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _626_ (.A1(net59),
    .A2(_220_),
    .A3(_266_),
    .B(_268_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _627_ (.A1(net59),
    .A2(_265_),
    .Z(_269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _628_ (.A1(_261_),
    .A2(_269_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _629_ (.A1(_261_),
    .A2(_269_),
    .B(_141_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _630_ (.A1(_212_),
    .A2(_213_),
    .A3(_271_),
    .B(net60),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _631_ (.A1(net60),
    .A2(_220_),
    .A3(_270_),
    .B(_272_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _632_ (.A1(net57),
    .A2(net58),
    .A3(net59),
    .A4(net60),
    .Z(_273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _633_ (.A1(_257_),
    .A2(_273_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _634_ (.I(_159_),
    .Z(_275_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _635_ (.I(_180_),
    .Z(_276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _636_ (.A1(_257_),
    .A2(_273_),
    .B(_141_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _637_ (.A1(_275_),
    .A2(_276_),
    .A3(_277_),
    .B(net61),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _638_ (.A1(net61),
    .A2(_220_),
    .A3(_274_),
    .B(_278_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _639_ (.A1(net61),
    .A2(_273_),
    .Z(_279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _640_ (.A1(_261_),
    .A2(_279_),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _641_ (.A1(_261_),
    .A2(_279_),
    .B(_141_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _642_ (.A1(_275_),
    .A2(_276_),
    .A3(_281_),
    .B(net62),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _643_ (.A1(net62),
    .A2(_220_),
    .A3(_280_),
    .B(_282_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _644_ (.A1(net61),
    .A2(net62),
    .A3(_273_),
    .Z(_283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _645_ (.A1(_257_),
    .A2(_283_),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _646_ (.A1(_257_),
    .A2(_283_),
    .B(_141_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _647_ (.A1(_275_),
    .A2(_276_),
    .A3(_285_),
    .B(net63),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _648_ (.A1(net63),
    .A2(_174_),
    .A3(_284_),
    .B(_286_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _649_ (.I(_357_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _650_ (.A1(_287_),
    .A2(_188_),
    .Z(_288_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _651_ (.A1(_275_),
    .A2(_276_),
    .A3(_288_),
    .B(net64),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _652_ (.A1(_287_),
    .A2(net64),
    .A3(_174_),
    .B(_289_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _653_ (.A1(net63),
    .A2(_283_),
    .Z(_290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _654_ (.A1(_261_),
    .A2(_290_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _655_ (.A1(_261_),
    .A2(_290_),
    .B(_141_),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _656_ (.A1(_275_),
    .A2(_276_),
    .A3(_292_),
    .B(net65),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _657_ (.A1(net65),
    .A2(_174_),
    .A3(_291_),
    .B(_293_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _658_ (.A1(net63),
    .A2(net65),
    .A3(_283_),
    .Z(_294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _659_ (.A1(_257_),
    .A2(_294_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _660_ (.A1(_257_),
    .A2(_294_),
    .B(_141_),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _661_ (.A1(_275_),
    .A2(_276_),
    .A3(_296_),
    .B(net66),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _662_ (.A1(net66),
    .A2(_174_),
    .A3(_295_),
    .B(_297_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _663_ (.A1(net64),
    .A2(_192_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _664_ (.A1(net67),
    .A2(_224_),
    .A3(_298_),
    .Z(_299_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _665_ (.A1(_176_),
    .A2(_181_),
    .B(net67),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _666_ (.A1(net67),
    .A2(_189_),
    .A3(_298_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _667_ (.A1(_237_),
    .A2(_299_),
    .B(_300_),
    .C(_301_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _668_ (.A1(_357_),
    .A2(net64),
    .A3(net67),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _669_ (.A1(net68),
    .A2(_224_),
    .A3(_302_),
    .Z(_303_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _670_ (.A1(_176_),
    .A2(_181_),
    .B(net68),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _671_ (.A1(net68),
    .A2(_189_),
    .A3(_302_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _672_ (.A1(_237_),
    .A2(_303_),
    .B(_304_),
    .C(_305_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _673_ (.A1(_183_),
    .A2(_192_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _674_ (.A1(_188_),
    .A2(_306_),
    .Z(_307_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _675_ (.A1(_275_),
    .A2(_276_),
    .A3(_307_),
    .B(net69),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _676_ (.A1(net69),
    .A2(_174_),
    .A3(_306_),
    .B(_308_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _677_ (.A1(_357_),
    .A2(net69),
    .A3(_183_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _678_ (.A1(_188_),
    .A2(_309_),
    .Z(_310_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _679_ (.A1(_275_),
    .A2(_276_),
    .A3(_310_),
    .B(net70),
    .ZN(_311_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _680_ (.A1(net70),
    .A2(_174_),
    .A3(_309_),
    .B(_311_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _681_ (.A1(_183_),
    .A2(_192_),
    .A3(_193_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _682_ (.A1(_188_),
    .A2(_312_),
    .Z(_313_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _683_ (.A1(_275_),
    .A2(_276_),
    .A3(_313_),
    .B(net71),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _684_ (.A1(net71),
    .A2(_174_),
    .A3(_312_),
    .B(_314_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _685_ (.I(_185_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _686_ (.A1(_188_),
    .A2(_315_),
    .Z(_316_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _687_ (.A1(_275_),
    .A2(_276_),
    .A3(_316_),
    .B(net72),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _688_ (.A1(net72),
    .A2(_174_),
    .A3(_315_),
    .B(_317_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _689_ (.A1(net72),
    .A2(_194_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _690_ (.A1(_188_),
    .A2(_318_),
    .Z(_319_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _691_ (.A1(_159_),
    .A2(_180_),
    .A3(_319_),
    .B(net73),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _692_ (.A1(net73),
    .A2(_174_),
    .A3(_318_),
    .B(_320_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _693_ (.I0(phase_complete),
    .I1(_072_),
    .S(_065_),
    .Z(_321_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _694_ (.A1(_062_),
    .A2(_086_),
    .B1(_321_),
    .B2(_056_),
    .C(_085_),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _695_ (.A1(_100_),
    .A2(_322_),
    .Z(_323_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _696_ (.A1(_076_),
    .A2(_083_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _697_ (.I0(phase_complete),
    .I1(_323_),
    .S(_324_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _698_ (.A1(net112),
    .A2(_070_),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _699_ (.A1(_065_),
    .A2(_325_),
    .B(_144_),
    .ZN(_326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _700_ (.A1(_142_),
    .A2(_178_),
    .Z(_327_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _701_ (.A1(_116_),
    .A2(phase_complete),
    .A3(_326_),
    .A4(_327_),
    .Z(_328_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _702_ (.A1(_116_),
    .A2(_327_),
    .B(read_phase),
    .ZN(_329_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _703_ (.A1(read_phase),
    .A2(_328_),
    .B(_329_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _704_ (.A1(\state[2] ),
    .A2(_370_),
    .B(phase_complete),
    .ZN(_330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _705_ (.A1(_062_),
    .A2(_330_),
    .Z(_331_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _706_ (.A1(_056_),
    .A2(_065_),
    .A3(_146_),
    .Z(_332_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _707_ (.A1(_077_),
    .A2(_124_),
    .Z(_333_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _708_ (.A1(_331_),
    .A2(_332_),
    .A3(_333_),
    .B(_082_),
    .ZN(_334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _709_ (.A1(phase_complete),
    .A2(_370_),
    .B(_054_),
    .C(_055_),
    .ZN(_335_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _710_ (.A1(_054_),
    .A2(_055_),
    .A3(net2),
    .Z(_336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _711_ (.A1(_335_),
    .A2(_336_),
    .B(_057_),
    .ZN(_337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _712_ (.A1(_061_),
    .A2(_334_),
    .A3(_337_),
    .ZN(_338_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _713_ (.A1(_116_),
    .A2(_338_),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _714_ (.I0(_338_),
    .I1(_339_),
    .S(_142_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _715_ (.A1(_142_),
    .A2(_082_),
    .Z(_340_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _716_ (.A1(_338_),
    .A2(_340_),
    .B(_062_),
    .ZN(_341_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _717_ (.A1(_142_),
    .A2(_062_),
    .A3(_116_),
    .A4(_338_),
    .Z(_342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _718_ (.A1(_341_),
    .A2(_342_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _719_ (.A1(_056_),
    .A2(_062_),
    .A3(_061_),
    .A4(_334_),
    .ZN(_343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _720_ (.I0(_073_),
    .I1(_343_),
    .S(_055_),
    .Z(_344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _721_ (.A1(_065_),
    .A2(_338_),
    .ZN(_345_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _722_ (.A1(_116_),
    .A2(_344_),
    .B(_345_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _723_ (.A1(_065_),
    .A2(_073_),
    .ZN(_346_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _724_ (.A1(_338_),
    .A2(_346_),
    .ZN(_347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _725_ (.I0(_125_),
    .I1(_347_),
    .S(_082_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _726_ (.A1(_062_),
    .A2(phase_complete),
    .ZN(_348_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _727_ (.A1(_327_),
    .A2(_348_),
    .Z(_349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _728_ (.A1(_081_),
    .A2(_346_),
    .B(_140_),
    .ZN(_350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _729_ (.A1(_065_),
    .A2(_073_),
    .B(_333_),
    .C(_116_),
    .ZN(_351_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _730_ (.A1(_116_),
    .A2(_349_),
    .A3(_350_),
    .B1(_351_),
    .B2(net112),
    .ZN(_352_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _731_ (.I(_352_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _732_ (.A1(_142_),
    .A2(_082_),
    .B(_078_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _733_ (.A1(_142_),
    .A2(_100_),
    .ZN(net104));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _734_ (.A(_353_),
    .B(_354_),
    .CO(_355_),
    .S(_356_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _735_ (.A(net42),
    .B(net53),
    .CO(_357_),
    .S(_358_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _736_ (.A(_359_),
    .B(_360_),
    .CO(_361_),
    .S(_362_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _737_ (.A(net74),
    .B(net75),
    .CO(_363_),
    .S(_364_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _738_ (.A(_365_),
    .B(_366_),
    .CO(_367_),
    .S(_368_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _739_ (.A(net78),
    .B(_369_),
    .CO(_370_),
    .S(_371_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _740_ (.I(net104),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _741_ (.I(net104),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _742_ (.I(net104),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _743_ (.I(net104),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _744_ (.I(net104),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _745_ (.I(net104),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _746_ (.I(net104),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _747_ (.I(net104),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _748_ (.I(net104),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _749_ (.I(net104),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _750_ (.I(net104),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _751_ (.I(net104),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _752_ (.I(net104),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _753_ (.I(net104),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _754_ (.I(net104),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _755_ (.I(net104),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _756_ (.I(net104),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _757_ (.I(net104),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _758_ (.I(net104),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _759_ (.I(net104),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _760_ (.I(net104),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _761_ (.I(net104),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _762_ (.I(net104),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _763_ (.I(net104),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _764_ (.I(net104),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _765_ (.I(net104),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _766_ (.I(net104),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _767_ (.I(net104),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _768_ (.I(net104),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _769_ (.I(net104),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _770_ (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \addr_counter[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \addr_counter[1]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \addr_counter[2]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net76));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \addr_counter[3]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net77));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \addr_counter[4]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net78));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bist_done$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net35));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bist_pass$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net36));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_addr[0]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_addr[1]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net38));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_addr[2]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net39));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_addr[3]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net40));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_addr[4]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[0]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[10]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[11]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net44));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[12]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[13]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[14]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[15]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[16]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[17]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[18]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[19]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[1]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[20]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[21]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[22]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[23]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[24]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[25]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[26]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[27]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[28]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[29]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[2]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[30]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[31]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[3]$_DFFE_PN0P_  (.D(_037_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[4]$_DFFE_PN0P_  (.D(_038_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[5]$_DFFE_PN0P_  (.D(_039_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[6]$_DFFE_PN0P_  (.D(_040_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[7]$_DFFE_PN0P_  (.D(_041_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[8]$_DFFE_PN0P_  (.D(_042_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error_count[9]$_DFFE_PN0P_  (.D(_043_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \phase_complete$_DFFE_PN0P_  (.D(_044_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(phase_complete));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \read_phase$_DFFE_PN0P_  (.D(_045_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(read_phase));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[0]$_DFFE_PN0P_  (.D(_046_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[1]$_DFFE_PN0P_  (.D(_047_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[2]$_DFFE_PN0P_  (.D(_048_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[3]$_DFFE_PN0P_  (.D(_049_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \write_phase$_DFFE_PN0P_  (.D(_050_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net113),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_90 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(bist_start),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(mem_rdata[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(mem_rdata[10]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(mem_rdata[11]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(mem_rdata[12]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(mem_rdata[13]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(mem_rdata[14]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(mem_rdata[15]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(mem_rdata[16]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(mem_rdata[17]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(mem_rdata[18]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(mem_rdata[19]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(mem_rdata[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(mem_rdata[20]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(mem_rdata[21]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(mem_rdata[22]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(mem_rdata[23]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(mem_rdata[24]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(mem_rdata[25]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(mem_rdata[26]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(mem_rdata[27]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(mem_rdata[28]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(mem_rdata[29]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(mem_rdata[2]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(mem_rdata[30]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(mem_rdata[31]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(mem_rdata[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(mem_rdata[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(mem_rdata[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(mem_rdata[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(mem_rdata[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(mem_rdata[8]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(mem_rdata[9]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output34 (.I(net35),
    .Z(bist_done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output35 (.I(net36),
    .Z(bist_pass));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output36 (.I(net37),
    .Z(error_addr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net38),
    .Z(error_addr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net39),
    .Z(error_addr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net40),
    .Z(error_addr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net41),
    .Z(error_addr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net42),
    .Z(error_count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net43),
    .Z(error_count[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net44),
    .Z(error_count[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net45),
    .Z(error_count[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net46),
    .Z(error_count[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net47),
    .Z(error_count[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net48),
    .Z(error_count[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net49),
    .Z(error_count[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net50),
    .Z(error_count[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net51),
    .Z(error_count[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net52),
    .Z(error_count[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net53),
    .Z(error_count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net54),
    .Z(error_count[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net55),
    .Z(error_count[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net56),
    .Z(error_count[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net57),
    .Z(error_count[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net58),
    .Z(error_count[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net59),
    .Z(error_count[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net60),
    .Z(error_count[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net61),
    .Z(error_count[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net62),
    .Z(error_count[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net63),
    .Z(error_count[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net64),
    .Z(error_count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net65),
    .Z(error_count[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net66),
    .Z(error_count[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net67),
    .Z(error_count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net68),
    .Z(error_count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net69),
    .Z(error_count[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(error_count[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(error_count[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net72),
    .Z(error_count[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net73),
    .Z(error_count[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net74),
    .Z(mem_addr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net75),
    .Z(mem_addr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net76),
    .Z(mem_addr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net77),
    .Z(mem_addr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net78),
    .Z(mem_addr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net79),
    .Z(mem_enable));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net80),
    .Z(mem_wdata[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net81),
    .Z(mem_wdata[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net82),
    .Z(mem_wdata[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net83),
    .Z(mem_wdata[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net84),
    .Z(mem_wdata[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net85),
    .Z(mem_wdata[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net86),
    .Z(mem_wdata[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net87),
    .Z(mem_wdata[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net88),
    .Z(mem_wdata[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net89),
    .Z(mem_wdata[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net90),
    .Z(mem_wdata[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net91),
    .Z(mem_wdata[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net92),
    .Z(mem_wdata[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net93),
    .Z(mem_wdata[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net94),
    .Z(mem_wdata[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net95),
    .Z(mem_wdata[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net96),
    .Z(mem_wdata[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net97),
    .Z(mem_wdata[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net98),
    .Z(mem_wdata[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net99),
    .Z(mem_wdata[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net100),
    .Z(mem_wdata[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net101),
    .Z(mem_wdata[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net102),
    .Z(mem_wdata[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net103),
    .Z(mem_wdata[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net104),
    .Z(mem_wdata[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net105),
    .Z(mem_wdata[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net106),
    .Z(mem_wdata[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net107),
    .Z(mem_wdata[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net108),
    .Z(mem_wdata[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net109),
    .Z(mem_wdata[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net110),
    .Z(mem_wdata[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net111),
    .Z(mem_wdata[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net112),
    .Z(mem_write));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload1 (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_374 ();
endmodule
