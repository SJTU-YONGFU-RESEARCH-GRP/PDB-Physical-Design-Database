module fixed_point_sqrt (clk,
    enable,
    reset,
    x,
    y);
 input clk;
 input enable;
 input reset;
 input [15:0] x;
 output [15:0] y;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _137_ (.A(reset),
    .Z(_068_));
 CLKBUF_X2 _138_ (.A(enable),
    .Z(_069_));
 INV_X1 _139_ (.A(_069_),
    .ZN(_070_));
 CLKBUF_X3 _140_ (.A(x[13]),
    .Z(_071_));
 BUF_X4 _141_ (.A(x[12]),
    .Z(_072_));
 NOR4_X4 _142_ (.A1(_071_),
    .A2(_072_),
    .A3(net1),
    .A4(net2),
    .ZN(_073_));
 NOR2_X1 _143_ (.A1(_070_),
    .A2(_073_),
    .ZN(_074_));
 AOI21_X1 _144_ (.A(_074_),
    .B1(_070_),
    .B2(net6),
    .ZN(_075_));
 NOR2_X1 _145_ (.A1(_068_),
    .A2(_075_),
    .ZN(_000_));
 CLKBUF_X3 _146_ (.A(x[8]),
    .Z(_076_));
 BUF_X2 _147_ (.A(x[0]),
    .Z(_077_));
 CLKBUF_X3 _148_ (.A(x[3]),
    .Z(_078_));
 BUF_X2 _149_ (.A(x[4]),
    .Z(_079_));
 NOR3_X2 _150_ (.A1(_077_),
    .A2(_078_),
    .A3(_079_),
    .ZN(_080_));
 CLKBUF_X3 _151_ (.A(x[1]),
    .Z(_081_));
 BUF_X2 _152_ (.A(x[2]),
    .Z(_082_));
 BUF_X2 _153_ (.A(x[5]),
    .Z(_083_));
 NOR3_X2 _154_ (.A1(_081_),
    .A2(_082_),
    .A3(_083_),
    .ZN(_084_));
 BUF_X2 _155_ (.A(x[6]),
    .Z(_085_));
 NOR3_X1 _156_ (.A1(net3),
    .A2(_085_),
    .A3(net4),
    .ZN(_086_));
 AND3_X1 _157_ (.A1(_080_),
    .A2(_084_),
    .A3(_086_),
    .ZN(_087_));
 CLKBUF_X3 _158_ (.A(x[10]),
    .Z(_088_));
 INV_X2 _159_ (.A(_088_),
    .ZN(_089_));
 CLKBUF_X3 _160_ (.A(x[11]),
    .Z(_090_));
 INV_X1 _161_ (.A(_090_),
    .ZN(_091_));
 AND3_X2 _162_ (.A1(_089_),
    .A2(_091_),
    .A3(_073_),
    .ZN(_092_));
 NAND3_X1 _163_ (.A1(_076_),
    .A2(_087_),
    .A3(_092_),
    .ZN(_093_));
 AND2_X1 _164_ (.A1(_069_),
    .A2(_093_),
    .ZN(_094_));
 NAND2_X2 _165_ (.A1(net3),
    .A2(net4),
    .ZN(_095_));
 NOR3_X1 _166_ (.A1(_085_),
    .A2(_076_),
    .A3(_095_),
    .ZN(_096_));
 NAND4_X2 _167_ (.A1(_080_),
    .A2(_084_),
    .A3(_092_),
    .A4(_096_),
    .ZN(_097_));
 NAND4_X1 _168_ (.A1(_079_),
    .A2(_072_),
    .A3(net1),
    .A4(net2),
    .ZN(_098_));
 NAND4_X1 _169_ (.A1(_076_),
    .A2(_088_),
    .A3(_090_),
    .A4(_071_),
    .ZN(_099_));
 OR2_X1 _170_ (.A1(_098_),
    .A2(_099_),
    .ZN(_100_));
 NAND2_X2 _171_ (.A1(_082_),
    .A2(_083_),
    .ZN(_101_));
 NAND4_X2 _172_ (.A1(_077_),
    .A2(_081_),
    .A3(_078_),
    .A4(_085_),
    .ZN(_102_));
 NOR4_X4 _173_ (.A1(_095_),
    .A2(_100_),
    .A3(_101_),
    .A4(_102_),
    .ZN(_103_));
 INV_X1 _174_ (.A(_103_),
    .ZN(_104_));
 NAND2_X2 _175_ (.A1(_097_),
    .A2(_104_),
    .ZN(_105_));
 AOI22_X1 _176_ (.A1(_070_),
    .A2(net8),
    .B1(_094_),
    .B2(_105_),
    .ZN(_106_));
 NOR2_X1 _177_ (.A1(_068_),
    .A2(_106_),
    .ZN(_001_));
 AOI22_X1 _178_ (.A1(_070_),
    .A2(net7),
    .B1(_094_),
    .B2(_103_),
    .ZN(_107_));
 NOR2_X1 _179_ (.A1(_068_),
    .A2(_107_),
    .ZN(_002_));
 NOR2_X1 _180_ (.A1(_082_),
    .A2(_083_),
    .ZN(_108_));
 OR2_X2 _181_ (.A1(net3),
    .A2(_085_),
    .ZN(_109_));
 INV_X1 _182_ (.A(net4),
    .ZN(_110_));
 INV_X1 _183_ (.A(_076_),
    .ZN(_111_));
 NAND3_X2 _184_ (.A1(_110_),
    .A2(_111_),
    .A3(_092_),
    .ZN(_112_));
 NOR3_X4 _185_ (.A1(_081_),
    .A2(_109_),
    .A3(_112_),
    .ZN(_113_));
 AND4_X1 _186_ (.A1(_077_),
    .A2(_078_),
    .A3(_108_),
    .A4(_113_),
    .ZN(_114_));
 OAI21_X1 _187_ (.A(_094_),
    .B1(_105_),
    .B2(_114_),
    .ZN(_115_));
 NAND2_X1 _188_ (.A1(_070_),
    .A2(net11),
    .ZN(_116_));
 AOI21_X1 _189_ (.A(_068_),
    .B1(_115_),
    .B2(_116_),
    .ZN(_003_));
 NOR2_X1 _190_ (.A1(_069_),
    .A2(_068_),
    .ZN(_117_));
 NAND2_X1 _191_ (.A1(net12),
    .A2(_117_),
    .ZN(_118_));
 INV_X1 _192_ (.A(_068_),
    .ZN(_119_));
 NAND2_X1 _193_ (.A1(_119_),
    .A2(_094_),
    .ZN(_120_));
 INV_X1 _194_ (.A(_112_),
    .ZN(_121_));
 NOR3_X2 _195_ (.A1(_078_),
    .A2(_079_),
    .A3(_101_),
    .ZN(_122_));
 NOR2_X1 _196_ (.A1(_081_),
    .A2(net3),
    .ZN(_123_));
 XOR2_X1 _197_ (.A(_077_),
    .B(_085_),
    .Z(_124_));
 NAND3_X1 _198_ (.A1(_122_),
    .A2(_123_),
    .A3(_124_),
    .ZN(_125_));
 INV_X1 _199_ (.A(_082_),
    .ZN(_126_));
 NOR4_X2 _200_ (.A1(_081_),
    .A2(_083_),
    .A3(_079_),
    .A4(_109_),
    .ZN(_009_));
 NAND4_X1 _201_ (.A1(_077_),
    .A2(_078_),
    .A3(_126_),
    .A4(_009_),
    .ZN(_010_));
 NOR2_X1 _202_ (.A1(_077_),
    .A2(_078_),
    .ZN(_011_));
 NAND3_X1 _203_ (.A1(_082_),
    .A2(_009_),
    .A3(_011_),
    .ZN(_012_));
 NAND3_X1 _204_ (.A1(_125_),
    .A2(_010_),
    .A3(_012_),
    .ZN(_013_));
 NOR2_X1 _205_ (.A1(_109_),
    .A2(_112_),
    .ZN(_014_));
 NOR2_X1 _206_ (.A1(net1),
    .A2(net2),
    .ZN(_015_));
 NAND2_X2 _207_ (.A1(_015_),
    .A2(_087_),
    .ZN(_016_));
 NOR2_X1 _208_ (.A1(_111_),
    .A2(_072_),
    .ZN(_017_));
 NOR3_X1 _209_ (.A1(_088_),
    .A2(_091_),
    .A3(_071_),
    .ZN(_018_));
 INV_X2 _210_ (.A(_071_),
    .ZN(_019_));
 NOR3_X2 _211_ (.A1(_089_),
    .A2(_090_),
    .A3(_019_),
    .ZN(_020_));
 OAI21_X2 _212_ (.A(_017_),
    .B1(_018_),
    .B2(_020_),
    .ZN(_021_));
 NOR4_X4 _213_ (.A1(_076_),
    .A2(_088_),
    .A3(_090_),
    .A4(_071_),
    .ZN(_022_));
 NOR4_X2 _214_ (.A1(_076_),
    .A2(_089_),
    .A3(_090_),
    .A4(_072_),
    .ZN(_023_));
 AOI22_X4 _215_ (.A1(_072_),
    .A2(_022_),
    .B1(_023_),
    .B2(_019_),
    .ZN(_024_));
 AOI21_X4 _216_ (.A(_016_),
    .B1(_021_),
    .B2(_024_),
    .ZN(_025_));
 INV_X1 _217_ (.A(_077_),
    .ZN(_026_));
 INV_X1 _218_ (.A(_078_),
    .ZN(_027_));
 AOI21_X1 _219_ (.A(_026_),
    .B1(_027_),
    .B2(_079_),
    .ZN(_028_));
 OAI21_X1 _220_ (.A(_108_),
    .B1(_011_),
    .B2(_028_),
    .ZN(_029_));
 INV_X1 _221_ (.A(_083_),
    .ZN(_030_));
 AOI22_X1 _222_ (.A1(_030_),
    .A2(_080_),
    .B1(_122_),
    .B2(_077_),
    .ZN(_031_));
 NAND2_X1 _223_ (.A1(_029_),
    .A2(_031_),
    .ZN(_032_));
 AOI21_X1 _224_ (.A(_025_),
    .B1(_032_),
    .B2(_113_),
    .ZN(_033_));
 AOI221_X2 _225_ (.A(_103_),
    .B1(_121_),
    .B2(_013_),
    .C1(_014_),
    .C2(_033_),
    .ZN(_034_));
 OAI21_X1 _226_ (.A(_118_),
    .B1(_120_),
    .B2(_034_),
    .ZN(_004_));
 INV_X1 _227_ (.A(net13),
    .ZN(_035_));
 NOR3_X1 _228_ (.A1(_105_),
    .A2(_121_),
    .A3(_025_),
    .ZN(_036_));
 AND2_X1 _229_ (.A1(_079_),
    .A2(_108_),
    .ZN(_037_));
 NAND2_X1 _230_ (.A1(_011_),
    .A2(_037_),
    .ZN(_038_));
 AOI21_X1 _231_ (.A(_122_),
    .B1(_037_),
    .B2(_078_),
    .ZN(_039_));
 OAI21_X1 _232_ (.A(_038_),
    .B1(_039_),
    .B2(_026_),
    .ZN(_040_));
 XNOR2_X1 _233_ (.A(_082_),
    .B(_083_),
    .ZN(_041_));
 NAND4_X1 _234_ (.A1(_085_),
    .A2(_080_),
    .A3(_123_),
    .A4(_041_),
    .ZN(_042_));
 NOR2_X1 _235_ (.A1(_112_),
    .A2(_042_),
    .ZN(_043_));
 AOI211_X2 _236_ (.A(_025_),
    .B(_043_),
    .C1(_032_),
    .C2(_113_),
    .ZN(_044_));
 AOI221_X2 _237_ (.A(_103_),
    .B1(_113_),
    .B2(_040_),
    .C1(_044_),
    .C2(_097_),
    .ZN(_045_));
 OAI33_X1 _238_ (.A1(_069_),
    .A2(_035_),
    .A3(_068_),
    .B1(_120_),
    .B2(_036_),
    .B3(_045_),
    .ZN(_005_));
 NAND2_X1 _239_ (.A1(net14),
    .A2(_117_),
    .ZN(_046_));
 OR2_X1 _240_ (.A1(net1),
    .A2(net2),
    .ZN(_047_));
 NOR2_X1 _241_ (.A1(_090_),
    .A2(_072_),
    .ZN(_048_));
 OAI21_X1 _242_ (.A(_088_),
    .B1(_076_),
    .B2(net4),
    .ZN(_049_));
 AOI21_X1 _243_ (.A(_019_),
    .B1(_048_),
    .B2(_049_),
    .ZN(_050_));
 NOR4_X1 _244_ (.A1(_047_),
    .A2(_014_),
    .A3(_025_),
    .A4(_050_),
    .ZN(_051_));
 NOR3_X1 _245_ (.A1(_105_),
    .A2(_043_),
    .A3(_051_),
    .ZN(_052_));
 OAI21_X1 _246_ (.A(_046_),
    .B1(_052_),
    .B2(_120_),
    .ZN(_006_));
 OAI21_X1 _247_ (.A(_119_),
    .B1(net15),
    .B2(_069_),
    .ZN(_053_));
 NAND2_X1 _248_ (.A1(_088_),
    .A2(_091_),
    .ZN(_054_));
 NAND3_X1 _249_ (.A1(_110_),
    .A2(_111_),
    .A3(_089_),
    .ZN(_055_));
 NAND4_X1 _250_ (.A1(_073_),
    .A2(_054_),
    .A3(_044_),
    .A4(_055_),
    .ZN(_056_));
 NOR2_X1 _251_ (.A1(_088_),
    .A2(_071_),
    .ZN(_057_));
 OAI21_X1 _252_ (.A(_017_),
    .B1(_057_),
    .B2(_020_),
    .ZN(_058_));
 OAI21_X1 _253_ (.A(_069_),
    .B1(_016_),
    .B2(_058_),
    .ZN(_059_));
 NOR2_X1 _254_ (.A1(_105_),
    .A2(_059_),
    .ZN(_060_));
 AOI21_X1 _255_ (.A(_053_),
    .B1(_056_),
    .B2(_060_),
    .ZN(_007_));
 NAND2_X1 _256_ (.A1(net16),
    .A2(_117_),
    .ZN(_061_));
 NOR3_X1 _257_ (.A1(_047_),
    .A2(_073_),
    .A3(_050_),
    .ZN(_062_));
 NOR3_X1 _258_ (.A1(_092_),
    .A2(_103_),
    .A3(_062_),
    .ZN(_063_));
 NAND3_X1 _259_ (.A1(_076_),
    .A2(_089_),
    .A3(_090_),
    .ZN(_064_));
 OAI21_X1 _260_ (.A(_064_),
    .B1(_054_),
    .B2(_076_),
    .ZN(_065_));
 AND2_X1 _261_ (.A1(_073_),
    .A2(_065_),
    .ZN(_066_));
 AOI221_X2 _262_ (.A(_103_),
    .B1(_044_),
    .B2(_063_),
    .C1(_066_),
    .C2(_087_),
    .ZN(_067_));
 OAI21_X1 _263_ (.A(_061_),
    .B1(_067_),
    .B2(_120_),
    .ZN(_008_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X1 _265_ (.A(net7),
    .Z(net5));
 BUF_X1 _266_ (.A(net7),
    .Z(net9));
 BUF_X1 _267_ (.A(net7),
    .Z(net10));
 BUF_X1 _268_ (.A(net17),
    .Z(y[12]));
 BUF_X1 _269_ (.A(net18),
    .Z(y[13]));
 BUF_X1 _270_ (.A(net19),
    .Z(y[14]));
 BUF_X1 _271_ (.A(net20),
    .Z(y[15]));
 DFF_X1 \y[10]$_SDFFE_PP0P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net6),
    .QN(_135_));
 DFF_X1 \y[1]$_SDFFE_PP0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net8),
    .QN(_134_));
 DFF_X1 \y[3]$_SDFFE_PP0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net7),
    .QN(_133_));
 DFF_X1 \y[4]$_SDFFE_PP0P_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net11),
    .QN(_132_));
 DFF_X1 \y[5]$_SDFFE_PP0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_131_));
 DFF_X1 \y[6]$_SDFFE_PP0P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_130_));
 DFF_X1 \y[7]$_SDFFE_PP0P_  (.D(_006_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_129_));
 DFF_X1 \y[8]$_SDFFE_PP0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_128_));
 DFF_X1 \y[9]$_SDFFE_PP0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_127_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_59 ();
 CLKBUF_X2 input1 (.A(x[14]),
    .Z(net1));
 CLKBUF_X2 input2 (.A(x[15]),
    .Z(net2));
 BUF_X1 input3 (.A(x[7]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(x[9]),
    .Z(net4));
 BUF_X1 output5 (.A(net5),
    .Z(y[0]));
 BUF_X1 output6 (.A(net6),
    .Z(y[10]));
 BUF_X1 output7 (.A(net7),
    .Z(y[11]));
 BUF_X1 output8 (.A(net8),
    .Z(y[1]));
 BUF_X1 output9 (.A(net9),
    .Z(y[2]));
 BUF_X1 output10 (.A(net10),
    .Z(y[3]));
 BUF_X1 output11 (.A(net11),
    .Z(y[4]));
 BUF_X1 output12 (.A(net12),
    .Z(y[5]));
 BUF_X1 output13 (.A(net13),
    .Z(y[6]));
 BUF_X1 output14 (.A(net14),
    .Z(y[7]));
 BUF_X1 output15 (.A(net15),
    .Z(y[8]));
 BUF_X1 output16 (.A(net16),
    .Z(y[9]));
 LOGIC0_X1 _268__17 (.Z(net17));
 LOGIC0_X1 _269__18 (.Z(net18));
 LOGIC0_X1 _270__19 (.Z(net19));
 LOGIC0_X1 _271__20 (.Z(net20));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X2 FILLER_0_73 ();
 FILLCELL_X1 FILLER_0_75 ();
 FILLCELL_X8 FILLER_0_80 ();
 FILLCELL_X16 FILLER_0_92 ();
 FILLCELL_X8 FILLER_0_108 ();
 FILLCELL_X4 FILLER_0_116 ();
 FILLCELL_X2 FILLER_0_120 ();
 FILLCELL_X16 FILLER_0_127 ();
 FILLCELL_X4 FILLER_0_143 ();
 FILLCELL_X2 FILLER_0_147 ();
 FILLCELL_X32 FILLER_0_154 ();
 FILLCELL_X32 FILLER_0_186 ();
 FILLCELL_X8 FILLER_0_218 ();
 FILLCELL_X2 FILLER_0_226 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_81 ();
 FILLCELL_X2 FILLER_1_89 ();
 FILLCELL_X1 FILLER_1_95 ();
 FILLCELL_X32 FILLER_1_103 ();
 FILLCELL_X32 FILLER_1_135 ();
 FILLCELL_X32 FILLER_1_167 ();
 FILLCELL_X16 FILLER_1_199 ();
 FILLCELL_X8 FILLER_1_215 ();
 FILLCELL_X4 FILLER_1_223 ();
 FILLCELL_X1 FILLER_1_227 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X16 FILLER_2_97 ();
 FILLCELL_X8 FILLER_2_113 ();
 FILLCELL_X4 FILLER_2_121 ();
 FILLCELL_X2 FILLER_2_125 ();
 FILLCELL_X1 FILLER_2_127 ();
 FILLCELL_X8 FILLER_2_130 ();
 FILLCELL_X4 FILLER_2_138 ();
 FILLCELL_X2 FILLER_2_142 ();
 FILLCELL_X32 FILLER_2_148 ();
 FILLCELL_X32 FILLER_2_180 ();
 FILLCELL_X16 FILLER_2_212 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X2 FILLER_3_97 ();
 FILLCELL_X1 FILLER_3_99 ();
 FILLCELL_X8 FILLER_3_111 ();
 FILLCELL_X32 FILLER_3_133 ();
 FILLCELL_X32 FILLER_3_165 ();
 FILLCELL_X16 FILLER_3_197 ();
 FILLCELL_X8 FILLER_3_213 ();
 FILLCELL_X4 FILLER_3_221 ();
 FILLCELL_X2 FILLER_3_225 ();
 FILLCELL_X1 FILLER_3_227 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X4 FILLER_4_97 ();
 FILLCELL_X2 FILLER_4_101 ();
 FILLCELL_X8 FILLER_4_110 ();
 FILLCELL_X4 FILLER_4_118 ();
 FILLCELL_X1 FILLER_4_122 ();
 FILLCELL_X32 FILLER_4_131 ();
 FILLCELL_X32 FILLER_4_163 ();
 FILLCELL_X32 FILLER_4_195 ();
 FILLCELL_X1 FILLER_4_227 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X2 FILLER_5_97 ();
 FILLCELL_X1 FILLER_5_99 ();
 FILLCELL_X8 FILLER_5_106 ();
 FILLCELL_X4 FILLER_5_114 ();
 FILLCELL_X2 FILLER_5_118 ();
 FILLCELL_X1 FILLER_5_120 ();
 FILLCELL_X32 FILLER_5_124 ();
 FILLCELL_X32 FILLER_5_156 ();
 FILLCELL_X32 FILLER_5_188 ();
 FILLCELL_X8 FILLER_5_220 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X4 FILLER_6_97 ();
 FILLCELL_X2 FILLER_6_101 ();
 FILLCELL_X1 FILLER_6_103 ();
 FILLCELL_X4 FILLER_6_109 ();
 FILLCELL_X1 FILLER_6_113 ();
 FILLCELL_X4 FILLER_6_116 ();
 FILLCELL_X2 FILLER_6_120 ();
 FILLCELL_X1 FILLER_6_122 ();
 FILLCELL_X32 FILLER_6_133 ();
 FILLCELL_X32 FILLER_6_165 ();
 FILLCELL_X16 FILLER_6_197 ();
 FILLCELL_X8 FILLER_6_213 ();
 FILLCELL_X4 FILLER_6_221 ();
 FILLCELL_X2 FILLER_6_225 ();
 FILLCELL_X1 FILLER_6_227 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X2 FILLER_7_89 ();
 FILLCELL_X1 FILLER_7_91 ();
 FILLCELL_X2 FILLER_7_97 ();
 FILLCELL_X4 FILLER_7_118 ();
 FILLCELL_X2 FILLER_7_122 ();
 FILLCELL_X4 FILLER_7_136 ();
 FILLCELL_X32 FILLER_7_142 ();
 FILLCELL_X32 FILLER_7_174 ();
 FILLCELL_X16 FILLER_7_206 ();
 FILLCELL_X4 FILLER_7_222 ();
 FILLCELL_X2 FILLER_7_226 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X1 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_105 ();
 FILLCELL_X4 FILLER_8_113 ();
 FILLCELL_X2 FILLER_8_117 ();
 FILLCELL_X4 FILLER_8_122 ();
 FILLCELL_X2 FILLER_8_126 ();
 FILLCELL_X1 FILLER_8_128 ();
 FILLCELL_X32 FILLER_8_135 ();
 FILLCELL_X32 FILLER_8_167 ();
 FILLCELL_X16 FILLER_8_199 ();
 FILLCELL_X8 FILLER_8_215 ();
 FILLCELL_X4 FILLER_8_223 ();
 FILLCELL_X1 FILLER_8_227 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X16 FILLER_9_108 ();
 FILLCELL_X1 FILLER_9_124 ();
 FILLCELL_X32 FILLER_9_131 ();
 FILLCELL_X32 FILLER_9_163 ();
 FILLCELL_X32 FILLER_9_195 ();
 FILLCELL_X1 FILLER_9_227 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X16 FILLER_10_65 ();
 FILLCELL_X8 FILLER_10_81 ();
 FILLCELL_X4 FILLER_10_89 ();
 FILLCELL_X8 FILLER_10_102 ();
 FILLCELL_X4 FILLER_10_110 ();
 FILLCELL_X2 FILLER_10_114 ();
 FILLCELL_X1 FILLER_10_116 ();
 FILLCELL_X32 FILLER_10_131 ();
 FILLCELL_X32 FILLER_10_163 ();
 FILLCELL_X32 FILLER_10_195 ();
 FILLCELL_X1 FILLER_10_227 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X1 FILLER_11_13 ();
 FILLCELL_X32 FILLER_11_19 ();
 FILLCELL_X32 FILLER_11_51 ();
 FILLCELL_X8 FILLER_11_83 ();
 FILLCELL_X2 FILLER_11_91 ();
 FILLCELL_X1 FILLER_11_93 ();
 FILLCELL_X4 FILLER_11_103 ();
 FILLCELL_X32 FILLER_11_113 ();
 FILLCELL_X32 FILLER_11_145 ();
 FILLCELL_X32 FILLER_11_177 ();
 FILLCELL_X16 FILLER_11_209 ();
 FILLCELL_X2 FILLER_11_225 ();
 FILLCELL_X1 FILLER_11_227 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_5 ();
 FILLCELL_X16 FILLER_12_14 ();
 FILLCELL_X4 FILLER_12_30 ();
 FILLCELL_X16 FILLER_12_38 ();
 FILLCELL_X4 FILLER_12_54 ();
 FILLCELL_X2 FILLER_12_58 ();
 FILLCELL_X16 FILLER_12_69 ();
 FILLCELL_X2 FILLER_12_85 ();
 FILLCELL_X2 FILLER_12_94 ();
 FILLCELL_X16 FILLER_12_105 ();
 FILLCELL_X4 FILLER_12_121 ();
 FILLCELL_X2 FILLER_12_125 ();
 FILLCELL_X4 FILLER_12_129 ();
 FILLCELL_X8 FILLER_12_144 ();
 FILLCELL_X4 FILLER_12_152 ();
 FILLCELL_X2 FILLER_12_156 ();
 FILLCELL_X8 FILLER_12_175 ();
 FILLCELL_X4 FILLER_12_183 ();
 FILLCELL_X2 FILLER_12_187 ();
 FILLCELL_X1 FILLER_12_189 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X2 FILLER_12_225 ();
 FILLCELL_X1 FILLER_12_227 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_9 ();
 FILLCELL_X1 FILLER_13_11 ();
 FILLCELL_X4 FILLER_13_16 ();
 FILLCELL_X16 FILLER_13_24 ();
 FILLCELL_X4 FILLER_13_40 ();
 FILLCELL_X8 FILLER_13_48 ();
 FILLCELL_X2 FILLER_13_74 ();
 FILLCELL_X1 FILLER_13_78 ();
 FILLCELL_X2 FILLER_13_86 ();
 FILLCELL_X1 FILLER_13_88 ();
 FILLCELL_X4 FILLER_13_91 ();
 FILLCELL_X2 FILLER_13_95 ();
 FILLCELL_X16 FILLER_13_102 ();
 FILLCELL_X1 FILLER_13_118 ();
 FILLCELL_X1 FILLER_13_123 ();
 FILLCELL_X16 FILLER_13_139 ();
 FILLCELL_X4 FILLER_13_155 ();
 FILLCELL_X2 FILLER_13_159 ();
 FILLCELL_X4 FILLER_13_165 ();
 FILLCELL_X1 FILLER_13_169 ();
 FILLCELL_X2 FILLER_13_180 ();
 FILLCELL_X1 FILLER_13_182 ();
 FILLCELL_X4 FILLER_13_200 ();
 FILLCELL_X1 FILLER_13_204 ();
 FILLCELL_X16 FILLER_13_208 ();
 FILLCELL_X4 FILLER_13_224 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_33 ();
 FILLCELL_X8 FILLER_14_53 ();
 FILLCELL_X16 FILLER_14_66 ();
 FILLCELL_X4 FILLER_14_82 ();
 FILLCELL_X1 FILLER_14_86 ();
 FILLCELL_X1 FILLER_14_96 ();
 FILLCELL_X16 FILLER_14_101 ();
 FILLCELL_X2 FILLER_14_117 ();
 FILLCELL_X1 FILLER_14_119 ();
 FILLCELL_X2 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_142 ();
 FILLCELL_X1 FILLER_14_174 ();
 FILLCELL_X32 FILLER_14_183 ();
 FILLCELL_X8 FILLER_14_215 ();
 FILLCELL_X4 FILLER_14_223 ();
 FILLCELL_X1 FILLER_14_227 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_33 ();
 FILLCELL_X2 FILLER_15_55 ();
 FILLCELL_X1 FILLER_15_57 ();
 FILLCELL_X16 FILLER_15_61 ();
 FILLCELL_X4 FILLER_15_77 ();
 FILLCELL_X2 FILLER_15_81 ();
 FILLCELL_X1 FILLER_15_83 ();
 FILLCELL_X4 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_105 ();
 FILLCELL_X4 FILLER_15_137 ();
 FILLCELL_X4 FILLER_15_170 ();
 FILLCELL_X1 FILLER_15_174 ();
 FILLCELL_X8 FILLER_15_178 ();
 FILLCELL_X2 FILLER_15_186 ();
 FILLCELL_X1 FILLER_15_188 ();
 FILLCELL_X32 FILLER_15_192 ();
 FILLCELL_X4 FILLER_15_224 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_33 ();
 FILLCELL_X1 FILLER_16_56 ();
 FILLCELL_X16 FILLER_16_64 ();
 FILLCELL_X8 FILLER_16_80 ();
 FILLCELL_X4 FILLER_16_88 ();
 FILLCELL_X4 FILLER_16_101 ();
 FILLCELL_X1 FILLER_16_105 ();
 FILLCELL_X16 FILLER_16_117 ();
 FILLCELL_X8 FILLER_16_133 ();
 FILLCELL_X4 FILLER_16_141 ();
 FILLCELL_X16 FILLER_16_147 ();
 FILLCELL_X4 FILLER_16_163 ();
 FILLCELL_X2 FILLER_16_167 ();
 FILLCELL_X1 FILLER_16_169 ();
 FILLCELL_X4 FILLER_16_191 ();
 FILLCELL_X2 FILLER_16_195 ();
 FILLCELL_X1 FILLER_16_197 ();
 FILLCELL_X16 FILLER_16_201 ();
 FILLCELL_X8 FILLER_16_217 ();
 FILLCELL_X2 FILLER_16_225 ();
 FILLCELL_X1 FILLER_16_227 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_17 ();
 FILLCELL_X8 FILLER_17_28 ();
 FILLCELL_X4 FILLER_17_36 ();
 FILLCELL_X1 FILLER_17_40 ();
 FILLCELL_X1 FILLER_17_44 ();
 FILLCELL_X1 FILLER_17_52 ();
 FILLCELL_X2 FILLER_17_57 ();
 FILLCELL_X4 FILLER_17_63 ();
 FILLCELL_X1 FILLER_17_67 ();
 FILLCELL_X2 FILLER_17_74 ();
 FILLCELL_X1 FILLER_17_79 ();
 FILLCELL_X2 FILLER_17_86 ();
 FILLCELL_X1 FILLER_17_88 ();
 FILLCELL_X4 FILLER_17_93 ();
 FILLCELL_X2 FILLER_17_97 ();
 FILLCELL_X4 FILLER_17_103 ();
 FILLCELL_X1 FILLER_17_107 ();
 FILLCELL_X4 FILLER_17_112 ();
 FILLCELL_X2 FILLER_17_116 ();
 FILLCELL_X8 FILLER_17_149 ();
 FILLCELL_X4 FILLER_17_157 ();
 FILLCELL_X1 FILLER_17_161 ();
 FILLCELL_X16 FILLER_17_167 ();
 FILLCELL_X4 FILLER_17_183 ();
 FILLCELL_X2 FILLER_17_187 ();
 FILLCELL_X32 FILLER_17_192 ();
 FILLCELL_X4 FILLER_17_224 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_33 ();
 FILLCELL_X1 FILLER_18_37 ();
 FILLCELL_X32 FILLER_18_43 ();
 FILLCELL_X32 FILLER_18_75 ();
 FILLCELL_X16 FILLER_18_107 ();
 FILLCELL_X2 FILLER_18_123 ();
 FILLCELL_X4 FILLER_18_129 ();
 FILLCELL_X2 FILLER_18_133 ();
 FILLCELL_X1 FILLER_18_135 ();
 FILLCELL_X32 FILLER_18_138 ();
 FILLCELL_X16 FILLER_18_170 ();
 FILLCELL_X4 FILLER_18_186 ();
 FILLCELL_X2 FILLER_18_190 ();
 FILLCELL_X32 FILLER_18_196 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X4 FILLER_19_113 ();
 FILLCELL_X8 FILLER_19_120 ();
 FILLCELL_X4 FILLER_19_128 ();
 FILLCELL_X2 FILLER_19_132 ();
 FILLCELL_X1 FILLER_19_134 ();
 FILLCELL_X8 FILLER_19_139 ();
 FILLCELL_X4 FILLER_19_147 ();
 FILLCELL_X4 FILLER_19_156 ();
 FILLCELL_X1 FILLER_19_160 ();
 FILLCELL_X2 FILLER_19_164 ();
 FILLCELL_X32 FILLER_19_183 ();
 FILLCELL_X2 FILLER_19_215 ();
 FILLCELL_X1 FILLER_19_223 ();
 FILLCELL_X1 FILLER_19_227 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X2 FILLER_20_113 ();
 FILLCELL_X1 FILLER_20_115 ();
 FILLCELL_X1 FILLER_20_120 ();
 FILLCELL_X8 FILLER_20_141 ();
 FILLCELL_X2 FILLER_20_149 ();
 FILLCELL_X2 FILLER_20_156 ();
 FILLCELL_X1 FILLER_20_158 ();
 FILLCELL_X32 FILLER_20_179 ();
 FILLCELL_X4 FILLER_20_211 ();
 FILLCELL_X2 FILLER_20_215 ();
 FILLCELL_X2 FILLER_20_220 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X8 FILLER_21_129 ();
 FILLCELL_X2 FILLER_21_137 ();
 FILLCELL_X1 FILLER_21_139 ();
 FILLCELL_X1 FILLER_21_147 ();
 FILLCELL_X32 FILLER_21_153 ();
 FILLCELL_X8 FILLER_21_185 ();
 FILLCELL_X2 FILLER_21_193 ();
 FILLCELL_X1 FILLER_21_195 ();
 FILLCELL_X16 FILLER_21_199 ();
 FILLCELL_X4 FILLER_21_215 ();
 FILLCELL_X1 FILLER_21_219 ();
 FILLCELL_X4 FILLER_21_223 ();
 FILLCELL_X1 FILLER_21_227 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X4 FILLER_22_129 ();
 FILLCELL_X1 FILLER_22_133 ();
 FILLCELL_X32 FILLER_22_151 ();
 FILLCELL_X32 FILLER_22_183 ();
 FILLCELL_X8 FILLER_22_215 ();
 FILLCELL_X4 FILLER_22_223 ();
 FILLCELL_X1 FILLER_22_227 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X2 FILLER_23_225 ();
 FILLCELL_X1 FILLER_23_227 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X2 FILLER_24_225 ();
 FILLCELL_X1 FILLER_24_227 ();
 FILLCELL_X2 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_10 ();
 FILLCELL_X32 FILLER_25_42 ();
 FILLCELL_X32 FILLER_25_74 ();
 FILLCELL_X16 FILLER_25_106 ();
 FILLCELL_X4 FILLER_25_122 ();
 FILLCELL_X2 FILLER_25_126 ();
 FILLCELL_X1 FILLER_25_128 ();
 FILLCELL_X32 FILLER_25_133 ();
 FILLCELL_X32 FILLER_25_165 ();
 FILLCELL_X16 FILLER_25_197 ();
 FILLCELL_X8 FILLER_25_213 ();
 FILLCELL_X4 FILLER_25_221 ();
 FILLCELL_X2 FILLER_25_225 ();
 FILLCELL_X1 FILLER_25_227 ();
 FILLCELL_X2 FILLER_26_12 ();
 FILLCELL_X32 FILLER_26_16 ();
 FILLCELL_X32 FILLER_26_48 ();
 FILLCELL_X32 FILLER_26_80 ();
 FILLCELL_X32 FILLER_26_112 ();
 FILLCELL_X32 FILLER_26_144 ();
 FILLCELL_X32 FILLER_26_176 ();
 FILLCELL_X16 FILLER_26_208 ();
 FILLCELL_X4 FILLER_26_224 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X2 FILLER_27_225 ();
 FILLCELL_X1 FILLER_27_227 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X2 FILLER_28_225 ();
 FILLCELL_X1 FILLER_28_227 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X16 FILLER_29_97 ();
 FILLCELL_X8 FILLER_29_113 ();
 FILLCELL_X16 FILLER_29_124 ();
 FILLCELL_X8 FILLER_29_140 ();
 FILLCELL_X32 FILLER_29_151 ();
 FILLCELL_X32 FILLER_29_183 ();
 FILLCELL_X8 FILLER_29_215 ();
 FILLCELL_X4 FILLER_29_223 ();
 FILLCELL_X1 FILLER_29_227 ();
endmodule
