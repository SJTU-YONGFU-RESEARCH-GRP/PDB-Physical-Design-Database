module simple_spi (ack_o,
    clk_i,
    cyc_i,
    inta_o,
    miso_i,
    mosi_o,
    rst_i,
    sck_o,
    stb_i,
    we_i,
    adr_i,
    dat_i,
    dat_o);
 output ack_o;
 input clk_i;
 input cyc_i;
 output inta_o;
 input miso_i;
 output mosi_o;
 input rst_i;
 output sck_o;
 input stb_i;
 input we_i;
 input [1:0] adr_i;
 input [7:0] dat_i;
 output [7:0] dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire \bcnt[0] ;
 wire \bcnt[1] ;
 wire \bcnt[2] ;
 wire \clkcnt[0] ;
 wire \clkcnt[10] ;
 wire \clkcnt[11] ;
 wire \clkcnt[1] ;
 wire \clkcnt[2] ;
 wire \clkcnt[3] ;
 wire \clkcnt[4] ;
 wire \clkcnt[5] ;
 wire \clkcnt[6] ;
 wire \clkcnt[7] ;
 wire \clkcnt[8] ;
 wire \clkcnt[9] ;
 wire cpha;
 wire cpol;
 wire dwom;
 wire \espr[0] ;
 wire \espr[1] ;
 wire \espr[2] ;
 wire \espr[3] ;
 wire \icnt[0] ;
 wire \icnt[1] ;
 wire \rfifo.din[1] ;
 wire \rfifo.din[2] ;
 wire \rfifo.din[3] ;
 wire \rfifo.din[4] ;
 wire \rfifo.din[5] ;
 wire \rfifo.din[6] ;
 wire \rfifo.din[7] ;
 wire \rfifo.gb ;
 wire \rfifo.mem[0][0] ;
 wire \rfifo.mem[0][1] ;
 wire \rfifo.mem[0][2] ;
 wire \rfifo.mem[0][3] ;
 wire \rfifo.mem[0][4] ;
 wire \rfifo.mem[0][5] ;
 wire \rfifo.mem[0][6] ;
 wire \rfifo.mem[0][7] ;
 wire \rfifo.mem[1][0] ;
 wire \rfifo.mem[1][1] ;
 wire \rfifo.mem[1][2] ;
 wire \rfifo.mem[1][3] ;
 wire \rfifo.mem[1][4] ;
 wire \rfifo.mem[1][5] ;
 wire \rfifo.mem[1][6] ;
 wire \rfifo.mem[1][7] ;
 wire \rfifo.mem[2][0] ;
 wire \rfifo.mem[2][1] ;
 wire \rfifo.mem[2][2] ;
 wire \rfifo.mem[2][3] ;
 wire \rfifo.mem[2][4] ;
 wire \rfifo.mem[2][5] ;
 wire \rfifo.mem[2][6] ;
 wire \rfifo.mem[2][7] ;
 wire \rfifo.mem[3][0] ;
 wire \rfifo.mem[3][1] ;
 wire \rfifo.mem[3][2] ;
 wire \rfifo.mem[3][3] ;
 wire \rfifo.mem[3][4] ;
 wire \rfifo.mem[3][5] ;
 wire \rfifo.mem[3][6] ;
 wire \rfifo.mem[3][7] ;
 wire \rfifo.rp[0] ;
 wire \rfifo.rp[1] ;
 wire \rfifo.we ;
 wire \rfifo.wp[0] ;
 wire \rfifo.wp[1] ;
 wire spe;
 wire \sper[2] ;
 wire \sper[3] ;
 wire \sper[4] ;
 wire \sper[5] ;
 wire spie;
 wire spif;
 wire \state[0] ;
 wire \state[1] ;
 wire \tcnt[0] ;
 wire \tcnt[1] ;
 wire wcol;
 wire \wfifo.gb ;
 wire \wfifo.mem[0][0] ;
 wire \wfifo.mem[0][1] ;
 wire \wfifo.mem[0][2] ;
 wire \wfifo.mem[0][3] ;
 wire \wfifo.mem[0][4] ;
 wire \wfifo.mem[0][5] ;
 wire \wfifo.mem[0][6] ;
 wire \wfifo.mem[0][7] ;
 wire \wfifo.mem[1][0] ;
 wire \wfifo.mem[1][1] ;
 wire \wfifo.mem[1][2] ;
 wire \wfifo.mem[1][3] ;
 wire \wfifo.mem[1][4] ;
 wire \wfifo.mem[1][5] ;
 wire \wfifo.mem[1][6] ;
 wire \wfifo.mem[1][7] ;
 wire \wfifo.mem[2][0] ;
 wire \wfifo.mem[2][1] ;
 wire \wfifo.mem[2][2] ;
 wire \wfifo.mem[2][3] ;
 wire \wfifo.mem[2][4] ;
 wire \wfifo.mem[2][5] ;
 wire \wfifo.mem[2][6] ;
 wire \wfifo.mem[2][7] ;
 wire \wfifo.mem[3][0] ;
 wire \wfifo.mem[3][1] ;
 wire \wfifo.mem[3][2] ;
 wire \wfifo.mem[3][3] ;
 wire \wfifo.mem[3][4] ;
 wire \wfifo.mem[3][5] ;
 wire \wfifo.mem[3][6] ;
 wire \wfifo.mem[3][7] ;
 wire \wfifo.re ;
 wire \wfifo.rp[0] ;
 wire \wfifo.rp[1] ;
 wire \wfifo.wp[0] ;
 wire \wfifo.wp[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire clknet_0_clk_i;
 wire clknet_4_0_0_clk_i;
 wire clknet_4_1_0_clk_i;
 wire clknet_4_2_0_clk_i;
 wire clknet_4_3_0_clk_i;
 wire clknet_4_4_0_clk_i;
 wire clknet_4_5_0_clk_i;
 wire clknet_4_6_0_clk_i;
 wire clknet_4_7_0_clk_i;
 wire clknet_4_8_0_clk_i;
 wire clknet_4_9_0_clk_i;
 wire clknet_4_10_0_clk_i;
 wire clknet_4_11_0_clk_i;
 wire clknet_4_12_0_clk_i;
 wire clknet_4_13_0_clk_i;
 wire clknet_4_14_0_clk_i;
 wire clknet_4_15_0_clk_i;
 wire net29;
 wire net30;

 BUF_X4 _0615_ (.A(adr_i[0]),
    .Z(_0130_));
 INV_X2 _0616_ (.A(_0130_),
    .ZN(_0131_));
 CLKBUF_X3 _0617_ (.A(\rfifo.rp[1] ),
    .Z(_0132_));
 CLKBUF_X3 _0618_ (.A(_0132_),
    .Z(_0133_));
 MUX2_X1 _0619_ (.A(\rfifo.mem[0][0] ),
    .B(\rfifo.mem[2][0] ),
    .S(_0133_),
    .Z(_0134_));
 MUX2_X1 _0620_ (.A(\rfifo.mem[1][0] ),
    .B(\rfifo.mem[3][0] ),
    .S(_0133_),
    .Z(_0135_));
 BUF_X2 _0621_ (.A(\rfifo.rp[0] ),
    .Z(_0136_));
 CLKBUF_X3 _0622_ (.A(_0136_),
    .Z(_0137_));
 MUX2_X1 _0623_ (.A(_0134_),
    .B(_0135_),
    .S(_0137_),
    .Z(_0138_));
 CLKBUF_X3 _0624_ (.A(adr_i[1]),
    .Z(_0139_));
 CLKBUF_X3 _0625_ (.A(_0139_),
    .Z(_0140_));
 MUX2_X1 _0626_ (.A(\espr[0] ),
    .B(_0138_),
    .S(_0140_),
    .Z(_0141_));
 NAND2_X1 _0627_ (.A1(_0131_),
    .A2(_0141_),
    .ZN(_0142_));
 BUF_X1 _0628_ (.A(\espr[2] ),
    .Z(_0143_));
 CLKBUF_X3 _0629_ (.A(_0143_),
    .Z(_0144_));
 INV_X1 _0630_ (.A(\rfifo.gb ),
    .ZN(_0145_));
 XOR2_X1 _0631_ (.A(_0133_),
    .B(\rfifo.wp[1] ),
    .Z(_0146_));
 XOR2_X2 _0632_ (.A(\rfifo.wp[0] ),
    .B(_0136_),
    .Z(_0147_));
 NOR3_X1 _0633_ (.A1(_0139_),
    .A2(_0146_),
    .A3(_0147_),
    .ZN(_0148_));
 AOI22_X1 _0634_ (.A1(_0140_),
    .A2(_0144_),
    .B1(_0145_),
    .B2(_0148_),
    .ZN(_0149_));
 OAI21_X1 _0635_ (.A(_0142_),
    .B1(_0149_),
    .B2(_0131_),
    .ZN(_0453_));
 BUF_X2 _0636_ (.A(\espr[3] ),
    .Z(_0150_));
 AOI221_X1 _0637_ (.A(_0131_),
    .B1(_0139_),
    .B2(_0150_),
    .C1(\rfifo.gb ),
    .C2(_0148_),
    .ZN(_0151_));
 MUX2_X1 _0638_ (.A(\rfifo.mem[0][1] ),
    .B(\rfifo.mem[2][1] ),
    .S(_0133_),
    .Z(_0152_));
 MUX2_X1 _0639_ (.A(\rfifo.mem[1][1] ),
    .B(\rfifo.mem[3][1] ),
    .S(_0133_),
    .Z(_0153_));
 MUX2_X1 _0640_ (.A(_0152_),
    .B(_0153_),
    .S(_0137_),
    .Z(_0154_));
 AND2_X1 _0641_ (.A1(_0140_),
    .A2(_0154_),
    .ZN(_0155_));
 BUF_X2 _0642_ (.A(\espr[1] ),
    .Z(_0156_));
 INV_X2 _0643_ (.A(_0139_),
    .ZN(_0157_));
 AOI21_X1 _0644_ (.A(_0155_),
    .B1(_0156_),
    .B2(_0157_),
    .ZN(_0158_));
 AOI21_X1 _0645_ (.A(_0151_),
    .B1(_0158_),
    .B2(_0131_),
    .ZN(_0454_));
 MUX2_X1 _0646_ (.A(\rfifo.mem[0][2] ),
    .B(\rfifo.mem[2][2] ),
    .S(_0132_),
    .Z(_0159_));
 MUX2_X1 _0647_ (.A(\rfifo.mem[1][2] ),
    .B(\rfifo.mem[3][2] ),
    .S(_0132_),
    .Z(_0160_));
 MUX2_X1 _0648_ (.A(_0159_),
    .B(_0160_),
    .S(_0137_),
    .Z(_0161_));
 MUX2_X1 _0649_ (.A(cpha),
    .B(_0161_),
    .S(_0140_),
    .Z(_0162_));
 XNOR2_X2 _0650_ (.A(\wfifo.rp[0] ),
    .B(\wfifo.wp[0] ),
    .ZN(_0163_));
 CLKBUF_X3 _0651_ (.A(\wfifo.rp[1] ),
    .Z(_0164_));
 XNOR2_X2 _0652_ (.A(\wfifo.wp[1] ),
    .B(_0164_),
    .ZN(_0165_));
 AND3_X1 _0653_ (.A1(_0002_),
    .A2(_0163_),
    .A3(_0165_),
    .ZN(_0166_));
 MUX2_X1 _0654_ (.A(\sper[2] ),
    .B(_0166_),
    .S(_0157_),
    .Z(_0167_));
 MUX2_X1 _0655_ (.A(_0162_),
    .B(_0167_),
    .S(_0130_),
    .Z(_0455_));
 MUX2_X1 _0656_ (.A(\rfifo.mem[0][3] ),
    .B(\rfifo.mem[2][3] ),
    .S(_0132_),
    .Z(_0168_));
 MUX2_X1 _0657_ (.A(\rfifo.mem[1][3] ),
    .B(\rfifo.mem[3][3] ),
    .S(_0132_),
    .Z(_0169_));
 MUX2_X1 _0658_ (.A(_0168_),
    .B(_0169_),
    .S(_0137_),
    .Z(_0170_));
 MUX2_X1 _0659_ (.A(cpol),
    .B(_0170_),
    .S(_0140_),
    .Z(_0171_));
 NAND2_X1 _0660_ (.A1(_0163_),
    .A2(_0165_),
    .ZN(_0172_));
 NOR2_X1 _0661_ (.A1(_0002_),
    .A2(_0172_),
    .ZN(_0173_));
 MUX2_X1 _0662_ (.A(\sper[3] ),
    .B(_0173_),
    .S(_0157_),
    .Z(_0174_));
 MUX2_X1 _0663_ (.A(_0171_),
    .B(_0174_),
    .S(_0130_),
    .Z(_0456_));
 MUX2_X1 _0664_ (.A(\rfifo.mem[0][4] ),
    .B(\rfifo.mem[2][4] ),
    .S(_0133_),
    .Z(_0175_));
 MUX2_X1 _0665_ (.A(\rfifo.mem[1][4] ),
    .B(\rfifo.mem[3][4] ),
    .S(_0133_),
    .Z(_0176_));
 MUX2_X1 _0666_ (.A(_0175_),
    .B(_0176_),
    .S(_0137_),
    .Z(_0177_));
 OAI21_X1 _0667_ (.A(_0131_),
    .B1(_0157_),
    .B2(_0177_),
    .ZN(_0178_));
 NAND3_X1 _0668_ (.A1(_0130_),
    .A2(_0140_),
    .A3(\sper[4] ),
    .ZN(_0179_));
 NAND2_X1 _0669_ (.A1(_0178_),
    .A2(_0179_),
    .ZN(_0457_));
 NAND3_X1 _0670_ (.A1(_0130_),
    .A2(_0140_),
    .A3(\sper[5] ),
    .ZN(_0180_));
 MUX2_X1 _0671_ (.A(\rfifo.mem[0][5] ),
    .B(\rfifo.mem[2][5] ),
    .S(_0133_),
    .Z(_0181_));
 MUX2_X1 _0672_ (.A(\rfifo.mem[1][5] ),
    .B(\rfifo.mem[3][5] ),
    .S(_0133_),
    .Z(_0182_));
 MUX2_X1 _0673_ (.A(_0181_),
    .B(_0182_),
    .S(_0137_),
    .Z(_0183_));
 AND2_X1 _0674_ (.A1(_0140_),
    .A2(_0183_),
    .ZN(_0184_));
 AOI21_X1 _0675_ (.A(_0184_),
    .B1(dwom),
    .B2(_0157_),
    .ZN(_0185_));
 OAI21_X1 _0676_ (.A(_0180_),
    .B1(_0185_),
    .B2(_0130_),
    .ZN(_0458_));
 BUF_X1 _0677_ (.A(spe),
    .Z(_0186_));
 MUX2_X1 _0678_ (.A(\rfifo.mem[0][6] ),
    .B(\rfifo.mem[2][6] ),
    .S(_0132_),
    .Z(_0187_));
 MUX2_X1 _0679_ (.A(\rfifo.mem[1][6] ),
    .B(\rfifo.mem[3][6] ),
    .S(_0132_),
    .Z(_0188_));
 MUX2_X1 _0680_ (.A(_0187_),
    .B(_0188_),
    .S(_0136_),
    .Z(_0189_));
 MUX2_X1 _0681_ (.A(_0186_),
    .B(_0189_),
    .S(_0139_),
    .Z(_0190_));
 MUX2_X1 _0682_ (.A(wcol),
    .B(\icnt[0] ),
    .S(_0140_),
    .Z(_0191_));
 MUX2_X1 _0683_ (.A(_0190_),
    .B(_0191_),
    .S(_0130_),
    .Z(_0459_));
 MUX2_X1 _0684_ (.A(\rfifo.mem[0][7] ),
    .B(\rfifo.mem[2][7] ),
    .S(_0132_),
    .Z(_0192_));
 MUX2_X1 _0685_ (.A(\rfifo.mem[1][7] ),
    .B(\rfifo.mem[3][7] ),
    .S(_0132_),
    .Z(_0193_));
 MUX2_X1 _0686_ (.A(_0192_),
    .B(_0193_),
    .S(_0136_),
    .Z(_0194_));
 MUX2_X1 _0687_ (.A(spie),
    .B(_0194_),
    .S(_0139_),
    .Z(_0195_));
 MUX2_X1 _0688_ (.A(spif),
    .B(\icnt[1] ),
    .S(_0140_),
    .Z(_0196_));
 MUX2_X1 _0689_ (.A(_0195_),
    .B(_0196_),
    .S(_0130_),
    .Z(_0460_));
 AND3_X1 _0690_ (.A1(net15),
    .A2(net6),
    .A3(_0004_),
    .ZN(_0000_));
 AND2_X1 _0691_ (.A1(spif),
    .A2(spie),
    .ZN(_0001_));
 BUF_X2 _0692_ (.A(_0596_),
    .Z(_0197_));
 NOR2_X2 _0693_ (.A1(_0005_),
    .A2(_0197_),
    .ZN(_0198_));
 INV_X1 _0694_ (.A(\clkcnt[11] ),
    .ZN(_0199_));
 NOR3_X4 _0695_ (.A1(\clkcnt[9] ),
    .A2(\clkcnt[8] ),
    .A3(\clkcnt[10] ),
    .ZN(_0200_));
 NAND3_X2 _0696_ (.A1(_0199_),
    .A2(_0604_),
    .A3(_0200_),
    .ZN(_0201_));
 BUF_X2 _0697_ (.A(\clkcnt[2] ),
    .Z(_0202_));
 BUF_X2 _0698_ (.A(\clkcnt[4] ),
    .Z(_0203_));
 NOR4_X4 _0699_ (.A1(\clkcnt[3] ),
    .A2(_0202_),
    .A3(\clkcnt[5] ),
    .A4(_0203_),
    .ZN(_0204_));
 NOR2_X1 _0700_ (.A1(\clkcnt[7] ),
    .A2(\clkcnt[6] ),
    .ZN(_0205_));
 NAND2_X2 _0701_ (.A1(_0204_),
    .A2(_0205_),
    .ZN(_0206_));
 OAI21_X2 _0702_ (.A(_0198_),
    .B1(_0201_),
    .B2(_0206_),
    .ZN(_0207_));
 BUF_X2 _0703_ (.A(_0207_),
    .Z(_0208_));
 OR2_X1 _0704_ (.A1(_0150_),
    .A2(_0144_),
    .ZN(_0209_));
 OR2_X1 _0705_ (.A1(_0156_),
    .A2(\espr[0] ),
    .ZN(_0210_));
 NAND2_X2 _0706_ (.A1(_0150_),
    .A2(_0143_),
    .ZN(_0211_));
 OAI221_X1 _0707_ (.A(_0208_),
    .B1(_0209_),
    .B2(_0210_),
    .C1(_0211_),
    .C2(\clkcnt[0] ),
    .ZN(_0212_));
 INV_X1 _0708_ (.A(_0602_),
    .ZN(_0213_));
 OAI21_X1 _0709_ (.A(_0212_),
    .B1(_0208_),
    .B2(_0213_),
    .ZN(_0012_));
 AND2_X1 _0710_ (.A1(_0156_),
    .A2(\espr[0] ),
    .ZN(_0214_));
 OAI21_X1 _0711_ (.A(_0150_),
    .B1(_0143_),
    .B2(_0214_),
    .ZN(_0215_));
 BUF_X2 _0712_ (.A(_0606_),
    .Z(_0216_));
 AND2_X2 _0713_ (.A1(_0204_),
    .A2(_0205_),
    .ZN(_0217_));
 AND2_X1 _0714_ (.A1(_0216_),
    .A2(_0217_),
    .ZN(_0218_));
 NOR2_X1 _0715_ (.A1(\clkcnt[9] ),
    .A2(\clkcnt[8] ),
    .ZN(_0219_));
 AND3_X1 _0716_ (.A1(_0143_),
    .A2(_0219_),
    .A3(_0198_),
    .ZN(_0220_));
 INV_X1 _0717_ (.A(\clkcnt[10] ),
    .ZN(_0221_));
 AOI221_X1 _0718_ (.A(_0215_),
    .B1(_0218_),
    .B2(_0220_),
    .C1(_0144_),
    .C2(_0221_),
    .ZN(_0222_));
 NAND3_X1 _0719_ (.A1(_0216_),
    .A2(_0217_),
    .A3(_0219_),
    .ZN(_0223_));
 XNOR2_X1 _0720_ (.A(\clkcnt[10] ),
    .B(_0223_),
    .ZN(_0224_));
 INV_X2 _0721_ (.A(_0198_),
    .ZN(_0225_));
 AND3_X2 _0722_ (.A1(_0199_),
    .A2(_0604_),
    .A3(_0200_),
    .ZN(_0226_));
 AOI21_X4 _0723_ (.A(_0225_),
    .B1(_0226_),
    .B2(_0217_),
    .ZN(_0227_));
 BUF_X4 _0724_ (.A(_0227_),
    .Z(_0228_));
 MUX2_X1 _0725_ (.A(_0222_),
    .B(_0224_),
    .S(_0228_),
    .Z(_0013_));
 CLKBUF_X2 _0726_ (.A(\clkcnt[1] ),
    .Z(_0229_));
 NOR4_X2 _0727_ (.A1(\clkcnt[7] ),
    .A2(\clkcnt[6] ),
    .A3(_0229_),
    .A4(\clkcnt[0] ),
    .ZN(_0230_));
 NAND3_X1 _0728_ (.A1(_0204_),
    .A2(_0200_),
    .A3(_0230_),
    .ZN(_0231_));
 OR3_X1 _0729_ (.A1(\clkcnt[11] ),
    .A2(_0208_),
    .A3(_0231_),
    .ZN(_0232_));
 NAND3_X1 _0730_ (.A1(\clkcnt[11] ),
    .A2(_0198_),
    .A3(_0231_),
    .ZN(_0233_));
 AND2_X1 _0731_ (.A1(_0150_),
    .A2(_0143_),
    .ZN(_0234_));
 NAND3_X1 _0732_ (.A1(\clkcnt[11] ),
    .A2(_0225_),
    .A3(_0234_),
    .ZN(_0235_));
 NAND3_X1 _0733_ (.A1(_0232_),
    .A2(_0233_),
    .A3(_0235_),
    .ZN(_0014_));
 OAI221_X1 _0734_ (.A(_0208_),
    .B1(_0209_),
    .B2(_0156_),
    .C1(_0211_),
    .C2(_0229_),
    .ZN(_0236_));
 OAI21_X1 _0735_ (.A(_0236_),
    .B1(_0208_),
    .B2(_0605_),
    .ZN(_0015_));
 NOR3_X1 _0736_ (.A1(_0228_),
    .A2(_0209_),
    .A3(_0214_),
    .ZN(_0237_));
 AND3_X1 _0737_ (.A1(_0202_),
    .A2(_0216_),
    .A3(_0228_),
    .ZN(_0238_));
 NOR3_X1 _0738_ (.A1(_0202_),
    .A2(_0228_),
    .A3(_0211_),
    .ZN(_0239_));
 NOR3_X1 _0739_ (.A1(_0202_),
    .A2(_0216_),
    .A3(_0207_),
    .ZN(_0240_));
 NOR4_X1 _0740_ (.A1(_0237_),
    .A2(_0238_),
    .A3(_0239_),
    .A4(_0240_),
    .ZN(_0016_));
 INV_X1 _0741_ (.A(\clkcnt[3] ),
    .ZN(_0241_));
 OR3_X1 _0742_ (.A1(_0202_),
    .A2(_0229_),
    .A3(\clkcnt[0] ),
    .ZN(_0242_));
 NOR3_X1 _0743_ (.A1(_0241_),
    .A2(_0207_),
    .A3(_0242_),
    .ZN(_0243_));
 MUX2_X1 _0744_ (.A(_0234_),
    .B(_0242_),
    .S(_0227_),
    .Z(_0244_));
 INV_X1 _0745_ (.A(\espr[0] ),
    .ZN(_0245_));
 AOI21_X1 _0746_ (.A(_0214_),
    .B1(_0144_),
    .B2(_0245_),
    .ZN(_0246_));
 NOR2_X2 _0747_ (.A1(_0150_),
    .A2(_0227_),
    .ZN(_0247_));
 AOI221_X1 _0748_ (.A(_0243_),
    .B1(_0244_),
    .B2(_0241_),
    .C1(_0246_),
    .C2(_0247_),
    .ZN(_0017_));
 INV_X1 _0749_ (.A(_0150_),
    .ZN(_0248_));
 OAI21_X1 _0750_ (.A(_0144_),
    .B1(_0245_),
    .B2(_0156_),
    .ZN(_0249_));
 NAND2_X1 _0751_ (.A1(_0248_),
    .A2(_0249_),
    .ZN(_0250_));
 NOR2_X2 _0752_ (.A1(_0206_),
    .A2(_0201_),
    .ZN(_0251_));
 OAI221_X1 _0753_ (.A(_0250_),
    .B1(_0225_),
    .B2(_0251_),
    .C1(_0203_),
    .C2(_0211_),
    .ZN(_0252_));
 NOR2_X1 _0754_ (.A1(\clkcnt[3] ),
    .A2(_0202_),
    .ZN(_0253_));
 NAND2_X1 _0755_ (.A1(_0216_),
    .A2(_0253_),
    .ZN(_0254_));
 XOR2_X1 _0756_ (.A(_0203_),
    .B(_0254_),
    .Z(_0255_));
 OAI21_X1 _0757_ (.A(_0252_),
    .B1(_0255_),
    .B2(_0208_),
    .ZN(_0018_));
 INV_X1 _0758_ (.A(\clkcnt[5] ),
    .ZN(_0256_));
 NOR2_X1 _0759_ (.A1(_0203_),
    .A2(_0229_),
    .ZN(_0257_));
 NAND3_X1 _0760_ (.A1(_0602_),
    .A2(_0253_),
    .A3(_0257_),
    .ZN(_0258_));
 NOR3_X1 _0761_ (.A1(_0256_),
    .A2(_0207_),
    .A3(_0258_),
    .ZN(_0259_));
 MUX2_X1 _0762_ (.A(_0234_),
    .B(_0258_),
    .S(_0227_),
    .Z(_0260_));
 NAND2_X1 _0763_ (.A1(_0156_),
    .A2(_0144_),
    .ZN(_0261_));
 AOI221_X1 _0764_ (.A(_0259_),
    .B1(_0260_),
    .B2(_0256_),
    .C1(_0247_),
    .C2(_0261_),
    .ZN(_0019_));
 INV_X1 _0765_ (.A(\clkcnt[6] ),
    .ZN(_0262_));
 NAND2_X1 _0766_ (.A1(_0216_),
    .A2(_0204_),
    .ZN(_0263_));
 NOR3_X1 _0767_ (.A1(_0262_),
    .A2(_0225_),
    .A3(_0263_),
    .ZN(_0264_));
 NAND2_X1 _0768_ (.A1(_0144_),
    .A2(_0214_),
    .ZN(_0265_));
 MUX2_X1 _0769_ (.A(_0234_),
    .B(_0263_),
    .S(_0228_),
    .Z(_0266_));
 AOI221_X1 _0770_ (.A(_0264_),
    .B1(_0265_),
    .B2(_0247_),
    .C1(_0266_),
    .C2(_0262_),
    .ZN(_0020_));
 INV_X1 _0771_ (.A(\clkcnt[7] ),
    .ZN(_0267_));
 NOR3_X1 _0772_ (.A1(\clkcnt[6] ),
    .A2(_0229_),
    .A3(\clkcnt[0] ),
    .ZN(_0268_));
 NAND2_X1 _0773_ (.A1(_0204_),
    .A2(_0268_),
    .ZN(_0269_));
 NOR2_X1 _0774_ (.A1(_0267_),
    .A2(_0269_),
    .ZN(_0270_));
 MUX2_X1 _0775_ (.A(_0144_),
    .B(_0269_),
    .S(_0228_),
    .Z(_0271_));
 AOI221_X1 _0776_ (.A(_0247_),
    .B1(_0270_),
    .B2(_0228_),
    .C1(_0271_),
    .C2(_0267_),
    .ZN(_0021_));
 NOR2_X1 _0777_ (.A1(_0248_),
    .A2(_0144_),
    .ZN(_0272_));
 NAND3_X1 _0778_ (.A1(_0208_),
    .A2(_0210_),
    .A3(_0272_),
    .ZN(_0273_));
 INV_X1 _0779_ (.A(\clkcnt[8] ),
    .ZN(_0274_));
 NAND2_X1 _0780_ (.A1(_0274_),
    .A2(_0228_),
    .ZN(_0275_));
 NAND2_X1 _0781_ (.A1(_0216_),
    .A2(_0217_),
    .ZN(_0276_));
 MUX2_X1 _0782_ (.A(_0211_),
    .B(_0218_),
    .S(_0228_),
    .Z(_0277_));
 OAI221_X1 _0783_ (.A(_0273_),
    .B1(_0275_),
    .B2(_0276_),
    .C1(_0277_),
    .C2(_0274_),
    .ZN(_0022_));
 NAND3_X1 _0784_ (.A1(_0156_),
    .A2(_0208_),
    .A3(_0272_),
    .ZN(_0278_));
 NAND3_X1 _0785_ (.A1(\clkcnt[9] ),
    .A2(_0208_),
    .A3(_0234_),
    .ZN(_0279_));
 NAND2_X1 _0786_ (.A1(_0204_),
    .A2(_0230_),
    .ZN(_0280_));
 OAI21_X1 _0787_ (.A(\clkcnt[9] ),
    .B1(\clkcnt[8] ),
    .B2(_0280_),
    .ZN(_0281_));
 OR2_X1 _0788_ (.A1(_0208_),
    .A2(_0281_),
    .ZN(_0282_));
 NAND4_X1 _0789_ (.A1(_0204_),
    .A2(_0219_),
    .A3(_0228_),
    .A4(_0230_),
    .ZN(_0283_));
 NAND4_X1 _0790_ (.A1(_0278_),
    .A2(_0279_),
    .A3(_0282_),
    .A4(_0283_),
    .ZN(_0023_));
 BUF_X1 _0791_ (.A(\rfifo.din[1] ),
    .Z(_0284_));
 BUF_X4 _0792_ (.A(\rfifo.we ),
    .Z(_0285_));
 NAND2_X4 _0793_ (.A1(_0285_),
    .A2(_0576_),
    .ZN(_0286_));
 MUX2_X1 _0794_ (.A(_0284_),
    .B(\rfifo.mem[0][0] ),
    .S(_0286_),
    .Z(_0025_));
 CLKBUF_X2 _0795_ (.A(\rfifo.din[2] ),
    .Z(_0287_));
 MUX2_X1 _0796_ (.A(_0287_),
    .B(\rfifo.mem[0][1] ),
    .S(_0286_),
    .Z(_0026_));
 BUF_X1 _0797_ (.A(\rfifo.din[3] ),
    .Z(_0288_));
 MUX2_X1 _0798_ (.A(_0288_),
    .B(\rfifo.mem[0][2] ),
    .S(_0286_),
    .Z(_0027_));
 BUF_X1 _0799_ (.A(\rfifo.din[4] ),
    .Z(_0289_));
 MUX2_X1 _0800_ (.A(_0289_),
    .B(\rfifo.mem[0][3] ),
    .S(_0286_),
    .Z(_0028_));
 BUF_X1 _0801_ (.A(\rfifo.din[5] ),
    .Z(_0290_));
 MUX2_X1 _0802_ (.A(_0290_),
    .B(\rfifo.mem[0][4] ),
    .S(_0286_),
    .Z(_0029_));
 BUF_X1 _0803_ (.A(\rfifo.din[6] ),
    .Z(_0291_));
 MUX2_X1 _0804_ (.A(_0291_),
    .B(\rfifo.mem[0][5] ),
    .S(_0286_),
    .Z(_0030_));
 BUF_X1 _0805_ (.A(\rfifo.din[7] ),
    .Z(_0292_));
 MUX2_X1 _0806_ (.A(_0292_),
    .B(\rfifo.mem[0][6] ),
    .S(_0286_),
    .Z(_0031_));
 MUX2_X1 _0807_ (.A(net27),
    .B(\rfifo.mem[0][7] ),
    .S(_0286_),
    .Z(_0032_));
 NAND2_X4 _0808_ (.A1(_0285_),
    .A2(_0580_),
    .ZN(_0293_));
 MUX2_X1 _0809_ (.A(_0284_),
    .B(\rfifo.mem[1][0] ),
    .S(_0293_),
    .Z(_0033_));
 MUX2_X1 _0810_ (.A(_0287_),
    .B(\rfifo.mem[1][1] ),
    .S(_0293_),
    .Z(_0034_));
 MUX2_X1 _0811_ (.A(_0288_),
    .B(\rfifo.mem[1][2] ),
    .S(_0293_),
    .Z(_0035_));
 MUX2_X1 _0812_ (.A(_0289_),
    .B(\rfifo.mem[1][3] ),
    .S(_0293_),
    .Z(_0036_));
 MUX2_X1 _0813_ (.A(_0290_),
    .B(\rfifo.mem[1][4] ),
    .S(_0293_),
    .Z(_0037_));
 MUX2_X1 _0814_ (.A(_0291_),
    .B(\rfifo.mem[1][5] ),
    .S(_0293_),
    .Z(_0038_));
 MUX2_X1 _0815_ (.A(_0292_),
    .B(\rfifo.mem[1][6] ),
    .S(_0293_),
    .Z(_0039_));
 MUX2_X1 _0816_ (.A(net27),
    .B(\rfifo.mem[1][7] ),
    .S(_0293_),
    .Z(_0040_));
 NAND2_X4 _0817_ (.A1(_0285_),
    .A2(_0578_),
    .ZN(_0294_));
 MUX2_X1 _0818_ (.A(_0284_),
    .B(\rfifo.mem[2][0] ),
    .S(_0294_),
    .Z(_0041_));
 MUX2_X1 _0819_ (.A(_0287_),
    .B(\rfifo.mem[2][1] ),
    .S(_0294_),
    .Z(_0042_));
 MUX2_X1 _0820_ (.A(_0288_),
    .B(\rfifo.mem[2][2] ),
    .S(_0294_),
    .Z(_0043_));
 MUX2_X1 _0821_ (.A(_0289_),
    .B(\rfifo.mem[2][3] ),
    .S(_0294_),
    .Z(_0044_));
 MUX2_X1 _0822_ (.A(_0290_),
    .B(\rfifo.mem[2][4] ),
    .S(_0294_),
    .Z(_0045_));
 MUX2_X1 _0823_ (.A(_0291_),
    .B(\rfifo.mem[2][5] ),
    .S(_0294_),
    .Z(_0046_));
 MUX2_X1 _0824_ (.A(_0292_),
    .B(\rfifo.mem[2][6] ),
    .S(_0294_),
    .Z(_0047_));
 MUX2_X1 _0825_ (.A(net27),
    .B(\rfifo.mem[2][7] ),
    .S(_0294_),
    .Z(_0048_));
 NAND2_X4 _0826_ (.A1(_0285_),
    .A2(_0582_),
    .ZN(_0295_));
 MUX2_X1 _0827_ (.A(_0284_),
    .B(\rfifo.mem[3][0] ),
    .S(_0295_),
    .Z(_0049_));
 MUX2_X1 _0828_ (.A(_0287_),
    .B(\rfifo.mem[3][1] ),
    .S(_0295_),
    .Z(_0050_));
 MUX2_X1 _0829_ (.A(_0288_),
    .B(\rfifo.mem[3][2] ),
    .S(_0295_),
    .Z(_0051_));
 MUX2_X1 _0830_ (.A(_0289_),
    .B(\rfifo.mem[3][3] ),
    .S(_0295_),
    .Z(_0052_));
 MUX2_X1 _0831_ (.A(_0290_),
    .B(\rfifo.mem[3][4] ),
    .S(_0295_),
    .Z(_0053_));
 MUX2_X1 _0832_ (.A(_0291_),
    .B(\rfifo.mem[3][5] ),
    .S(_0295_),
    .Z(_0054_));
 MUX2_X1 _0833_ (.A(_0292_),
    .B(\rfifo.mem[3][6] ),
    .S(_0295_),
    .Z(_0055_));
 MUX2_X1 _0834_ (.A(net27),
    .B(\rfifo.mem[3][7] ),
    .S(_0295_),
    .Z(_0056_));
 INV_X1 _0835_ (.A(_0186_),
    .ZN(_0296_));
 CLKBUF_X3 _0836_ (.A(_0296_),
    .Z(_0297_));
 NOR2_X1 _0837_ (.A1(_0297_),
    .A2(_0137_),
    .ZN(_0298_));
 INV_X1 _0838_ (.A(_0005_),
    .ZN(_0299_));
 OR3_X2 _0839_ (.A1(_0130_),
    .A2(_0157_),
    .A3(_0004_),
    .ZN(_0300_));
 INV_X1 _0840_ (.A(net16),
    .ZN(_0301_));
 NAND3_X1 _0841_ (.A1(net15),
    .A2(net6),
    .A3(_0301_),
    .ZN(_0302_));
 OAI21_X2 _0842_ (.A(_0299_),
    .B1(_0300_),
    .B2(_0302_),
    .ZN(_0303_));
 MUX2_X1 _0843_ (.A(_0137_),
    .B(_0298_),
    .S(_0303_),
    .Z(_0057_));
 INV_X1 _0844_ (.A(_0133_),
    .ZN(_0304_));
 NOR2_X1 _0845_ (.A1(_0137_),
    .A2(_0304_),
    .ZN(_0305_));
 AND2_X1 _0846_ (.A1(_0137_),
    .A2(_0304_),
    .ZN(_0306_));
 AOI21_X1 _0847_ (.A(_0305_),
    .B1(_0306_),
    .B2(_0303_),
    .ZN(_0307_));
 OAI22_X1 _0848_ (.A1(_0304_),
    .A2(_0303_),
    .B1(_0307_),
    .B2(_0297_),
    .ZN(_0058_));
 XNOR2_X1 _0849_ (.A(\rfifo.wp[0] ),
    .B(_0285_),
    .ZN(_0308_));
 NOR2_X1 _0850_ (.A1(_0297_),
    .A2(_0308_),
    .ZN(_0059_));
 NAND2_X1 _0851_ (.A1(_0285_),
    .A2(_0577_),
    .ZN(_0309_));
 INV_X1 _0852_ (.A(_0285_),
    .ZN(_0310_));
 NAND2_X1 _0853_ (.A1(_0310_),
    .A2(\rfifo.wp[1] ),
    .ZN(_0311_));
 AOI21_X1 _0854_ (.A(_0297_),
    .B1(_0309_),
    .B2(_0311_),
    .ZN(_0060_));
 NAND3_X4 _0855_ (.A1(net15),
    .A2(net6),
    .A3(net16),
    .ZN(_0312_));
 NOR3_X4 _0856_ (.A1(_0130_),
    .A2(_0139_),
    .A3(_0312_),
    .ZN(_0313_));
 MUX2_X1 _0857_ (.A(\espr[0] ),
    .B(net7),
    .S(_0313_),
    .Z(_0063_));
 MUX2_X1 _0858_ (.A(_0156_),
    .B(net8),
    .S(_0313_),
    .Z(_0064_));
 MUX2_X1 _0859_ (.A(cpha),
    .B(net9),
    .S(_0313_),
    .Z(_0065_));
 MUX2_X1 _0860_ (.A(cpol),
    .B(net10),
    .S(_0313_),
    .Z(_0066_));
 MUX2_X1 _0861_ (.A(dwom),
    .B(net12),
    .S(_0313_),
    .Z(_0067_));
 CLKBUF_X3 _0862_ (.A(_0186_),
    .Z(_0314_));
 CLKBUF_X2 _0863_ (.A(dat_i[6]),
    .Z(_0315_));
 MUX2_X1 _0864_ (.A(_0314_),
    .B(_0315_),
    .S(_0313_),
    .Z(_0068_));
 CLKBUF_X2 _0865_ (.A(dat_i[7]),
    .Z(_0316_));
 MUX2_X1 _0866_ (.A(spie),
    .B(_0316_),
    .S(_0313_),
    .Z(_0069_));
 NOR3_X4 _0867_ (.A1(_0131_),
    .A2(_0157_),
    .A3(_0312_),
    .ZN(_0317_));
 MUX2_X1 _0868_ (.A(_0144_),
    .B(net7),
    .S(_0317_),
    .Z(_0070_));
 MUX2_X1 _0869_ (.A(_0150_),
    .B(net8),
    .S(_0317_),
    .Z(_0071_));
 MUX2_X1 _0870_ (.A(\sper[2] ),
    .B(net9),
    .S(_0317_),
    .Z(_0072_));
 MUX2_X1 _0871_ (.A(\sper[3] ),
    .B(net10),
    .S(_0317_),
    .Z(_0073_));
 MUX2_X1 _0872_ (.A(\sper[4] ),
    .B(net11),
    .S(_0317_),
    .Z(_0074_));
 MUX2_X1 _0873_ (.A(\sper[5] ),
    .B(net12),
    .S(_0317_),
    .Z(_0075_));
 MUX2_X1 _0874_ (.A(\icnt[0] ),
    .B(_0315_),
    .S(_0317_),
    .Z(_0076_));
 MUX2_X1 _0875_ (.A(\icnt[1] ),
    .B(_0316_),
    .S(_0317_),
    .Z(_0077_));
 NOR2_X1 _0876_ (.A1(\tcnt[1] ),
    .A2(\tcnt[0] ),
    .ZN(_0318_));
 INV_X1 _0877_ (.A(_0318_),
    .ZN(_0319_));
 AOI21_X1 _0878_ (.A(\icnt[0] ),
    .B1(_0319_),
    .B2(_0314_),
    .ZN(_0320_));
 OR3_X1 _0879_ (.A1(_0310_),
    .A2(_0008_),
    .A3(_0318_),
    .ZN(_0321_));
 OAI21_X1 _0880_ (.A(_0321_),
    .B1(\tcnt[0] ),
    .B2(_0285_),
    .ZN(_0322_));
 BUF_X2 _0881_ (.A(_0186_),
    .Z(_0323_));
 AOI21_X1 _0882_ (.A(_0320_),
    .B1(_0322_),
    .B2(_0323_),
    .ZN(_0081_));
 NAND2_X1 _0883_ (.A1(_0285_),
    .A2(_0318_),
    .ZN(_0324_));
 NAND2_X1 _0884_ (.A1(_0314_),
    .A2(_0324_),
    .ZN(_0325_));
 NAND2_X1 _0885_ (.A1(\icnt[1] ),
    .A2(_0325_),
    .ZN(_0326_));
 NOR2_X1 _0886_ (.A1(_0310_),
    .A2(\tcnt[0] ),
    .ZN(_0327_));
 NAND2_X1 _0887_ (.A1(_0323_),
    .A2(\tcnt[1] ),
    .ZN(_0328_));
 OAI21_X1 _0888_ (.A(_0326_),
    .B1(_0327_),
    .B2(_0328_),
    .ZN(_0082_));
 NOR2_X4 _0889_ (.A1(_0300_),
    .A2(_0312_),
    .ZN(_0329_));
 NAND2_X4 _0890_ (.A1(_0586_),
    .A2(_0329_),
    .ZN(_0330_));
 MUX2_X1 _0891_ (.A(net7),
    .B(\wfifo.mem[0][0] ),
    .S(_0330_),
    .Z(_0093_));
 MUX2_X1 _0892_ (.A(net8),
    .B(\wfifo.mem[0][1] ),
    .S(_0330_),
    .Z(_0094_));
 MUX2_X1 _0893_ (.A(net9),
    .B(\wfifo.mem[0][2] ),
    .S(_0330_),
    .Z(_0095_));
 MUX2_X1 _0894_ (.A(net10),
    .B(\wfifo.mem[0][3] ),
    .S(_0330_),
    .Z(_0096_));
 MUX2_X1 _0895_ (.A(net11),
    .B(\wfifo.mem[0][4] ),
    .S(_0330_),
    .Z(_0097_));
 MUX2_X1 _0896_ (.A(net12),
    .B(\wfifo.mem[0][5] ),
    .S(_0330_),
    .Z(_0098_));
 MUX2_X1 _0897_ (.A(_0315_),
    .B(\wfifo.mem[0][6] ),
    .S(_0330_),
    .Z(_0099_));
 MUX2_X1 _0898_ (.A(_0316_),
    .B(\wfifo.mem[0][7] ),
    .S(_0330_),
    .Z(_0100_));
 NAND2_X4 _0899_ (.A1(_0590_),
    .A2(_0329_),
    .ZN(_0331_));
 MUX2_X1 _0900_ (.A(net7),
    .B(\wfifo.mem[1][0] ),
    .S(_0331_),
    .Z(_0101_));
 MUX2_X1 _0901_ (.A(net8),
    .B(\wfifo.mem[1][1] ),
    .S(_0331_),
    .Z(_0102_));
 MUX2_X1 _0902_ (.A(net9),
    .B(\wfifo.mem[1][2] ),
    .S(_0331_),
    .Z(_0103_));
 MUX2_X1 _0903_ (.A(net10),
    .B(\wfifo.mem[1][3] ),
    .S(_0331_),
    .Z(_0104_));
 MUX2_X1 _0904_ (.A(net11),
    .B(\wfifo.mem[1][4] ),
    .S(_0331_),
    .Z(_0105_));
 MUX2_X1 _0905_ (.A(net12),
    .B(\wfifo.mem[1][5] ),
    .S(_0331_),
    .Z(_0106_));
 MUX2_X1 _0906_ (.A(_0315_),
    .B(\wfifo.mem[1][6] ),
    .S(_0331_),
    .Z(_0107_));
 MUX2_X1 _0907_ (.A(_0316_),
    .B(\wfifo.mem[1][7] ),
    .S(_0331_),
    .Z(_0108_));
 NAND2_X4 _0908_ (.A1(_0588_),
    .A2(_0329_),
    .ZN(_0332_));
 MUX2_X1 _0909_ (.A(net7),
    .B(\wfifo.mem[2][0] ),
    .S(_0332_),
    .Z(_0109_));
 MUX2_X1 _0910_ (.A(net8),
    .B(\wfifo.mem[2][1] ),
    .S(_0332_),
    .Z(_0110_));
 MUX2_X1 _0911_ (.A(net9),
    .B(\wfifo.mem[2][2] ),
    .S(_0332_),
    .Z(_0111_));
 MUX2_X1 _0912_ (.A(net10),
    .B(\wfifo.mem[2][3] ),
    .S(_0332_),
    .Z(_0112_));
 MUX2_X1 _0913_ (.A(net11),
    .B(\wfifo.mem[2][4] ),
    .S(_0332_),
    .Z(_0113_));
 MUX2_X1 _0914_ (.A(net12),
    .B(\wfifo.mem[2][5] ),
    .S(_0332_),
    .Z(_0114_));
 MUX2_X1 _0915_ (.A(_0315_),
    .B(\wfifo.mem[2][6] ),
    .S(_0332_),
    .Z(_0115_));
 MUX2_X1 _0916_ (.A(_0316_),
    .B(\wfifo.mem[2][7] ),
    .S(_0332_),
    .Z(_0116_));
 NAND2_X4 _0917_ (.A1(_0592_),
    .A2(_0329_),
    .ZN(_0333_));
 MUX2_X1 _0918_ (.A(net7),
    .B(\wfifo.mem[3][0] ),
    .S(_0333_),
    .Z(_0117_));
 MUX2_X1 _0919_ (.A(net8),
    .B(\wfifo.mem[3][1] ),
    .S(_0333_),
    .Z(_0118_));
 MUX2_X1 _0920_ (.A(net9),
    .B(\wfifo.mem[3][2] ),
    .S(_0333_),
    .Z(_0119_));
 MUX2_X1 _0921_ (.A(net10),
    .B(\wfifo.mem[3][3] ),
    .S(_0333_),
    .Z(_0120_));
 MUX2_X1 _0922_ (.A(net11),
    .B(\wfifo.mem[3][4] ),
    .S(_0333_),
    .Z(_0121_));
 MUX2_X1 _0923_ (.A(net12),
    .B(\wfifo.mem[3][5] ),
    .S(_0333_),
    .Z(_0122_));
 MUX2_X1 _0924_ (.A(_0315_),
    .B(\wfifo.mem[3][6] ),
    .S(_0333_),
    .Z(_0123_));
 MUX2_X1 _0925_ (.A(_0316_),
    .B(\wfifo.mem[3][7] ),
    .S(_0333_),
    .Z(_0124_));
 CLKBUF_X3 _0926_ (.A(\wfifo.rp[0] ),
    .Z(_0334_));
 XNOR2_X1 _0927_ (.A(_0334_),
    .B(\wfifo.re ),
    .ZN(_0335_));
 NOR2_X1 _0928_ (.A1(_0297_),
    .A2(_0335_),
    .ZN(_0125_));
 CLKBUF_X3 _0929_ (.A(_0164_),
    .Z(_0336_));
 NAND2_X1 _0930_ (.A1(_0334_),
    .A2(\wfifo.re ),
    .ZN(_0337_));
 XOR2_X1 _0931_ (.A(_0336_),
    .B(_0337_),
    .Z(_0338_));
 NOR2_X1 _0932_ (.A1(_0297_),
    .A2(_0338_),
    .ZN(_0126_));
 NOR2_X1 _0933_ (.A1(\wfifo.wp[0] ),
    .A2(_0297_),
    .ZN(_0339_));
 NOR2_X1 _0934_ (.A1(_0005_),
    .A2(_0329_),
    .ZN(_0340_));
 MUX2_X1 _0935_ (.A(_0339_),
    .B(\wfifo.wp[0] ),
    .S(_0340_),
    .Z(_0127_));
 AND2_X1 _0936_ (.A1(_0186_),
    .A2(_0587_),
    .ZN(_0341_));
 MUX2_X1 _0937_ (.A(_0341_),
    .B(\wfifo.wp[1] ),
    .S(_0340_),
    .Z(_0128_));
 CLKBUF_X3 _0938_ (.A(_0600_),
    .Z(_0342_));
 CLKBUF_X3 _0939_ (.A(_0342_),
    .Z(_0343_));
 AND4_X1 _0940_ (.A1(_0343_),
    .A2(_0314_),
    .A3(_0613_),
    .A4(_0251_),
    .ZN(_0061_));
 OR2_X1 _0941_ (.A1(_0342_),
    .A2(_0197_),
    .ZN(_0344_));
 OAI21_X1 _0942_ (.A(_0314_),
    .B1(\bcnt[0] ),
    .B2(_0344_),
    .ZN(_0345_));
 XNOR2_X1 _0943_ (.A(\bcnt[0] ),
    .B(_0251_),
    .ZN(_0346_));
 AOI21_X1 _0944_ (.A(_0345_),
    .B1(_0346_),
    .B2(_0343_),
    .ZN(_0009_));
 OAI21_X1 _0945_ (.A(_0314_),
    .B1(\bcnt[1] ),
    .B2(_0344_),
    .ZN(_0347_));
 NOR3_X1 _0946_ (.A1(_0611_),
    .A2(_0206_),
    .A3(_0201_),
    .ZN(_0348_));
 NAND2_X1 _0947_ (.A1(_0217_),
    .A2(_0226_),
    .ZN(_0349_));
 AOI21_X1 _0948_ (.A(_0348_),
    .B1(_0349_),
    .B2(\bcnt[1] ),
    .ZN(_0350_));
 AOI21_X1 _0949_ (.A(_0347_),
    .B1(_0350_),
    .B2(_0343_),
    .ZN(_0010_));
 OAI21_X1 _0950_ (.A(_0314_),
    .B1(\bcnt[2] ),
    .B2(_0344_),
    .ZN(_0351_));
 NOR3_X1 _0951_ (.A1(_0614_),
    .A2(_0206_),
    .A3(_0201_),
    .ZN(_0352_));
 AOI21_X1 _0952_ (.A(_0352_),
    .B1(_0349_),
    .B2(\bcnt[2] ),
    .ZN(_0353_));
 AOI21_X1 _0953_ (.A(_0351_),
    .B1(_0353_),
    .B2(_0343_),
    .ZN(_0011_));
 NAND2_X1 _0954_ (.A1(_0314_),
    .A2(net14),
    .ZN(_0354_));
 XOR2_X1 _0955_ (.A(_0003_),
    .B(_0577_),
    .Z(_0355_));
 NAND3_X1 _0956_ (.A1(_0285_),
    .A2(_0147_),
    .A3(_0355_),
    .ZN(_0356_));
 OAI21_X1 _0957_ (.A(\rfifo.gb ),
    .B1(_0300_),
    .B2(_0302_),
    .ZN(_0357_));
 AOI21_X1 _0958_ (.A(_0354_),
    .B1(_0356_),
    .B2(_0357_),
    .ZN(_0024_));
 INV_X1 _0959_ (.A(net28),
    .ZN(_0358_));
 MUX2_X1 _0960_ (.A(_0007_),
    .B(cpol),
    .S(_0613_),
    .Z(_0359_));
 AOI22_X1 _0961_ (.A1(_0598_),
    .A2(_0358_),
    .B1(_0359_),
    .B2(_0342_),
    .ZN(_0360_));
 INV_X1 _0962_ (.A(_0595_),
    .ZN(_0361_));
 NAND4_X1 _0963_ (.A1(_0199_),
    .A2(\state[0] ),
    .A3(_0604_),
    .A4(_0200_),
    .ZN(_0362_));
 OAI22_X2 _0964_ (.A1(_0361_),
    .A2(\state[0] ),
    .B1(_0206_),
    .B2(_0362_),
    .ZN(_0363_));
 MUX2_X1 _0965_ (.A(_0358_),
    .B(_0360_),
    .S(_0363_),
    .Z(_0364_));
 INV_X1 _0966_ (.A(cpol),
    .ZN(_0365_));
 INV_X1 _0967_ (.A(_0007_),
    .ZN(_0366_));
 INV_X1 _0968_ (.A(cpha),
    .ZN(_0367_));
 NOR2_X1 _0969_ (.A1(_0367_),
    .A2(_0166_),
    .ZN(_0368_));
 MUX2_X1 _0970_ (.A(_0365_),
    .B(_0366_),
    .S(_0368_),
    .Z(_0369_));
 NOR2_X1 _0971_ (.A1(_0342_),
    .A2(_0598_),
    .ZN(_0370_));
 NAND3_X1 _0972_ (.A1(_0314_),
    .A2(_0363_),
    .A3(_0370_),
    .ZN(_0371_));
 OAI22_X1 _0973_ (.A1(_0297_),
    .A2(_0364_),
    .B1(_0369_),
    .B2(_0371_),
    .ZN(_0062_));
 INV_X1 _0974_ (.A(spif),
    .ZN(_0372_));
 NOR3_X1 _0975_ (.A1(_0131_),
    .A2(_0139_),
    .A3(_0312_),
    .ZN(_0373_));
 AOI221_X1 _0976_ (.A(_0297_),
    .B1(_0372_),
    .B2(_0324_),
    .C1(_0373_),
    .C2(_0316_),
    .ZN(_0078_));
 AOI21_X1 _0977_ (.A(_0370_),
    .B1(_0226_),
    .B2(_0217_),
    .ZN(_0374_));
 NAND4_X2 _0978_ (.A1(_0002_),
    .A2(_0197_),
    .A3(_0163_),
    .A4(_0165_),
    .ZN(_0375_));
 INV_X1 _0979_ (.A(_0197_),
    .ZN(_0376_));
 INV_X1 _0980_ (.A(_0613_),
    .ZN(_0377_));
 NAND3_X1 _0981_ (.A1(_0342_),
    .A2(_0377_),
    .A3(\state[1] ),
    .ZN(_0378_));
 AOI21_X1 _0982_ (.A(_0296_),
    .B1(_0376_),
    .B2(_0378_),
    .ZN(_0379_));
 NAND2_X1 _0983_ (.A1(_0375_),
    .A2(_0379_),
    .ZN(_0380_));
 NAND2_X1 _0984_ (.A1(_0314_),
    .A2(\state[0] ),
    .ZN(_0381_));
 NAND2_X1 _0985_ (.A1(\state[1] ),
    .A2(_0375_),
    .ZN(_0382_));
 NOR2_X1 _0986_ (.A1(_0374_),
    .A2(_0382_),
    .ZN(_0383_));
 OAI22_X1 _0987_ (.A1(_0374_),
    .A2(_0380_),
    .B1(_0381_),
    .B2(_0383_),
    .ZN(_0079_));
 AOI21_X1 _0988_ (.A(\state[1] ),
    .B1(_0251_),
    .B2(_0375_),
    .ZN(_0384_));
 AOI221_X2 _0989_ (.A(_0598_),
    .B1(_0166_),
    .B2(_0197_),
    .C1(_0349_),
    .C2(_0342_),
    .ZN(_0385_));
 NOR3_X1 _0990_ (.A1(_0297_),
    .A2(_0384_),
    .A3(_0385_),
    .ZN(_0080_));
 BUF_X2 _0991_ (.A(_0342_),
    .Z(_0386_));
 NAND2_X1 _0992_ (.A1(_0386_),
    .A2(net13),
    .ZN(_0387_));
 MUX2_X1 _0993_ (.A(\wfifo.mem[0][0] ),
    .B(\wfifo.mem[2][0] ),
    .S(_0336_),
    .Z(_0388_));
 MUX2_X1 _0994_ (.A(\wfifo.mem[1][0] ),
    .B(\wfifo.mem[3][0] ),
    .S(_0336_),
    .Z(_0389_));
 MUX2_X1 _0995_ (.A(_0388_),
    .B(_0389_),
    .S(_0334_),
    .Z(_0390_));
 INV_X1 _0996_ (.A(_0390_),
    .ZN(_0391_));
 AND3_X2 _0997_ (.A1(_0342_),
    .A2(_0217_),
    .A3(_0226_),
    .ZN(_0392_));
 BUF_X4 _0998_ (.A(_0392_),
    .Z(_0393_));
 NOR2_X2 _0999_ (.A1(_0342_),
    .A2(_0376_),
    .ZN(_0394_));
 BUF_X2 _1000_ (.A(_0394_),
    .Z(_0395_));
 OAI221_X1 _1001_ (.A(_0387_),
    .B1(_0391_),
    .B2(_0343_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0396_));
 OR3_X1 _1002_ (.A1(_0284_),
    .A2(_0393_),
    .A3(_0395_),
    .ZN(_0397_));
 AND3_X1 _1003_ (.A1(_0323_),
    .A2(_0396_),
    .A3(_0397_),
    .ZN(_0083_));
 NAND2_X1 _1004_ (.A1(_0386_),
    .A2(_0284_),
    .ZN(_0398_));
 MUX2_X1 _1005_ (.A(\wfifo.mem[0][1] ),
    .B(\wfifo.mem[2][1] ),
    .S(_0164_),
    .Z(_0399_));
 MUX2_X1 _1006_ (.A(\wfifo.mem[1][1] ),
    .B(\wfifo.mem[3][1] ),
    .S(_0336_),
    .Z(_0400_));
 MUX2_X1 _1007_ (.A(_0399_),
    .B(_0400_),
    .S(_0334_),
    .Z(_0401_));
 INV_X1 _1008_ (.A(_0401_),
    .ZN(_0402_));
 OAI221_X1 _1009_ (.A(_0398_),
    .B1(_0402_),
    .B2(_0343_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0403_));
 OR3_X1 _1010_ (.A1(_0287_),
    .A2(_0393_),
    .A3(_0395_),
    .ZN(_0404_));
 AND3_X1 _1011_ (.A1(_0323_),
    .A2(_0403_),
    .A3(_0404_),
    .ZN(_0084_));
 NAND2_X1 _1012_ (.A1(_0386_),
    .A2(_0287_),
    .ZN(_0405_));
 MUX2_X1 _1013_ (.A(\wfifo.mem[0][2] ),
    .B(\wfifo.mem[2][2] ),
    .S(_0164_),
    .Z(_0406_));
 MUX2_X1 _1014_ (.A(\wfifo.mem[1][2] ),
    .B(\wfifo.mem[3][2] ),
    .S(_0336_),
    .Z(_0407_));
 MUX2_X1 _1015_ (.A(_0406_),
    .B(_0407_),
    .S(_0334_),
    .Z(_0408_));
 INV_X1 _1016_ (.A(_0408_),
    .ZN(_0409_));
 OAI221_X1 _1017_ (.A(_0405_),
    .B1(_0409_),
    .B2(_0343_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0410_));
 OR3_X1 _1018_ (.A1(_0288_),
    .A2(_0392_),
    .A3(_0394_),
    .ZN(_0411_));
 AND3_X1 _1019_ (.A1(_0323_),
    .A2(_0410_),
    .A3(_0411_),
    .ZN(_0085_));
 NAND2_X1 _1020_ (.A1(_0386_),
    .A2(_0288_),
    .ZN(_0412_));
 MUX2_X1 _1021_ (.A(\wfifo.mem[0][3] ),
    .B(\wfifo.mem[2][3] ),
    .S(_0164_),
    .Z(_0413_));
 MUX2_X1 _1022_ (.A(\wfifo.mem[1][3] ),
    .B(\wfifo.mem[3][3] ),
    .S(_0336_),
    .Z(_0414_));
 MUX2_X1 _1023_ (.A(_0413_),
    .B(_0414_),
    .S(_0334_),
    .Z(_0415_));
 INV_X1 _1024_ (.A(_0415_),
    .ZN(_0416_));
 OAI221_X1 _1025_ (.A(_0412_),
    .B1(_0416_),
    .B2(_0343_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0417_));
 OR3_X1 _1026_ (.A1(_0289_),
    .A2(_0392_),
    .A3(_0394_),
    .ZN(_0418_));
 AND3_X1 _1027_ (.A1(_0323_),
    .A2(_0417_),
    .A3(_0418_),
    .ZN(_0086_));
 NAND2_X1 _1028_ (.A1(_0386_),
    .A2(_0289_),
    .ZN(_0419_));
 MUX2_X1 _1029_ (.A(\wfifo.mem[0][4] ),
    .B(\wfifo.mem[2][4] ),
    .S(_0164_),
    .Z(_0420_));
 MUX2_X1 _1030_ (.A(\wfifo.mem[1][4] ),
    .B(\wfifo.mem[3][4] ),
    .S(_0336_),
    .Z(_0421_));
 MUX2_X1 _1031_ (.A(_0420_),
    .B(_0421_),
    .S(_0334_),
    .Z(_0422_));
 INV_X1 _1032_ (.A(_0422_),
    .ZN(_0423_));
 OAI221_X1 _1033_ (.A(_0419_),
    .B1(_0423_),
    .B2(_0343_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0424_));
 OR3_X1 _1034_ (.A1(_0290_),
    .A2(_0392_),
    .A3(_0394_),
    .ZN(_0425_));
 AND3_X1 _1035_ (.A1(_0323_),
    .A2(_0424_),
    .A3(_0425_),
    .ZN(_0087_));
 NAND2_X1 _1036_ (.A1(_0386_),
    .A2(_0290_),
    .ZN(_0426_));
 MUX2_X1 _1037_ (.A(\wfifo.mem[0][5] ),
    .B(\wfifo.mem[2][5] ),
    .S(_0164_),
    .Z(_0427_));
 MUX2_X1 _1038_ (.A(\wfifo.mem[1][5] ),
    .B(\wfifo.mem[3][5] ),
    .S(_0336_),
    .Z(_0428_));
 MUX2_X1 _1039_ (.A(_0427_),
    .B(_0428_),
    .S(_0334_),
    .Z(_0429_));
 INV_X1 _1040_ (.A(_0429_),
    .ZN(_0430_));
 OAI221_X1 _1041_ (.A(_0426_),
    .B1(_0430_),
    .B2(_0343_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0431_));
 OR3_X1 _1042_ (.A1(_0291_),
    .A2(_0392_),
    .A3(_0394_),
    .ZN(_0432_));
 AND3_X1 _1043_ (.A1(_0323_),
    .A2(_0431_),
    .A3(_0432_),
    .ZN(_0088_));
 NAND2_X1 _1044_ (.A1(_0386_),
    .A2(_0291_),
    .ZN(_0433_));
 MUX2_X1 _1045_ (.A(\wfifo.mem[0][6] ),
    .B(\wfifo.mem[2][6] ),
    .S(_0164_),
    .Z(_0434_));
 MUX2_X1 _1046_ (.A(\wfifo.mem[1][6] ),
    .B(\wfifo.mem[3][6] ),
    .S(_0336_),
    .Z(_0435_));
 MUX2_X1 _1047_ (.A(_0434_),
    .B(_0435_),
    .S(_0334_),
    .Z(_0436_));
 INV_X1 _1048_ (.A(_0436_),
    .ZN(_0437_));
 OAI221_X1 _1049_ (.A(_0433_),
    .B1(_0437_),
    .B2(_0386_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0438_));
 OR3_X1 _1050_ (.A1(_0292_),
    .A2(_0392_),
    .A3(_0394_),
    .ZN(_0439_));
 AND3_X1 _1051_ (.A1(_0323_),
    .A2(_0438_),
    .A3(_0439_),
    .ZN(_0089_));
 NAND2_X1 _1052_ (.A1(_0386_),
    .A2(_0292_),
    .ZN(_0440_));
 MUX2_X1 _1053_ (.A(\wfifo.mem[0][7] ),
    .B(\wfifo.mem[2][7] ),
    .S(_0164_),
    .Z(_0441_));
 MUX2_X1 _1054_ (.A(\wfifo.mem[1][7] ),
    .B(\wfifo.mem[3][7] ),
    .S(_0336_),
    .Z(_0442_));
 MUX2_X1 _1055_ (.A(_0441_),
    .B(_0442_),
    .S(_0334_),
    .Z(_0443_));
 INV_X1 _1056_ (.A(_0443_),
    .ZN(_0444_));
 OAI221_X1 _1057_ (.A(_0440_),
    .B1(_0444_),
    .B2(_0386_),
    .C1(_0393_),
    .C2(_0395_),
    .ZN(_0445_));
 OR3_X1 _1058_ (.A1(net27),
    .A2(_0392_),
    .A3(_0394_),
    .ZN(_0446_));
 AND3_X1 _1059_ (.A1(_0323_),
    .A2(_0445_),
    .A3(_0446_),
    .ZN(_0090_));
 NAND2_X1 _1060_ (.A1(_0173_),
    .A2(_0329_),
    .ZN(_0447_));
 INV_X1 _1061_ (.A(wcol),
    .ZN(_0448_));
 AOI221_X1 _1062_ (.A(_0296_),
    .B1(_0315_),
    .B2(_0373_),
    .C1(_0447_),
    .C2(_0448_),
    .ZN(_0091_));
 INV_X1 _1063_ (.A(\wfifo.re ),
    .ZN(_0449_));
 XNOR2_X1 _1064_ (.A(_0006_),
    .B(_0587_),
    .ZN(_0450_));
 NOR2_X1 _1065_ (.A1(_0163_),
    .A2(_0450_),
    .ZN(_0451_));
 AOI22_X1 _1066_ (.A1(_0449_),
    .A2(\wfifo.gb ),
    .B1(_0329_),
    .B2(_0451_),
    .ZN(_0452_));
 NOR2_X1 _1067_ (.A1(_0354_),
    .A2(_0452_),
    .ZN(_0092_));
 NOR3_X1 _1068_ (.A1(_0005_),
    .A2(_0376_),
    .A3(_0166_),
    .ZN(_0129_));
 HA_X1 _1069_ (.A(_0574_),
    .B(_0575_),
    .CO(_0576_),
    .S(_0577_));
 HA_X1 _1070_ (.A(_0574_),
    .B(\rfifo.wp[1] ),
    .CO(_0578_),
    .S(_0579_));
 HA_X1 _1071_ (.A(\rfifo.wp[0] ),
    .B(_0575_),
    .CO(_0580_),
    .S(_0581_));
 HA_X1 _1072_ (.A(\rfifo.wp[0] ),
    .B(\rfifo.wp[1] ),
    .CO(_0582_),
    .S(_0583_));
 HA_X1 _1073_ (.A(_0584_),
    .B(_0585_),
    .CO(_0586_),
    .S(_0587_));
 HA_X1 _1074_ (.A(_0584_),
    .B(\wfifo.wp[1] ),
    .CO(_0588_),
    .S(_0589_));
 HA_X1 _1075_ (.A(\wfifo.wp[0] ),
    .B(_0585_),
    .CO(_0590_),
    .S(_0591_));
 HA_X1 _1076_ (.A(\wfifo.wp[0] ),
    .B(\wfifo.wp[1] ),
    .CO(_0592_),
    .S(_0593_));
 HA_X1 _1077_ (.A(_0594_),
    .B(_0595_),
    .CO(_0596_),
    .S(_0597_));
 HA_X1 _1078_ (.A(\state[0] ),
    .B(_0595_),
    .CO(_0598_),
    .S(_0599_));
 HA_X1 _1079_ (.A(\state[0] ),
    .B(\state[1] ),
    .CO(_0600_),
    .S(_0601_));
 HA_X1 _1080_ (.A(_0602_),
    .B(_0603_),
    .CO(_0604_),
    .S(_0605_));
 HA_X1 _1081_ (.A(_0602_),
    .B(_0603_),
    .CO(_0606_),
    .S(_0607_));
 HA_X1 _1082_ (.A(_0608_),
    .B(_0609_),
    .CO(_0610_),
    .S(_0611_));
 HA_X1 _1083_ (.A(_0612_),
    .B(_0610_),
    .CO(_0613_),
    .S(_0614_));
 DFFR_X1 \ack_o$_DFF_PN0_  (.D(_0000_),
    .RN(net3),
    .CK(clknet_4_9_0_clk_i),
    .Q(net17),
    .QN(_0004_));
 DFF_X1 \bcnt[0]$_SDFFE_PN0P_  (.D(_0009_),
    .CK(clknet_4_9_0_clk_i),
    .Q(\bcnt[0] ),
    .QN(_0608_));
 DFF_X1 \bcnt[1]$_SDFFE_PN0P_  (.D(_0010_),
    .CK(clknet_4_9_0_clk_i),
    .Q(\bcnt[1] ),
    .QN(_0609_));
 DFF_X1 \bcnt[2]$_SDFFE_PN0P_  (.D(_0011_),
    .CK(clknet_4_9_0_clk_i),
    .Q(\bcnt[2] ),
    .QN(_0612_));
 DFF_X2 \clkcnt[0]$_DFFE_PP_  (.D(_0012_),
    .CK(clknet_4_10_0_clk_i),
    .Q(\clkcnt[0] ),
    .QN(_0602_));
 DFF_X2 \clkcnt[10]$_DFFE_PP_  (.D(_0013_),
    .CK(clknet_4_11_0_clk_i),
    .Q(\clkcnt[10] ),
    .QN(_0564_));
 DFF_X1 \clkcnt[11]$_SDFFCE_PP0P_  (.D(_0014_),
    .CK(clknet_4_8_0_clk_i),
    .Q(\clkcnt[11] ),
    .QN(_0563_));
 DFF_X1 \clkcnt[1]$_DFFE_PP_  (.D(_0015_),
    .CK(clknet_4_8_0_clk_i),
    .Q(\clkcnt[1] ),
    .QN(_0603_));
 DFF_X1 \clkcnt[2]$_DFFE_PP_  (.D(_0016_),
    .CK(clknet_4_10_0_clk_i),
    .Q(\clkcnt[2] ),
    .QN(_0562_));
 DFF_X2 \clkcnt[3]$_DFFE_PP_  (.D(_0017_),
    .CK(clknet_4_10_0_clk_i),
    .Q(\clkcnt[3] ),
    .QN(_0561_));
 DFF_X1 \clkcnt[4]$_DFFE_PP_  (.D(_0018_),
    .CK(clknet_4_10_0_clk_i),
    .Q(\clkcnt[4] ),
    .QN(_0560_));
 DFF_X1 \clkcnt[5]$_DFFE_PP_  (.D(_0019_),
    .CK(clknet_4_10_0_clk_i),
    .Q(\clkcnt[5] ),
    .QN(_0559_));
 DFF_X2 \clkcnt[6]$_DFFE_PP_  (.D(_0020_),
    .CK(clknet_4_10_0_clk_i),
    .Q(\clkcnt[6] ),
    .QN(_0558_));
 DFF_X1 \clkcnt[7]$_DFFE_PP_  (.D(_0021_),
    .CK(clknet_4_11_0_clk_i),
    .Q(\clkcnt[7] ),
    .QN(_0557_));
 DFF_X2 \clkcnt[8]$_DFFE_PP_  (.D(_0022_),
    .CK(clknet_4_11_0_clk_i),
    .Q(\clkcnt[8] ),
    .QN(_0556_));
 DFF_X2 \clkcnt[9]$_DFFE_PP_  (.D(_0023_),
    .CK(clknet_4_11_0_clk_i),
    .Q(\clkcnt[9] ),
    .QN(_0565_));
 DFF_X1 \dat_o[0]$_DFF_P_  (.D(_0453_),
    .CK(clknet_4_9_0_clk_i),
    .Q(net18),
    .QN(_0566_));
 DFF_X1 \dat_o[1]$_DFF_P_  (.D(_0454_),
    .CK(clknet_4_11_0_clk_i),
    .Q(net19),
    .QN(_0567_));
 DFF_X1 \dat_o[2]$_DFF_P_  (.D(_0455_),
    .CK(clknet_4_5_0_clk_i),
    .Q(net20),
    .QN(_0568_));
 DFF_X1 \dat_o[3]$_DFF_P_  (.D(_0456_),
    .CK(clknet_4_5_0_clk_i),
    .Q(net21),
    .QN(_0569_));
 DFF_X1 \dat_o[4]$_DFF_P_  (.D(_0457_),
    .CK(clknet_4_5_0_clk_i),
    .Q(net22),
    .QN(_0570_));
 DFF_X1 \dat_o[5]$_DFF_P_  (.D(_0458_),
    .CK(clknet_4_5_0_clk_i),
    .Q(net23),
    .QN(_0571_));
 DFF_X1 \dat_o[6]$_DFF_P_  (.D(_0459_),
    .CK(clknet_4_15_0_clk_i),
    .Q(net24),
    .QN(_0572_));
 DFF_X1 \dat_o[7]$_DFF_P_  (.D(_0460_),
    .CK(clknet_4_5_0_clk_i),
    .Q(net25),
    .QN(_0573_));
 DFF_X1 \inta_o$_DFF_P_  (.D(_0001_),
    .CK(clknet_4_5_0_clk_i),
    .Q(net26),
    .QN(_0555_));
 DFF_X1 \rfifo.gb$_SDFFE_PN0P_  (.D(_0024_),
    .CK(clknet_4_12_0_clk_i),
    .Q(\rfifo.gb ),
    .QN(_0554_));
 DFF_X1 \rfifo.mem[0][0]$_DFFE_PP_  (.D(_0025_),
    .CK(clknet_4_13_0_clk_i),
    .Q(\rfifo.mem[0][0] ),
    .QN(_0553_));
 DFF_X1 \rfifo.mem[0][1]$_DFFE_PP_  (.D(_0026_),
    .CK(clknet_4_14_0_clk_i),
    .Q(\rfifo.mem[0][1] ),
    .QN(_0552_));
 DFF_X1 \rfifo.mem[0][2]$_DFFE_PP_  (.D(_0027_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.mem[0][2] ),
    .QN(_0551_));
 DFF_X1 \rfifo.mem[0][3]$_DFFE_PP_  (.D(_0028_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[0][3] ),
    .QN(_0550_));
 DFF_X1 \rfifo.mem[0][4]$_DFFE_PP_  (.D(_0029_),
    .CK(clknet_4_15_0_clk_i),
    .Q(\rfifo.mem[0][4] ),
    .QN(_0549_));
 DFF_X1 \rfifo.mem[0][5]$_DFFE_PP_  (.D(_0030_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.mem[0][5] ),
    .QN(_0548_));
 DFF_X1 \rfifo.mem[0][6]$_DFFE_PP_  (.D(_0031_),
    .CK(clknet_4_15_0_clk_i),
    .Q(\rfifo.mem[0][6] ),
    .QN(_0547_));
 DFF_X1 \rfifo.mem[0][7]$_DFFE_PP_  (.D(_0032_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[0][7] ),
    .QN(_0546_));
 DFF_X1 \rfifo.mem[1][0]$_DFFE_PP_  (.D(_0033_),
    .CK(clknet_4_14_0_clk_i),
    .Q(\rfifo.mem[1][0] ),
    .QN(_0545_));
 DFF_X1 \rfifo.mem[1][1]$_DFFE_PP_  (.D(_0034_),
    .CK(clknet_4_15_0_clk_i),
    .Q(\rfifo.mem[1][1] ),
    .QN(_0544_));
 DFF_X1 \rfifo.mem[1][2]$_DFFE_PP_  (.D(_0035_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.mem[1][2] ),
    .QN(_0543_));
 DFF_X1 \rfifo.mem[1][3]$_DFFE_PP_  (.D(_0036_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[1][3] ),
    .QN(_0542_));
 DFF_X1 \rfifo.mem[1][4]$_DFFE_PP_  (.D(_0037_),
    .CK(clknet_4_15_0_clk_i),
    .Q(\rfifo.mem[1][4] ),
    .QN(_0541_));
 DFF_X1 \rfifo.mem[1][5]$_DFFE_PP_  (.D(_0038_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[1][5] ),
    .QN(_0540_));
 DFF_X1 \rfifo.mem[1][6]$_DFFE_PP_  (.D(_0039_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[1][6] ),
    .QN(_0539_));
 DFF_X1 \rfifo.mem[1][7]$_DFFE_PP_  (.D(_0040_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[1][7] ),
    .QN(_0538_));
 DFF_X1 \rfifo.mem[2][0]$_DFFE_PP_  (.D(_0041_),
    .CK(clknet_4_14_0_clk_i),
    .Q(\rfifo.mem[2][0] ),
    .QN(_0537_));
 DFF_X1 \rfifo.mem[2][1]$_DFFE_PP_  (.D(_0042_),
    .CK(clknet_4_14_0_clk_i),
    .Q(\rfifo.mem[2][1] ),
    .QN(_0536_));
 DFF_X1 \rfifo.mem[2][2]$_DFFE_PP_  (.D(_0043_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.mem[2][2] ),
    .QN(_0535_));
 DFF_X1 \rfifo.mem[2][3]$_DFFE_PP_  (.D(_0044_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[2][3] ),
    .QN(_0534_));
 DFF_X1 \rfifo.mem[2][4]$_DFFE_PP_  (.D(_0045_),
    .CK(clknet_4_15_0_clk_i),
    .Q(\rfifo.mem[2][4] ),
    .QN(_0533_));
 DFF_X1 \rfifo.mem[2][5]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.mem[2][5] ),
    .QN(_0532_));
 DFF_X1 \rfifo.mem[2][6]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[2][6] ),
    .QN(_0531_));
 DFF_X1 \rfifo.mem[2][7]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[2][7] ),
    .QN(_0530_));
 DFF_X1 \rfifo.mem[3][0]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_4_14_0_clk_i),
    .Q(\rfifo.mem[3][0] ),
    .QN(_0529_));
 DFF_X1 \rfifo.mem[3][1]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_4_14_0_clk_i),
    .Q(\rfifo.mem[3][1] ),
    .QN(_0528_));
 DFF_X1 \rfifo.mem[3][2]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.mem[3][2] ),
    .QN(_0527_));
 DFF_X1 \rfifo.mem[3][3]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[3][3] ),
    .QN(_0526_));
 DFF_X1 \rfifo.mem[3][4]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_4_15_0_clk_i),
    .Q(\rfifo.mem[3][4] ),
    .QN(_0525_));
 DFF_X1 \rfifo.mem[3][5]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[3][5] ),
    .QN(_0524_));
 DFF_X1 \rfifo.mem[3][6]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[3][6] ),
    .QN(_0523_));
 DFF_X1 \rfifo.mem[3][7]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_4_7_0_clk_i),
    .Q(\rfifo.mem[3][7] ),
    .QN(_0522_));
 DFFR_X1 \rfifo.rp[0]$_DFFE_PN0P_  (.D(_0057_),
    .RN(net3),
    .CK(clknet_4_13_0_clk_i),
    .Q(\rfifo.rp[0] ),
    .QN(_0521_));
 DFFR_X1 \rfifo.rp[1]$_DFFE_PN0P_  (.D(_0058_),
    .RN(net3),
    .CK(clknet_4_13_0_clk_i),
    .Q(\rfifo.rp[1] ),
    .QN(_0003_));
 DFFR_X2 \rfifo.wp[0]$_DFFE_PN0P_  (.D(_0059_),
    .RN(net3),
    .CK(clknet_4_13_0_clk_i),
    .Q(\rfifo.wp[0] ),
    .QN(_0574_));
 DFFR_X2 \rfifo.wp[1]$_DFFE_PN0P_  (.D(_0060_),
    .RN(net3),
    .CK(clknet_4_13_0_clk_i),
    .Q(\rfifo.wp[1] ),
    .QN(_0575_));
 DFF_X1 \rfwe$_SDFF_PP0_  (.D(_0061_),
    .CK(clknet_4_12_0_clk_i),
    .Q(\rfifo.we ),
    .QN(_0520_));
 DFF_X1 \sck_o$_SDFFE_PN0P_  (.D(_0062_),
    .CK(clknet_4_12_0_clk_i),
    .Q(net28),
    .QN(_0007_));
 DFFR_X1 \spcr[0]$_DFFE_PN0P_  (.D(_0063_),
    .RN(net3),
    .CK(clknet_4_8_0_clk_i),
    .Q(\espr[0] ),
    .QN(_0519_));
 DFFR_X1 \spcr[1]$_DFFE_PN0P_  (.D(_0064_),
    .RN(net3),
    .CK(clknet_4_8_0_clk_i),
    .Q(\espr[1] ),
    .QN(_0518_));
 DFFR_X1 \spcr[2]$_DFFE_PN0P_  (.D(_0065_),
    .RN(net3),
    .CK(clknet_4_4_0_clk_i),
    .Q(cpha),
    .QN(_0517_));
 DFFR_X1 \spcr[3]$_DFFE_PN0P_  (.D(_0066_),
    .RN(net3),
    .CK(clknet_4_3_0_clk_i),
    .Q(cpol),
    .QN(_0516_));
 DFFR_X1 \spcr[5]$_DFFE_PN0P_  (.D(_0067_),
    .RN(net3),
    .CK(clknet_4_4_0_clk_i),
    .Q(dwom),
    .QN(_0515_));
 DFFR_X2 \spcr[6]$_DFFE_PN0P_  (.D(_0068_),
    .RN(net3),
    .CK(clknet_4_3_0_clk_i),
    .Q(spe),
    .QN(_0005_));
 DFFR_X1 \spcr[7]$_DFFE_PN0P_  (.D(_0069_),
    .RN(net3),
    .CK(clknet_4_5_0_clk_i),
    .Q(spie),
    .QN(_0514_));
 DFFR_X1 \sper[0]$_DFFE_PN0P_  (.D(_0070_),
    .RN(net3),
    .CK(clknet_4_8_0_clk_i),
    .Q(\espr[2] ),
    .QN(_0513_));
 DFFR_X1 \sper[1]$_DFFE_PN0P_  (.D(_0071_),
    .RN(net3),
    .CK(clknet_4_8_0_clk_i),
    .Q(\espr[3] ),
    .QN(_0512_));
 DFFR_X1 \sper[2]$_DFFE_PN0P_  (.D(_0072_),
    .RN(net3),
    .CK(clknet_4_1_0_clk_i),
    .Q(\sper[2] ),
    .QN(_0511_));
 DFFR_X1 \sper[3]$_DFFE_PN0P_  (.D(_0073_),
    .RN(net3),
    .CK(clknet_4_1_0_clk_i),
    .Q(\sper[3] ),
    .QN(_0510_));
 DFFR_X1 \sper[4]$_DFFE_PN0P_  (.D(_0074_),
    .RN(net3),
    .CK(clknet_4_5_0_clk_i),
    .Q(\sper[4] ),
    .QN(_0509_));
 DFFR_X1 \sper[5]$_DFFE_PN0P_  (.D(_0075_),
    .RN(net3),
    .CK(clknet_4_5_0_clk_i),
    .Q(\sper[5] ),
    .QN(_0508_));
 DFFR_X1 \sper[6]$_DFFE_PN0P_  (.D(_0076_),
    .RN(net3),
    .CK(clknet_4_12_0_clk_i),
    .Q(\icnt[0] ),
    .QN(_0507_));
 DFFR_X1 \sper[7]$_DFFE_PN0P_  (.D(_0077_),
    .RN(net3),
    .CK(clknet_4_4_0_clk_i),
    .Q(\icnt[1] ),
    .QN(_0506_));
 DFF_X1 \spif$_SDFF_PN0_  (.D(_0078_),
    .CK(clknet_4_12_0_clk_i),
    .Q(spif),
    .QN(_0505_));
 DFF_X2 \state[0]$_SDFFE_PN0P_  (.D(_0079_),
    .CK(clknet_4_9_0_clk_i),
    .Q(\state[0] ),
    .QN(_0594_));
 DFF_X2 \state[1]$_SDFFE_PN0P_  (.D(_0080_),
    .CK(clknet_4_8_0_clk_i),
    .Q(\state[1] ),
    .QN(_0595_));
 DFF_X1 \tcnt[0]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_4_13_0_clk_i),
    .Q(\tcnt[0] ),
    .QN(_0008_));
 DFF_X1 \tcnt[1]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_4_13_0_clk_i),
    .Q(\tcnt[1] ),
    .QN(_0504_));
 DFF_X1 \treg[0]$_SDFFE_PN0P_  (.D(_0083_),
    .CK(clknet_4_12_0_clk_i),
    .Q(\rfifo.din[1] ),
    .QN(_0503_));
 DFF_X1 \treg[1]$_SDFFE_PN0P_  (.D(_0084_),
    .CK(clknet_4_4_0_clk_i),
    .Q(\rfifo.din[2] ),
    .QN(_0502_));
 DFF_X1 \treg[2]$_SDFFE_PN0P_  (.D(_0085_),
    .CK(clknet_4_4_0_clk_i),
    .Q(\rfifo.din[3] ),
    .QN(_0501_));
 DFF_X1 \treg[3]$_SDFFE_PN0P_  (.D(_0086_),
    .CK(clknet_4_4_0_clk_i),
    .Q(\rfifo.din[4] ),
    .QN(_0500_));
 DFF_X1 \treg[4]$_SDFFE_PN0P_  (.D(_0087_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.din[5] ),
    .QN(_0499_));
 DFF_X1 \treg[5]$_SDFFE_PN0P_  (.D(_0088_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.din[6] ),
    .QN(_0498_));
 DFF_X1 \treg[6]$_SDFFE_PN0P_  (.D(_0089_),
    .CK(clknet_4_6_0_clk_i),
    .Q(\rfifo.din[7] ),
    .QN(_0497_));
 DFF_X2 \treg[7]$_SDFFE_PN0P_  (.D(_0090_),
    .CK(clknet_4_4_0_clk_i),
    .Q(net27),
    .QN(_0496_));
 DFF_X1 \wcol$_SDFF_PN0_  (.D(_0091_),
    .CK(clknet_4_12_0_clk_i),
    .Q(wcol),
    .QN(_0495_));
 DFF_X1 \wfifo.gb$_SDFFE_PN0P_  (.D(_0092_),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.gb ),
    .QN(_0002_));
 DFF_X1 \wfifo.mem[0][0]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[0][0] ),
    .QN(_0494_));
 DFF_X1 \wfifo.mem[0][1]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[0][1] ),
    .QN(_0493_));
 DFF_X1 \wfifo.mem[0][2]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[0][2] ),
    .QN(_0492_));
 DFF_X1 \wfifo.mem[0][3]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[0][3] ),
    .QN(_0491_));
 DFF_X1 \wfifo.mem[0][4]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[0][4] ),
    .QN(_0490_));
 DFF_X1 \wfifo.mem[0][5]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[0][5] ),
    .QN(_0489_));
 DFF_X1 \wfifo.mem[0][6]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.mem[0][6] ),
    .QN(_0488_));
 DFF_X1 \wfifo.mem[0][7]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[0][7] ),
    .QN(_0487_));
 DFF_X1 \wfifo.mem[1][0]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[1][0] ),
    .QN(_0486_));
 DFF_X1 \wfifo.mem[1][1]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[1][1] ),
    .QN(_0485_));
 DFF_X1 \wfifo.mem[1][2]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[1][2] ),
    .QN(_0484_));
 DFF_X1 \wfifo.mem[1][3]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[1][3] ),
    .QN(_0483_));
 DFF_X1 \wfifo.mem[1][4]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[1][4] ),
    .QN(_0482_));
 DFF_X1 \wfifo.mem[1][5]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[1][5] ),
    .QN(_0481_));
 DFF_X1 \wfifo.mem[1][6]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.mem[1][6] ),
    .QN(_0480_));
 DFF_X1 \wfifo.mem[1][7]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[1][7] ),
    .QN(_0479_));
 DFF_X1 \wfifo.mem[2][0]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[2][0] ),
    .QN(_0478_));
 DFF_X1 \wfifo.mem[2][1]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[2][1] ),
    .QN(_0477_));
 DFF_X1 \wfifo.mem[2][2]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[2][2] ),
    .QN(_0476_));
 DFF_X1 \wfifo.mem[2][3]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[2][3] ),
    .QN(_0475_));
 DFF_X1 \wfifo.mem[2][4]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[2][4] ),
    .QN(_0474_));
 DFF_X1 \wfifo.mem[2][5]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[2][5] ),
    .QN(_0473_));
 DFF_X1 \wfifo.mem[2][6]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.mem[2][6] ),
    .QN(_0472_));
 DFF_X1 \wfifo.mem[2][7]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[2][7] ),
    .QN(_0471_));
 DFF_X1 \wfifo.mem[3][0]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[3][0] ),
    .QN(_0470_));
 DFF_X1 \wfifo.mem[3][1]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.mem[3][1] ),
    .QN(_0469_));
 DFF_X1 \wfifo.mem[3][2]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[3][2] ),
    .QN(_0468_));
 DFF_X1 \wfifo.mem[3][3]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[3][3] ),
    .QN(_0467_));
 DFF_X1 \wfifo.mem[3][4]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_4_0_0_clk_i),
    .Q(\wfifo.mem[3][4] ),
    .QN(_0466_));
 DFF_X1 \wfifo.mem[3][5]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[3][5] ),
    .QN(_0465_));
 DFF_X1 \wfifo.mem[3][6]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.mem[3][6] ),
    .QN(_0464_));
 DFF_X1 \wfifo.mem[3][7]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_4_1_0_clk_i),
    .Q(\wfifo.mem[3][7] ),
    .QN(_0463_));
 DFFR_X1 \wfifo.rp[0]$_DFFE_PN0P_  (.D(_0125_),
    .RN(net3),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.rp[0] ),
    .QN(_0462_));
 DFFR_X1 \wfifo.rp[1]$_DFFE_PN0P_  (.D(_0126_),
    .RN(net3),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.rp[1] ),
    .QN(_0006_));
 DFFR_X2 \wfifo.wp[0]$_DFFE_PN0P_  (.D(_0127_),
    .RN(net3),
    .CK(clknet_4_8_0_clk_i),
    .Q(\wfifo.wp[0] ),
    .QN(_0584_));
 DFFR_X2 \wfifo.wp[1]$_DFFE_PN0P_  (.D(_0128_),
    .RN(net3),
    .CK(clknet_4_2_0_clk_i),
    .Q(\wfifo.wp[1] ),
    .QN(_0585_));
 DFF_X1 \wfre$_SDFF_PN0_  (.D(_0129_),
    .CK(clknet_4_3_0_clk_i),
    .Q(\wfifo.re ),
    .QN(_0461_));
 CLKBUF_X1 hold1 (.A(net5),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(net4),
    .Z(net2));
 BUF_X8 hold3 (.A(net1),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(net30),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(net2),
    .Z(net5));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_77 ();
 CLKBUF_X2 input1 (.A(cyc_i),
    .Z(net6));
 BUF_X1 input2 (.A(dat_i[0]),
    .Z(net7));
 BUF_X1 input3 (.A(dat_i[1]),
    .Z(net8));
 BUF_X1 input4 (.A(dat_i[2]),
    .Z(net9));
 BUF_X1 input5 (.A(dat_i[3]),
    .Z(net10));
 BUF_X1 input6 (.A(dat_i[4]),
    .Z(net11));
 BUF_X1 input7 (.A(dat_i[5]),
    .Z(net12));
 BUF_X1 input8 (.A(miso_i),
    .Z(net13));
 BUF_X1 input9 (.A(net29),
    .Z(net14));
 CLKBUF_X2 input10 (.A(stb_i),
    .Z(net15));
 CLKBUF_X2 input11 (.A(we_i),
    .Z(net16));
 BUF_X1 output12 (.A(net17),
    .Z(ack_o));
 BUF_X1 output13 (.A(net18),
    .Z(dat_o[0]));
 BUF_X1 output14 (.A(net19),
    .Z(dat_o[1]));
 BUF_X1 output15 (.A(net20),
    .Z(dat_o[2]));
 BUF_X1 output16 (.A(net21),
    .Z(dat_o[3]));
 BUF_X1 output17 (.A(net22),
    .Z(dat_o[4]));
 BUF_X1 output18 (.A(net23),
    .Z(dat_o[5]));
 BUF_X1 output19 (.A(net24),
    .Z(dat_o[6]));
 BUF_X1 output20 (.A(net25),
    .Z(dat_o[7]));
 BUF_X1 output21 (.A(net26),
    .Z(inta_o));
 BUF_X1 output22 (.A(net27),
    .Z(mosi_o));
 BUF_X1 output23 (.A(net28),
    .Z(sck_o));
 CLKBUF_X3 clkbuf_0_clk_i (.A(clk_i),
    .Z(clknet_0_clk_i));
 CLKBUF_X3 clkbuf_4_0_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_0_0_clk_i));
 CLKBUF_X3 clkbuf_4_1_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_1_0_clk_i));
 CLKBUF_X3 clkbuf_4_2_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_2_0_clk_i));
 CLKBUF_X3 clkbuf_4_3_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_3_0_clk_i));
 CLKBUF_X3 clkbuf_4_4_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_4_0_clk_i));
 CLKBUF_X3 clkbuf_4_5_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_5_0_clk_i));
 CLKBUF_X3 clkbuf_4_6_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_6_0_clk_i));
 CLKBUF_X3 clkbuf_4_7_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_7_0_clk_i));
 CLKBUF_X3 clkbuf_4_8_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_8_0_clk_i));
 CLKBUF_X3 clkbuf_4_9_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_9_0_clk_i));
 CLKBUF_X3 clkbuf_4_10_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_10_0_clk_i));
 CLKBUF_X3 clkbuf_4_11_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_11_0_clk_i));
 CLKBUF_X3 clkbuf_4_12_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_12_0_clk_i));
 CLKBUF_X3 clkbuf_4_13_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_13_0_clk_i));
 CLKBUF_X3 clkbuf_4_14_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_14_0_clk_i));
 CLKBUF_X3 clkbuf_4_15_0_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_4_15_0_clk_i));
 INV_X2 clkload0 (.A(clknet_4_0_0_clk_i));
 CLKBUF_X1 clkload1 (.A(clknet_4_1_0_clk_i));
 CLKBUF_X1 clkload2 (.A(clknet_4_2_0_clk_i));
 INV_X2 clkload3 (.A(clknet_4_3_0_clk_i));
 INV_X4 clkload4 (.A(clknet_4_4_0_clk_i));
 INV_X2 clkload5 (.A(clknet_4_5_0_clk_i));
 INV_X2 clkload6 (.A(clknet_4_6_0_clk_i));
 INV_X2 clkload7 (.A(clknet_4_8_0_clk_i));
 INV_X4 clkload8 (.A(clknet_4_9_0_clk_i));
 INV_X4 clkload9 (.A(clknet_4_10_0_clk_i));
 INV_X4 clkload10 (.A(clknet_4_11_0_clk_i));
 INV_X4 clkload11 (.A(clknet_4_12_0_clk_i));
 INV_X4 clkload12 (.A(clknet_4_13_0_clk_i));
 INV_X4 clkload13 (.A(clknet_4_14_0_clk_i));
 INV_X4 clkload14 (.A(clknet_4_15_0_clk_i));
 CLKBUF_X1 hold6 (.A(rst_i),
    .Z(net29));
 CLKBUF_X1 hold7 (.A(net14),
    .Z(net30));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X4 FILLER_0_57 ();
 FILLCELL_X1 FILLER_0_61 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_73 ();
 FILLCELL_X2 FILLER_0_77 ();
 FILLCELL_X1 FILLER_0_79 ();
 FILLCELL_X2 FILLER_0_97 ();
 FILLCELL_X1 FILLER_0_99 ();
 FILLCELL_X16 FILLER_0_103 ();
 FILLCELL_X8 FILLER_0_119 ();
 FILLCELL_X4 FILLER_0_127 ();
 FILLCELL_X2 FILLER_0_131 ();
 FILLCELL_X1 FILLER_0_133 ();
 FILLCELL_X8 FILLER_0_138 ();
 FILLCELL_X2 FILLER_0_146 ();
 FILLCELL_X1 FILLER_0_148 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X1 FILLER_0_174 ();
 FILLCELL_X1 FILLER_0_178 ();
 FILLCELL_X4 FILLER_0_182 ();
 FILLCELL_X2 FILLER_0_186 ();
 FILLCELL_X1 FILLER_0_188 ();
 FILLCELL_X32 FILLER_0_209 ();
 FILLCELL_X32 FILLER_0_241 ();
 FILLCELL_X16 FILLER_0_273 ();
 FILLCELL_X4 FILLER_0_289 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X16 FILLER_1_33 ();
 FILLCELL_X1 FILLER_1_49 ();
 FILLCELL_X8 FILLER_1_74 ();
 FILLCELL_X1 FILLER_1_82 ();
 FILLCELL_X1 FILLER_1_97 ();
 FILLCELL_X16 FILLER_1_105 ();
 FILLCELL_X2 FILLER_1_121 ();
 FILLCELL_X1 FILLER_1_123 ();
 FILLCELL_X8 FILLER_1_144 ();
 FILLCELL_X4 FILLER_1_152 ();
 FILLCELL_X2 FILLER_1_156 ();
 FILLCELL_X1 FILLER_1_158 ();
 FILLCELL_X4 FILLER_1_179 ();
 FILLCELL_X2 FILLER_1_183 ();
 FILLCELL_X4 FILLER_1_190 ();
 FILLCELL_X2 FILLER_1_194 ();
 FILLCELL_X1 FILLER_1_196 ();
 FILLCELL_X32 FILLER_1_200 ();
 FILLCELL_X32 FILLER_1_232 ();
 FILLCELL_X16 FILLER_1_264 ();
 FILLCELL_X8 FILLER_1_280 ();
 FILLCELL_X4 FILLER_1_288 ();
 FILLCELL_X1 FILLER_1_292 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_57 ();
 FILLCELL_X4 FILLER_2_76 ();
 FILLCELL_X2 FILLER_2_80 ();
 FILLCELL_X1 FILLER_2_99 ();
 FILLCELL_X4 FILLER_2_117 ();
 FILLCELL_X2 FILLER_2_121 ();
 FILLCELL_X1 FILLER_2_123 ();
 FILLCELL_X8 FILLER_2_144 ();
 FILLCELL_X4 FILLER_2_169 ();
 FILLCELL_X4 FILLER_2_180 ();
 FILLCELL_X1 FILLER_2_184 ();
 FILLCELL_X32 FILLER_2_202 ();
 FILLCELL_X32 FILLER_2_234 ();
 FILLCELL_X16 FILLER_2_266 ();
 FILLCELL_X8 FILLER_2_282 ();
 FILLCELL_X2 FILLER_2_290 ();
 FILLCELL_X1 FILLER_2_292 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_49 ();
 FILLCELL_X4 FILLER_3_57 ();
 FILLCELL_X8 FILLER_3_75 ();
 FILLCELL_X4 FILLER_3_83 ();
 FILLCELL_X8 FILLER_3_111 ();
 FILLCELL_X2 FILLER_3_119 ();
 FILLCELL_X4 FILLER_3_135 ();
 FILLCELL_X2 FILLER_3_139 ();
 FILLCELL_X1 FILLER_3_141 ();
 FILLCELL_X2 FILLER_3_150 ();
 FILLCELL_X1 FILLER_3_169 ();
 FILLCELL_X4 FILLER_3_177 ();
 FILLCELL_X32 FILLER_3_197 ();
 FILLCELL_X32 FILLER_3_229 ();
 FILLCELL_X32 FILLER_3_261 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_41 ();
 FILLCELL_X16 FILLER_4_62 ();
 FILLCELL_X8 FILLER_4_78 ();
 FILLCELL_X4 FILLER_4_86 ();
 FILLCELL_X8 FILLER_4_97 ();
 FILLCELL_X1 FILLER_4_105 ();
 FILLCELL_X16 FILLER_4_113 ();
 FILLCELL_X2 FILLER_4_129 ();
 FILLCELL_X1 FILLER_4_131 ();
 FILLCELL_X16 FILLER_4_139 ();
 FILLCELL_X8 FILLER_4_155 ();
 FILLCELL_X2 FILLER_4_163 ();
 FILLCELL_X1 FILLER_4_165 ();
 FILLCELL_X32 FILLER_4_200 ();
 FILLCELL_X32 FILLER_4_232 ();
 FILLCELL_X16 FILLER_4_264 ();
 FILLCELL_X8 FILLER_4_280 ();
 FILLCELL_X4 FILLER_4_288 ();
 FILLCELL_X1 FILLER_4_292 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_33 ();
 FILLCELL_X2 FILLER_5_41 ();
 FILLCELL_X1 FILLER_5_43 ();
 FILLCELL_X16 FILLER_5_58 ();
 FILLCELL_X32 FILLER_5_91 ();
 FILLCELL_X2 FILLER_5_130 ();
 FILLCELL_X1 FILLER_5_156 ();
 FILLCELL_X8 FILLER_5_199 ();
 FILLCELL_X4 FILLER_5_207 ();
 FILLCELL_X1 FILLER_5_211 ();
 FILLCELL_X32 FILLER_5_229 ();
 FILLCELL_X4 FILLER_5_261 ();
 FILLCELL_X8 FILLER_5_282 ();
 FILLCELL_X2 FILLER_5_290 ();
 FILLCELL_X1 FILLER_5_292 ();
 FILLCELL_X2 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_3 ();
 FILLCELL_X4 FILLER_6_21 ();
 FILLCELL_X2 FILLER_6_25 ();
 FILLCELL_X4 FILLER_6_44 ();
 FILLCELL_X2 FILLER_6_48 ();
 FILLCELL_X4 FILLER_6_67 ();
 FILLCELL_X1 FILLER_6_71 ();
 FILLCELL_X1 FILLER_6_79 ();
 FILLCELL_X1 FILLER_6_87 ();
 FILLCELL_X8 FILLER_6_100 ();
 FILLCELL_X2 FILLER_6_135 ();
 FILLCELL_X2 FILLER_6_144 ();
 FILLCELL_X1 FILLER_6_146 ();
 FILLCELL_X32 FILLER_6_164 ();
 FILLCELL_X8 FILLER_6_196 ();
 FILLCELL_X1 FILLER_6_204 ();
 FILLCELL_X4 FILLER_6_236 ();
 FILLCELL_X1 FILLER_6_240 ();
 FILLCELL_X4 FILLER_6_258 ();
 FILLCELL_X4 FILLER_6_269 ();
 FILLCELL_X2 FILLER_6_273 ();
 FILLCELL_X1 FILLER_6_275 ();
 FILLCELL_X8 FILLER_6_279 ();
 FILLCELL_X4 FILLER_6_287 ();
 FILLCELL_X2 FILLER_6_291 ();
 FILLCELL_X2 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_3 ();
 FILLCELL_X4 FILLER_7_11 ();
 FILLCELL_X1 FILLER_7_15 ();
 FILLCELL_X2 FILLER_7_33 ();
 FILLCELL_X1 FILLER_7_71 ();
 FILLCELL_X8 FILLER_7_113 ();
 FILLCELL_X2 FILLER_7_121 ();
 FILLCELL_X1 FILLER_7_123 ();
 FILLCELL_X4 FILLER_7_144 ();
 FILLCELL_X1 FILLER_7_148 ();
 FILLCELL_X1 FILLER_7_156 ();
 FILLCELL_X8 FILLER_7_176 ();
 FILLCELL_X4 FILLER_7_184 ();
 FILLCELL_X1 FILLER_7_188 ();
 FILLCELL_X16 FILLER_7_193 ();
 FILLCELL_X1 FILLER_7_250 ();
 FILLCELL_X2 FILLER_7_258 ();
 FILLCELL_X1 FILLER_7_267 ();
 FILLCELL_X1 FILLER_7_275 ();
 FILLCELL_X8 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_9 ();
 FILLCELL_X2 FILLER_8_13 ();
 FILLCELL_X2 FILLER_8_22 ();
 FILLCELL_X1 FILLER_8_24 ();
 FILLCELL_X8 FILLER_8_32 ();
 FILLCELL_X4 FILLER_8_40 ();
 FILLCELL_X2 FILLER_8_44 ();
 FILLCELL_X1 FILLER_8_46 ();
 FILLCELL_X4 FILLER_8_78 ();
 FILLCELL_X2 FILLER_8_82 ();
 FILLCELL_X1 FILLER_8_84 ();
 FILLCELL_X32 FILLER_8_112 ();
 FILLCELL_X16 FILLER_8_181 ();
 FILLCELL_X8 FILLER_8_197 ();
 FILLCELL_X4 FILLER_8_205 ();
 FILLCELL_X2 FILLER_8_240 ();
 FILLCELL_X8 FILLER_8_256 ();
 FILLCELL_X4 FILLER_8_264 ();
 FILLCELL_X16 FILLER_8_275 ();
 FILLCELL_X2 FILLER_8_291 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_33 ();
 FILLCELL_X2 FILLER_9_37 ();
 FILLCELL_X32 FILLER_9_44 ();
 FILLCELL_X4 FILLER_9_76 ();
 FILLCELL_X2 FILLER_9_80 ();
 FILLCELL_X4 FILLER_9_84 ();
 FILLCELL_X2 FILLER_9_88 ();
 FILLCELL_X1 FILLER_9_111 ();
 FILLCELL_X8 FILLER_9_114 ();
 FILLCELL_X1 FILLER_9_122 ();
 FILLCELL_X8 FILLER_9_125 ();
 FILLCELL_X2 FILLER_9_133 ();
 FILLCELL_X1 FILLER_9_135 ();
 FILLCELL_X4 FILLER_9_138 ();
 FILLCELL_X2 FILLER_9_142 ();
 FILLCELL_X1 FILLER_9_144 ();
 FILLCELL_X2 FILLER_9_176 ();
 FILLCELL_X16 FILLER_9_195 ();
 FILLCELL_X4 FILLER_9_211 ();
 FILLCELL_X8 FILLER_9_229 ();
 FILLCELL_X2 FILLER_9_237 ();
 FILLCELL_X1 FILLER_9_244 ();
 FILLCELL_X2 FILLER_9_264 ();
 FILLCELL_X1 FILLER_9_266 ();
 FILLCELL_X8 FILLER_9_281 ();
 FILLCELL_X4 FILLER_9_289 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_9 ();
 FILLCELL_X8 FILLER_10_27 ();
 FILLCELL_X4 FILLER_10_35 ();
 FILLCELL_X32 FILLER_10_56 ();
 FILLCELL_X8 FILLER_10_88 ();
 FILLCELL_X1 FILLER_10_96 ();
 FILLCELL_X8 FILLER_10_99 ();
 FILLCELL_X4 FILLER_10_107 ();
 FILLCELL_X2 FILLER_10_111 ();
 FILLCELL_X1 FILLER_10_113 ();
 FILLCELL_X2 FILLER_10_134 ();
 FILLCELL_X2 FILLER_10_173 ();
 FILLCELL_X1 FILLER_10_175 ();
 FILLCELL_X8 FILLER_10_186 ();
 FILLCELL_X1 FILLER_10_194 ();
 FILLCELL_X4 FILLER_10_198 ();
 FILLCELL_X16 FILLER_10_210 ();
 FILLCELL_X4 FILLER_10_226 ();
 FILLCELL_X1 FILLER_10_230 ();
 FILLCELL_X1 FILLER_10_248 ();
 FILLCELL_X4 FILLER_10_266 ();
 FILLCELL_X2 FILLER_10_270 ();
 FILLCELL_X1 FILLER_10_272 ();
 FILLCELL_X2 FILLER_10_290 ();
 FILLCELL_X1 FILLER_10_292 ();
 FILLCELL_X1 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_5 ();
 FILLCELL_X2 FILLER_11_9 ();
 FILLCELL_X2 FILLER_11_25 ();
 FILLCELL_X1 FILLER_11_27 ();
 FILLCELL_X1 FILLER_11_35 ();
 FILLCELL_X1 FILLER_11_67 ();
 FILLCELL_X8 FILLER_11_101 ();
 FILLCELL_X2 FILLER_11_109 ();
 FILLCELL_X16 FILLER_11_118 ();
 FILLCELL_X2 FILLER_11_141 ();
 FILLCELL_X8 FILLER_11_150 ();
 FILLCELL_X2 FILLER_11_158 ();
 FILLCELL_X32 FILLER_11_174 ();
 FILLCELL_X2 FILLER_11_223 ();
 FILLCELL_X1 FILLER_11_225 ();
 FILLCELL_X1 FILLER_11_233 ();
 FILLCELL_X4 FILLER_11_241 ();
 FILLCELL_X2 FILLER_11_245 ();
 FILLCELL_X1 FILLER_11_247 ();
 FILLCELL_X16 FILLER_11_262 ();
 FILLCELL_X8 FILLER_11_278 ();
 FILLCELL_X4 FILLER_11_286 ();
 FILLCELL_X2 FILLER_11_290 ();
 FILLCELL_X1 FILLER_11_292 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X2 FILLER_12_13 ();
 FILLCELL_X1 FILLER_12_15 ();
 FILLCELL_X8 FILLER_12_33 ();
 FILLCELL_X1 FILLER_12_41 ();
 FILLCELL_X1 FILLER_12_49 ();
 FILLCELL_X1 FILLER_12_57 ();
 FILLCELL_X1 FILLER_12_75 ();
 FILLCELL_X2 FILLER_12_83 ();
 FILLCELL_X1 FILLER_12_92 ();
 FILLCELL_X2 FILLER_12_107 ();
 FILLCELL_X2 FILLER_12_136 ();
 FILLCELL_X4 FILLER_12_140 ();
 FILLCELL_X2 FILLER_12_144 ();
 FILLCELL_X1 FILLER_12_146 ();
 FILLCELL_X4 FILLER_12_150 ();
 FILLCELL_X4 FILLER_12_158 ();
 FILLCELL_X2 FILLER_12_162 ();
 FILLCELL_X1 FILLER_12_164 ();
 FILLCELL_X2 FILLER_12_168 ();
 FILLCELL_X1 FILLER_12_197 ();
 FILLCELL_X2 FILLER_12_201 ();
 FILLCELL_X4 FILLER_12_224 ();
 FILLCELL_X2 FILLER_12_228 ();
 FILLCELL_X8 FILLER_12_247 ();
 FILLCELL_X16 FILLER_12_272 ();
 FILLCELL_X4 FILLER_12_288 ();
 FILLCELL_X1 FILLER_12_292 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X16 FILLER_13_20 ();
 FILLCELL_X8 FILLER_13_53 ();
 FILLCELL_X4 FILLER_13_61 ();
 FILLCELL_X2 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_67 ();
 FILLCELL_X32 FILLER_13_109 ();
 FILLCELL_X2 FILLER_13_141 ();
 FILLCELL_X1 FILLER_13_152 ();
 FILLCELL_X1 FILLER_13_158 ();
 FILLCELL_X16 FILLER_13_173 ();
 FILLCELL_X8 FILLER_13_189 ();
 FILLCELL_X2 FILLER_13_197 ();
 FILLCELL_X1 FILLER_13_199 ();
 FILLCELL_X4 FILLER_13_217 ();
 FILLCELL_X2 FILLER_13_221 ();
 FILLCELL_X16 FILLER_13_237 ();
 FILLCELL_X4 FILLER_13_253 ();
 FILLCELL_X2 FILLER_13_262 ();
 FILLCELL_X16 FILLER_13_271 ();
 FILLCELL_X4 FILLER_13_287 ();
 FILLCELL_X2 FILLER_13_291 ();
 FILLCELL_X2 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_3 ();
 FILLCELL_X4 FILLER_14_7 ();
 FILLCELL_X1 FILLER_14_11 ();
 FILLCELL_X2 FILLER_14_19 ();
 FILLCELL_X1 FILLER_14_21 ();
 FILLCELL_X2 FILLER_14_36 ();
 FILLCELL_X2 FILLER_14_45 ();
 FILLCELL_X1 FILLER_14_47 ();
 FILLCELL_X32 FILLER_14_62 ();
 FILLCELL_X1 FILLER_14_94 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X8 FILLER_14_129 ();
 FILLCELL_X1 FILLER_14_137 ();
 FILLCELL_X2 FILLER_14_160 ();
 FILLCELL_X1 FILLER_14_177 ();
 FILLCELL_X16 FILLER_14_198 ();
 FILLCELL_X8 FILLER_14_214 ();
 FILLCELL_X1 FILLER_14_222 ();
 FILLCELL_X8 FILLER_14_247 ();
 FILLCELL_X1 FILLER_14_272 ();
 FILLCELL_X2 FILLER_14_290 ();
 FILLCELL_X1 FILLER_14_292 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_9 ();
 FILLCELL_X2 FILLER_15_13 ();
 FILLCELL_X4 FILLER_15_32 ();
 FILLCELL_X1 FILLER_15_36 ();
 FILLCELL_X4 FILLER_15_61 ();
 FILLCELL_X2 FILLER_15_65 ();
 FILLCELL_X1 FILLER_15_67 ();
 FILLCELL_X4 FILLER_15_74 ();
 FILLCELL_X1 FILLER_15_78 ();
 FILLCELL_X8 FILLER_15_99 ();
 FILLCELL_X1 FILLER_15_107 ();
 FILLCELL_X4 FILLER_15_129 ();
 FILLCELL_X4 FILLER_15_142 ();
 FILLCELL_X2 FILLER_15_150 ();
 FILLCELL_X1 FILLER_15_152 ();
 FILLCELL_X4 FILLER_15_166 ();
 FILLCELL_X1 FILLER_15_170 ();
 FILLCELL_X4 FILLER_15_174 ();
 FILLCELL_X2 FILLER_15_178 ();
 FILLCELL_X1 FILLER_15_180 ();
 FILLCELL_X32 FILLER_15_200 ();
 FILLCELL_X8 FILLER_15_232 ();
 FILLCELL_X4 FILLER_15_240 ();
 FILLCELL_X8 FILLER_15_275 ();
 FILLCELL_X4 FILLER_15_283 ();
 FILLCELL_X2 FILLER_15_287 ();
 FILLCELL_X1 FILLER_15_289 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X1 FILLER_16_21 ();
 FILLCELL_X2 FILLER_16_56 ();
 FILLCELL_X1 FILLER_16_83 ();
 FILLCELL_X4 FILLER_16_103 ();
 FILLCELL_X2 FILLER_16_107 ();
 FILLCELL_X1 FILLER_16_109 ();
 FILLCELL_X4 FILLER_16_112 ();
 FILLCELL_X2 FILLER_16_143 ();
 FILLCELL_X8 FILLER_16_153 ();
 FILLCELL_X16 FILLER_16_187 ();
 FILLCELL_X8 FILLER_16_203 ();
 FILLCELL_X2 FILLER_16_211 ();
 FILLCELL_X1 FILLER_16_213 ();
 FILLCELL_X1 FILLER_16_219 ();
 FILLCELL_X4 FILLER_16_244 ();
 FILLCELL_X2 FILLER_16_265 ();
 FILLCELL_X2 FILLER_16_291 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X1 FILLER_17_25 ();
 FILLCELL_X2 FILLER_17_33 ();
 FILLCELL_X1 FILLER_17_35 ();
 FILLCELL_X16 FILLER_17_50 ();
 FILLCELL_X4 FILLER_17_66 ();
 FILLCELL_X4 FILLER_17_79 ();
 FILLCELL_X4 FILLER_17_89 ();
 FILLCELL_X4 FILLER_17_103 ();
 FILLCELL_X4 FILLER_17_122 ();
 FILLCELL_X2 FILLER_17_126 ();
 FILLCELL_X1 FILLER_17_130 ();
 FILLCELL_X1 FILLER_17_136 ();
 FILLCELL_X4 FILLER_17_178 ();
 FILLCELL_X2 FILLER_17_182 ();
 FILLCELL_X1 FILLER_17_184 ();
 FILLCELL_X8 FILLER_17_199 ();
 FILLCELL_X1 FILLER_17_207 ();
 FILLCELL_X1 FILLER_17_212 ();
 FILLCELL_X2 FILLER_17_222 ();
 FILLCELL_X1 FILLER_17_224 ();
 FILLCELL_X2 FILLER_17_250 ();
 FILLCELL_X16 FILLER_17_273 ();
 FILLCELL_X4 FILLER_17_289 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_9 ();
 FILLCELL_X2 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_30 ();
 FILLCELL_X16 FILLER_18_55 ();
 FILLCELL_X2 FILLER_18_71 ();
 FILLCELL_X1 FILLER_18_76 ();
 FILLCELL_X2 FILLER_18_91 ();
 FILLCELL_X1 FILLER_18_128 ();
 FILLCELL_X16 FILLER_18_132 ();
 FILLCELL_X8 FILLER_18_148 ();
 FILLCELL_X1 FILLER_18_181 ();
 FILLCELL_X1 FILLER_18_185 ();
 FILLCELL_X1 FILLER_18_189 ();
 FILLCELL_X1 FILLER_18_197 ();
 FILLCELL_X4 FILLER_18_209 ();
 FILLCELL_X2 FILLER_18_213 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X2 FILLER_18_257 ();
 FILLCELL_X4 FILLER_18_266 ();
 FILLCELL_X2 FILLER_18_270 ();
 FILLCELL_X8 FILLER_18_279 ();
 FILLCELL_X4 FILLER_18_287 ();
 FILLCELL_X2 FILLER_18_291 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X2 FILLER_19_13 ();
 FILLCELL_X1 FILLER_19_15 ();
 FILLCELL_X16 FILLER_19_47 ();
 FILLCELL_X4 FILLER_19_122 ();
 FILLCELL_X1 FILLER_19_132 ();
 FILLCELL_X4 FILLER_19_142 ();
 FILLCELL_X2 FILLER_19_146 ();
 FILLCELL_X16 FILLER_19_153 ();
 FILLCELL_X8 FILLER_19_169 ();
 FILLCELL_X1 FILLER_19_177 ();
 FILLCELL_X1 FILLER_19_210 ();
 FILLCELL_X16 FILLER_19_218 ();
 FILLCELL_X2 FILLER_19_234 ();
 FILLCELL_X1 FILLER_19_236 ();
 FILLCELL_X8 FILLER_19_246 ();
 FILLCELL_X2 FILLER_19_254 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X16 FILLER_20_33 ();
 FILLCELL_X4 FILLER_20_49 ();
 FILLCELL_X2 FILLER_20_53 ();
 FILLCELL_X16 FILLER_20_96 ();
 FILLCELL_X2 FILLER_20_112 ();
 FILLCELL_X1 FILLER_20_114 ();
 FILLCELL_X1 FILLER_20_124 ();
 FILLCELL_X1 FILLER_20_129 ();
 FILLCELL_X4 FILLER_20_132 ();
 FILLCELL_X2 FILLER_20_136 ();
 FILLCELL_X16 FILLER_20_143 ();
 FILLCELL_X8 FILLER_20_159 ();
 FILLCELL_X2 FILLER_20_167 ();
 FILLCELL_X1 FILLER_20_173 ();
 FILLCELL_X1 FILLER_20_204 ();
 FILLCELL_X2 FILLER_20_248 ();
 FILLCELL_X1 FILLER_20_250 ();
 FILLCELL_X8 FILLER_20_285 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X16 FILLER_21_33 ();
 FILLCELL_X8 FILLER_21_49 ();
 FILLCELL_X8 FILLER_21_86 ();
 FILLCELL_X4 FILLER_21_94 ();
 FILLCELL_X1 FILLER_21_105 ();
 FILLCELL_X1 FILLER_21_110 ();
 FILLCELL_X1 FILLER_21_121 ();
 FILLCELL_X16 FILLER_21_176 ();
 FILLCELL_X4 FILLER_21_192 ();
 FILLCELL_X4 FILLER_21_287 ();
 FILLCELL_X2 FILLER_21_291 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_65 ();
 FILLCELL_X4 FILLER_22_73 ();
 FILLCELL_X8 FILLER_22_84 ();
 FILLCELL_X2 FILLER_22_92 ();
 FILLCELL_X2 FILLER_22_122 ();
 FILLCELL_X1 FILLER_22_124 ();
 FILLCELL_X8 FILLER_22_141 ();
 FILLCELL_X4 FILLER_22_149 ();
 FILLCELL_X1 FILLER_22_153 ();
 FILLCELL_X4 FILLER_22_197 ();
 FILLCELL_X2 FILLER_22_201 ();
 FILLCELL_X1 FILLER_22_203 ();
 FILLCELL_X2 FILLER_22_208 ();
 FILLCELL_X1 FILLER_22_210 ();
 FILLCELL_X2 FILLER_22_227 ();
 FILLCELL_X4 FILLER_22_257 ();
 FILLCELL_X4 FILLER_22_278 ();
 FILLCELL_X8 FILLER_22_285 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X8 FILLER_23_80 ();
 FILLCELL_X4 FILLER_23_88 ();
 FILLCELL_X1 FILLER_23_121 ();
 FILLCELL_X2 FILLER_23_126 ();
 FILLCELL_X16 FILLER_23_141 ();
 FILLCELL_X2 FILLER_23_157 ();
 FILLCELL_X1 FILLER_23_159 ();
 FILLCELL_X2 FILLER_23_163 ();
 FILLCELL_X1 FILLER_23_165 ();
 FILLCELL_X32 FILLER_23_192 ();
 FILLCELL_X16 FILLER_23_224 ();
 FILLCELL_X1 FILLER_23_240 ();
 FILLCELL_X8 FILLER_23_260 ();
 FILLCELL_X2 FILLER_23_268 ();
 FILLCELL_X1 FILLER_23_270 ();
 FILLCELL_X8 FILLER_23_278 ();
 FILLCELL_X4 FILLER_23_286 ();
 FILLCELL_X2 FILLER_23_290 ();
 FILLCELL_X1 FILLER_23_292 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_33 ();
 FILLCELL_X8 FILLER_24_49 ();
 FILLCELL_X1 FILLER_24_57 ();
 FILLCELL_X4 FILLER_24_98 ();
 FILLCELL_X1 FILLER_24_102 ();
 FILLCELL_X2 FILLER_24_113 ();
 FILLCELL_X1 FILLER_24_115 ();
 FILLCELL_X1 FILLER_24_121 ();
 FILLCELL_X1 FILLER_24_127 ();
 FILLCELL_X2 FILLER_24_132 ();
 FILLCELL_X1 FILLER_24_134 ();
 FILLCELL_X16 FILLER_24_142 ();
 FILLCELL_X1 FILLER_24_158 ();
 FILLCELL_X4 FILLER_24_173 ();
 FILLCELL_X16 FILLER_24_194 ();
 FILLCELL_X8 FILLER_24_210 ();
 FILLCELL_X2 FILLER_24_218 ();
 FILLCELL_X2 FILLER_24_234 ();
 FILLCELL_X2 FILLER_24_270 ();
 FILLCELL_X1 FILLER_24_272 ();
 FILLCELL_X2 FILLER_24_290 ();
 FILLCELL_X1 FILLER_24_292 ();
 FILLCELL_X1 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_5 ();
 FILLCELL_X2 FILLER_25_9 ();
 FILLCELL_X32 FILLER_25_14 ();
 FILLCELL_X4 FILLER_25_46 ();
 FILLCELL_X2 FILLER_25_57 ();
 FILLCELL_X1 FILLER_25_59 ();
 FILLCELL_X4 FILLER_25_67 ();
 FILLCELL_X2 FILLER_25_71 ();
 FILLCELL_X2 FILLER_25_84 ();
 FILLCELL_X16 FILLER_25_90 ();
 FILLCELL_X8 FILLER_25_106 ();
 FILLCELL_X1 FILLER_25_123 ();
 FILLCELL_X1 FILLER_25_141 ();
 FILLCELL_X2 FILLER_25_156 ();
 FILLCELL_X1 FILLER_25_158 ();
 FILLCELL_X8 FILLER_25_194 ();
 FILLCELL_X4 FILLER_25_202 ();
 FILLCELL_X1 FILLER_25_213 ();
 FILLCELL_X4 FILLER_25_228 ();
 FILLCELL_X2 FILLER_25_239 ();
 FILLCELL_X1 FILLER_25_241 ();
 FILLCELL_X2 FILLER_25_263 ();
 FILLCELL_X1 FILLER_25_265 ();
 FILLCELL_X2 FILLER_25_290 ();
 FILLCELL_X1 FILLER_25_292 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X16 FILLER_26_33 ();
 FILLCELL_X4 FILLER_26_49 ();
 FILLCELL_X1 FILLER_26_53 ();
 FILLCELL_X8 FILLER_26_99 ();
 FILLCELL_X2 FILLER_26_107 ();
 FILLCELL_X1 FILLER_26_109 ();
 FILLCELL_X1 FILLER_26_137 ();
 FILLCELL_X1 FILLER_26_142 ();
 FILLCELL_X2 FILLER_26_157 ();
 FILLCELL_X4 FILLER_26_169 ();
 FILLCELL_X2 FILLER_26_176 ();
 FILLCELL_X1 FILLER_26_178 ();
 FILLCELL_X8 FILLER_26_187 ();
 FILLCELL_X4 FILLER_26_195 ();
 FILLCELL_X8 FILLER_26_250 ();
 FILLCELL_X2 FILLER_26_258 ();
 FILLCELL_X16 FILLER_26_274 ();
 FILLCELL_X2 FILLER_26_290 ();
 FILLCELL_X1 FILLER_26_292 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X4 FILLER_27_81 ();
 FILLCELL_X2 FILLER_27_85 ();
 FILLCELL_X4 FILLER_27_90 ();
 FILLCELL_X8 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_105 ();
 FILLCELL_X2 FILLER_27_109 ();
 FILLCELL_X1 FILLER_27_111 ();
 FILLCELL_X2 FILLER_27_135 ();
 FILLCELL_X1 FILLER_27_145 ();
 FILLCELL_X8 FILLER_27_163 ();
 FILLCELL_X2 FILLER_27_171 ();
 FILLCELL_X1 FILLER_27_173 ();
 FILLCELL_X16 FILLER_27_194 ();
 FILLCELL_X2 FILLER_27_210 ();
 FILLCELL_X32 FILLER_27_236 ();
 FILLCELL_X16 FILLER_27_268 ();
 FILLCELL_X8 FILLER_27_284 ();
 FILLCELL_X1 FILLER_27_292 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X16 FILLER_28_65 ();
 FILLCELL_X8 FILLER_28_81 ();
 FILLCELL_X4 FILLER_28_89 ();
 FILLCELL_X1 FILLER_28_93 ();
 FILLCELL_X8 FILLER_28_120 ();
 FILLCELL_X4 FILLER_28_128 ();
 FILLCELL_X2 FILLER_28_136 ();
 FILLCELL_X1 FILLER_28_138 ();
 FILLCELL_X8 FILLER_28_143 ();
 FILLCELL_X4 FILLER_28_151 ();
 FILLCELL_X2 FILLER_28_155 ();
 FILLCELL_X4 FILLER_28_170 ();
 FILLCELL_X1 FILLER_28_179 ();
 FILLCELL_X32 FILLER_28_197 ();
 FILLCELL_X32 FILLER_28_229 ();
 FILLCELL_X32 FILLER_28_261 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X16 FILLER_29_33 ();
 FILLCELL_X4 FILLER_29_49 ();
 FILLCELL_X1 FILLER_29_53 ();
 FILLCELL_X1 FILLER_29_116 ();
 FILLCELL_X4 FILLER_29_120 ();
 FILLCELL_X1 FILLER_29_124 ();
 FILLCELL_X16 FILLER_29_139 ();
 FILLCELL_X4 FILLER_29_155 ();
 FILLCELL_X2 FILLER_29_159 ();
 FILLCELL_X4 FILLER_29_163 ();
 FILLCELL_X4 FILLER_29_171 ();
 FILLCELL_X1 FILLER_29_175 ();
 FILLCELL_X4 FILLER_29_179 ();
 FILLCELL_X1 FILLER_29_183 ();
 FILLCELL_X1 FILLER_29_190 ();
 FILLCELL_X32 FILLER_29_207 ();
 FILLCELL_X32 FILLER_29_239 ();
 FILLCELL_X16 FILLER_29_271 ();
 FILLCELL_X4 FILLER_29_287 ();
 FILLCELL_X2 FILLER_29_291 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X16 FILLER_30_33 ();
 FILLCELL_X8 FILLER_30_49 ();
 FILLCELL_X1 FILLER_30_57 ();
 FILLCELL_X2 FILLER_30_85 ();
 FILLCELL_X1 FILLER_30_87 ();
 FILLCELL_X4 FILLER_30_92 ();
 FILLCELL_X1 FILLER_30_96 ();
 FILLCELL_X2 FILLER_30_102 ();
 FILLCELL_X1 FILLER_30_109 ();
 FILLCELL_X16 FILLER_30_147 ();
 FILLCELL_X8 FILLER_30_163 ();
 FILLCELL_X4 FILLER_30_171 ();
 FILLCELL_X1 FILLER_30_175 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X4 FILLER_30_289 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X4 FILLER_31_65 ();
 FILLCELL_X1 FILLER_31_104 ();
 FILLCELL_X2 FILLER_31_109 ();
 FILLCELL_X32 FILLER_31_169 ();
 FILLCELL_X32 FILLER_31_201 ();
 FILLCELL_X32 FILLER_31_233 ();
 FILLCELL_X16 FILLER_31_265 ();
 FILLCELL_X8 FILLER_31_281 ();
 FILLCELL_X4 FILLER_31_289 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X16 FILLER_32_33 ();
 FILLCELL_X8 FILLER_32_49 ();
 FILLCELL_X2 FILLER_32_92 ();
 FILLCELL_X2 FILLER_32_97 ();
 FILLCELL_X2 FILLER_32_105 ();
 FILLCELL_X1 FILLER_32_107 ();
 FILLCELL_X32 FILLER_32_172 ();
 FILLCELL_X32 FILLER_32_204 ();
 FILLCELL_X32 FILLER_32_236 ();
 FILLCELL_X16 FILLER_32_268 ();
 FILLCELL_X8 FILLER_32_284 ();
 FILLCELL_X1 FILLER_32_292 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X2 FILLER_33_65 ();
 FILLCELL_X1 FILLER_33_67 ();
 FILLCELL_X1 FILLER_33_71 ();
 FILLCELL_X1 FILLER_33_75 ();
 FILLCELL_X2 FILLER_33_82 ();
 FILLCELL_X4 FILLER_33_93 ();
 FILLCELL_X2 FILLER_33_97 ();
 FILLCELL_X1 FILLER_33_99 ();
 FILLCELL_X8 FILLER_33_114 ();
 FILLCELL_X1 FILLER_33_122 ();
 FILLCELL_X4 FILLER_33_126 ();
 FILLCELL_X2 FILLER_33_130 ();
 FILLCELL_X32 FILLER_33_151 ();
 FILLCELL_X32 FILLER_33_183 ();
 FILLCELL_X32 FILLER_33_215 ();
 FILLCELL_X32 FILLER_33_247 ();
 FILLCELL_X8 FILLER_33_279 ();
 FILLCELL_X4 FILLER_33_287 ();
 FILLCELL_X2 FILLER_33_291 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X2 FILLER_34_65 ();
 FILLCELL_X1 FILLER_34_67 ();
 FILLCELL_X2 FILLER_34_87 ();
 FILLCELL_X4 FILLER_34_94 ();
 FILLCELL_X2 FILLER_34_98 ();
 FILLCELL_X1 FILLER_34_100 ();
 FILLCELL_X2 FILLER_34_108 ();
 FILLCELL_X32 FILLER_34_132 ();
 FILLCELL_X4 FILLER_34_164 ();
 FILLCELL_X32 FILLER_34_171 ();
 FILLCELL_X32 FILLER_34_203 ();
 FILLCELL_X32 FILLER_34_235 ();
 FILLCELL_X16 FILLER_34_267 ();
 FILLCELL_X8 FILLER_34_283 ();
 FILLCELL_X2 FILLER_34_291 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X1 FILLER_35_65 ();
 FILLCELL_X1 FILLER_35_70 ();
 FILLCELL_X1 FILLER_35_77 ();
 FILLCELL_X1 FILLER_35_103 ();
 FILLCELL_X1 FILLER_35_121 ();
 FILLCELL_X4 FILLER_35_126 ();
 FILLCELL_X2 FILLER_35_130 ();
 FILLCELL_X32 FILLER_35_144 ();
 FILLCELL_X32 FILLER_35_176 ();
 FILLCELL_X32 FILLER_35_208 ();
 FILLCELL_X32 FILLER_35_240 ();
 FILLCELL_X16 FILLER_35_272 ();
 FILLCELL_X4 FILLER_35_288 ();
 FILLCELL_X1 FILLER_35_292 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X16 FILLER_36_33 ();
 FILLCELL_X8 FILLER_36_49 ();
 FILLCELL_X4 FILLER_36_57 ();
 FILLCELL_X2 FILLER_36_61 ();
 FILLCELL_X4 FILLER_36_92 ();
 FILLCELL_X1 FILLER_36_96 ();
 FILLCELL_X32 FILLER_36_141 ();
 FILLCELL_X32 FILLER_36_173 ();
 FILLCELL_X32 FILLER_36_205 ();
 FILLCELL_X32 FILLER_36_237 ();
 FILLCELL_X16 FILLER_36_269 ();
 FILLCELL_X8 FILLER_36_285 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X4 FILLER_37_65 ();
 FILLCELL_X8 FILLER_37_88 ();
 FILLCELL_X4 FILLER_37_96 ();
 FILLCELL_X1 FILLER_37_100 ();
 FILLCELL_X8 FILLER_37_122 ();
 FILLCELL_X1 FILLER_37_130 ();
 FILLCELL_X8 FILLER_37_148 ();
 FILLCELL_X2 FILLER_37_159 ();
 FILLCELL_X32 FILLER_37_165 ();
 FILLCELL_X32 FILLER_37_197 ();
 FILLCELL_X32 FILLER_37_229 ();
 FILLCELL_X32 FILLER_37_261 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X8 FILLER_38_129 ();
 FILLCELL_X4 FILLER_38_137 ();
 FILLCELL_X2 FILLER_38_141 ();
 FILLCELL_X1 FILLER_38_143 ();
 FILLCELL_X4 FILLER_38_147 ();
 FILLCELL_X2 FILLER_38_154 ();
 FILLCELL_X1 FILLER_38_160 ();
 FILLCELL_X16 FILLER_38_165 ();
 FILLCELL_X4 FILLER_38_181 ();
 FILLCELL_X2 FILLER_38_185 ();
 FILLCELL_X1 FILLER_38_187 ();
 FILLCELL_X32 FILLER_38_194 ();
 FILLCELL_X32 FILLER_38_226 ();
 FILLCELL_X32 FILLER_38_258 ();
 FILLCELL_X2 FILLER_38_290 ();
 FILLCELL_X1 FILLER_38_292 ();
endmodule
