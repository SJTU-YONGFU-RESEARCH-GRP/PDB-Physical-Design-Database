module parameterized_updown_counter (clk,
    enable,
    overflow,
    rst_n,
    up_down,
    count);
 input clk;
 input enable;
 output overflow;
 input rst_n;
 input up_down;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net9;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _32_ (.I(net4),
    .ZN(_26_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _33_ (.I(net5),
    .ZN(_27_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _34_ (.I(_28_),
    .ZN(_05_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _35_ (.A1(net6),
    .A2(net7),
    .A3(_05_),
    .A4(net3),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _36_ (.A1(net2),
    .A2(_06_),
    .Z(_07_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _37_ (.A1(net6),
    .A2(net7),
    .A3(_30_),
    .A4(net3),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _38_ (.I0(_26_),
    .I1(_08_),
    .S(net2),
    .Z(_09_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _39_ (.A1(net4),
    .A2(_07_),
    .B(_09_),
    .ZN(_00_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _40_ (.A1(net3),
    .A2(_29_),
    .ZN(_10_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _41_ (.I0(net5),
    .I1(_10_),
    .S(net2),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _42_ (.I(net6),
    .ZN(_11_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _43_ (.I0(_28_),
    .I1(_30_),
    .S(net3),
    .Z(_12_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _44_ (.A1(net2),
    .A2(_12_),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _45_ (.A1(_11_),
    .A2(_13_),
    .ZN(_02_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _46_ (.A1(net6),
    .A2(net5),
    .A3(net4),
    .ZN(_14_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _47_ (.A1(net7),
    .A2(net3),
    .A3(_14_),
    .ZN(_15_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _48_ (.A1(net7),
    .A2(net2),
    .ZN(_16_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _49_ (.I(net3),
    .ZN(_17_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _50_ (.A1(net7),
    .A2(_17_),
    .A3(net2),
    .A4(_14_),
    .Z(_18_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _51_ (.A1(_16_),
    .A2(_18_),
    .Z(_19_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _52_ (.A1(_11_),
    .A2(net7),
    .A3(_27_),
    .A4(_26_),
    .Z(_20_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _53_ (.A1(net5),
    .A2(net4),
    .B(_30_),
    .ZN(_21_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _54_ (.A1(_11_),
    .A2(_21_),
    .B(net7),
    .ZN(_22_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _55_ (.A1(net3),
    .A2(net2),
    .A3(_20_),
    .A4(_22_),
    .Z(_23_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _56_ (.A1(_07_),
    .A2(_15_),
    .B(_19_),
    .C(_23_),
    .ZN(_03_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _57_ (.A1(net6),
    .A2(net7),
    .A3(_30_),
    .A4(net3),
    .ZN(_24_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _58_ (.A1(net2),
    .A2(net8),
    .ZN(_25_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _59_ (.A1(_07_),
    .A2(_24_),
    .B(_25_),
    .ZN(_04_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _60_ (.A(_26_),
    .B(_27_),
    .CO(_28_),
    .S(_29_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _61_ (.A(net4),
    .B(net5),
    .CO(_30_),
    .S(_31_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \overflow_reg$_DFFE_PN0P_  (.D(_04_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 hold1 (.I(net9),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_60 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input2 (.I(up_down),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net4),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net5),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net7),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net8),
    .Z(overflow));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_220 ();
endmodule
