module basic_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \rx_shift_reg[7] ;
 wire spi_clk_en;
 wire \state[0] ;
 wire \state[1] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net26;

 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _131_ (.A1(\bit_count[2] ),
    .A2(_114_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _132_ (.A1(\bit_count[3] ),
    .A2(_111_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _133_ (.I(\state[0] ),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _134_ (.A1(\state[1] ),
    .A2(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _135_ (.I(_113_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _136_ (.I(\bit_count[3] ),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _137_ (.A1(\bit_count[2] ),
    .A2(\bit_count[0] ),
    .A3(\bit_count[1] ),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _138_ (.I(_125_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _139_ (.A1(\bit_count[3] ),
    .A2(_117_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _140_ (.I(\state[1] ),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _141_ (.I(\bit_count[0] ),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _142_ (.I(net22),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _143_ (.A1(spi_clk_en),
    .A2(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _144_ (.A1(_035_),
    .A2(spi_clk_en),
    .A3(_037_),
    .A4(_036_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _145_ (.A1(\bit_count[0] ),
    .A2(_038_),
    .B(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _146_ (.A1(_035_),
    .A2(_036_),
    .B1(_040_),
    .B2(_112_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _147_ (.A1(_035_),
    .A2(spi_clk_en),
    .A3(_037_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _148_ (.A1(\bit_count[1] ),
    .A2(_038_),
    .B1(_041_),
    .B2(_115_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _149_ (.A1(\state[1] ),
    .A2(\bit_count[1] ),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _150_ (.A1(_112_),
    .A2(_042_),
    .B(_043_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _151_ (.I(_114_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _152_ (.I(spi_clk_en),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _153_ (.A1(\state[1] ),
    .A2(\bit_count[2] ),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _154_ (.A1(_044_),
    .A2(_045_),
    .A3(net22),
    .A4(_046_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _155_ (.A1(_044_),
    .A2(_045_),
    .A3(net22),
    .B(\bit_count[2] ),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _156_ (.A1(_047_),
    .A2(_048_),
    .B(_112_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _157_ (.A1(\state[1] ),
    .A2(\bit_count[2] ),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _158_ (.A1(_049_),
    .A2(_050_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _159_ (.A1(\bit_count[3] ),
    .A2(_038_),
    .B1(_041_),
    .B2(_119_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _160_ (.A1(_035_),
    .A2(_116_),
    .B1(_051_),
    .B2(_112_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _161_ (.I0(\rx_shift_reg[0] ),
    .I1(net13),
    .S(_113_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _162_ (.I0(\rx_shift_reg[1] ),
    .I1(net14),
    .S(_113_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _163_ (.I0(\rx_shift_reg[2] ),
    .I1(net15),
    .S(_113_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _164_ (.I0(\rx_shift_reg[3] ),
    .I1(net16),
    .S(_113_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _165_ (.I0(\rx_shift_reg[4] ),
    .I1(net17),
    .S(_113_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _166_ (.I0(\rx_shift_reg[5] ),
    .I1(net18),
    .S(_113_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _167_ (.I0(\rx_shift_reg[6] ),
    .I1(net19),
    .S(_113_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _168_ (.I0(\rx_shift_reg[7] ),
    .I1(net20),
    .S(_113_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _169_ (.A1(_118_),
    .A2(_129_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _170_ (.A1(_122_),
    .A2(_130_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _171_ (.A1(_118_),
    .A2(_129_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _172_ (.A1(_122_),
    .A2(_130_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _173_ (.A1(_052_),
    .A2(_053_),
    .B1(_054_),
    .B2(_055_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _174_ (.A1(_126_),
    .A2(_123_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _175_ (.A1(\bit_count[0] ),
    .A2(_057_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _176_ (.A1(_035_),
    .A2(\state[0] ),
    .A3(spi_clk_en),
    .A4(_037_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _177_ (.I(_115_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _178_ (.A1(\bit_count[2] ),
    .A2(_114_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _179_ (.A1(_122_),
    .A2(_060_),
    .A3(_119_),
    .A4(_061_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _180_ (.A1(_056_),
    .A2(_058_),
    .A3(_059_),
    .A4(_062_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _181_ (.I0(\rx_shift_reg[0] ),
    .I1(net3),
    .S(_063_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _182_ (.I(_059_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _183_ (.I(_119_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _184_ (.A1(_115_),
    .A2(_065_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _185_ (.A1(_064_),
    .A2(_066_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _186_ (.A1(_118_),
    .A2(_129_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _187_ (.A1(_122_),
    .A2(_130_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _188_ (.A1(_036_),
    .A2(net3),
    .A3(_057_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _189_ (.A1(_068_),
    .A2(_069_),
    .A3(_070_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _190_ (.A1(\bit_count[2] ),
    .A2(_114_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _191_ (.A1(_116_),
    .A2(_036_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _192_ (.A1(_064_),
    .A2(_072_),
    .A3(_066_),
    .A4(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _193_ (.I(\rx_shift_reg[1] ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _194_ (.A1(_061_),
    .A2(_067_),
    .A3(_071_),
    .B1(_074_),
    .B2(_075_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _195_ (.A1(\bit_count[0] ),
    .A2(_068_),
    .A3(_069_),
    .A4(_057_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _196_ (.A1(_064_),
    .A2(_072_),
    .A3(_066_),
    .A4(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _197_ (.I0(\rx_shift_reg[2] ),
    .I1(net3),
    .S(_077_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _198_ (.A1(_060_),
    .A2(_065_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _199_ (.A1(_064_),
    .A2(_078_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _200_ (.A1(_064_),
    .A2(_072_),
    .A3(_073_),
    .A4(_078_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _201_ (.I(\rx_shift_reg[3] ),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _202_ (.A1(_061_),
    .A2(_071_),
    .A3(_079_),
    .B1(_080_),
    .B2(_081_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _203_ (.A1(_064_),
    .A2(_072_),
    .A3(_076_),
    .A4(_078_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _204_ (.I0(\rx_shift_reg[4] ),
    .I1(net3),
    .S(_082_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _205_ (.A1(_064_),
    .A2(_061_),
    .A3(_066_),
    .A4(_073_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _206_ (.I(\rx_shift_reg[5] ),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _207_ (.A1(_072_),
    .A2(_067_),
    .A3(_071_),
    .B1(_083_),
    .B2(_084_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _208_ (.A1(_064_),
    .A2(_061_),
    .A3(_066_),
    .A4(_076_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(\rx_shift_reg[6] ),
    .I1(net3),
    .S(_085_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _210_ (.A1(_064_),
    .A2(_061_),
    .A3(_073_),
    .A4(_078_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _211_ (.I(\rx_shift_reg[7] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _212_ (.A1(_072_),
    .A2(_071_),
    .A3(_079_),
    .B1(_086_),
    .B2(_087_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _213_ (.A1(_045_),
    .A2(net22),
    .B(_041_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _214_ (.A1(_035_),
    .A2(_037_),
    .B1(_088_),
    .B2(_112_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _215_ (.A1(_112_),
    .A2(net12),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _216_ (.A1(\state[0] ),
    .A2(spi_clk_en),
    .A3(net22),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _217_ (.I(_090_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _218_ (.A1(_089_),
    .A2(_091_),
    .B(\state[1] ),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _219_ (.A1(\bit_count[3] ),
    .A2(_111_),
    .B(_037_),
    .C(\state[0] ),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _220_ (.A1(_035_),
    .A2(_093_),
    .B(_045_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _221_ (.A1(_092_),
    .A2(_094_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _222_ (.A1(_035_),
    .A2(net12),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _223_ (.I0(net23),
    .I1(_095_),
    .S(_112_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _224_ (.I0(net11),
    .I1(\tx_shift_reg[6] ),
    .S(\state[0] ),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _225_ (.A1(_121_),
    .A2(_090_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _226_ (.A1(_089_),
    .A2(_097_),
    .B(\state[1] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _227_ (.I0(net24),
    .I1(_096_),
    .S(_098_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _228_ (.A1(\bit_count[3] ),
    .A2(_111_),
    .A3(_038_),
    .B(\state[0] ),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _229_ (.A1(_089_),
    .A2(_099_),
    .B(\state[1] ),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _230_ (.A1(_125_),
    .A2(_064_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _231_ (.I(net12),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _232_ (.A1(_035_),
    .A2(_112_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _233_ (.I0(_100_),
    .I1(net25),
    .S(_101_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _234_ (.I(\tx_shift_reg[0] ),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _235_ (.A1(net12),
    .A2(net4),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _236_ (.A1(_102_),
    .A2(_092_),
    .B1(_101_),
    .B2(_103_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _237_ (.A1(_035_),
    .A2(\state[0] ),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _238_ (.I0(net5),
    .I1(\tx_shift_reg[0] ),
    .S(_104_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _239_ (.I0(\tx_shift_reg[1] ),
    .I1(_105_),
    .S(_092_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _240_ (.I0(net6),
    .I1(\tx_shift_reg[1] ),
    .S(_104_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _241_ (.I0(\tx_shift_reg[2] ),
    .I1(_106_),
    .S(_092_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _242_ (.I0(net7),
    .I1(\tx_shift_reg[2] ),
    .S(_104_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _243_ (.I0(\tx_shift_reg[3] ),
    .I1(_107_),
    .S(_092_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _244_ (.I0(net8),
    .I1(\tx_shift_reg[3] ),
    .S(_104_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _245_ (.I0(\tx_shift_reg[4] ),
    .I1(_108_),
    .S(_092_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _246_ (.I0(net9),
    .I1(\tx_shift_reg[4] ),
    .S(_104_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _247_ (.I0(\tx_shift_reg[5] ),
    .I1(_109_),
    .S(_092_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _248_ (.I0(net10),
    .I1(\tx_shift_reg[5] ),
    .S(_104_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _249_ (.I0(\tx_shift_reg[6] ),
    .I1(_110_),
    .S(_092_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _250_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_114_),
    .S(_115_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _251_ (.A(_116_),
    .B(_117_),
    .CO(_118_),
    .S(_119_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _252_ (.A(_116_),
    .B(_120_),
    .CO(_121_),
    .S(_122_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _253_ (.A(\bit_count[3] ),
    .B(_120_),
    .CO(_123_),
    .S(_124_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _254_ (.A(\bit_count[3] ),
    .B(_125_),
    .CO(_126_),
    .S(_127_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _255_ (.A(_116_),
    .B(_128_),
    .CO(_129_),
    .S(_130_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[1]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[2]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[3]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[0]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[1]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[2]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[3]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rx_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[4]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[5]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[6]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[7]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_valid$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk_en$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(spi_clk_en));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \spi_cs_n$_DFFE_PN1P_  (.D(_023_),
    .SETN(net2),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_mosi$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[0]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[1]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx_ready$_DFFE_PN1P_  (.D(_027_),
    .SETN(net2),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[0]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[1]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[2]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[3]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[4]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[5]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[6]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net26),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input2 (.I(spi_miso),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(tx_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(tx_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(tx_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(tx_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(tx_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(tx_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tx_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input11 (.I(tx_valid),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(rx_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(rx_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rx_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rx_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rx_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rx_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rx_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(spi_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(spi_cs_n));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(spi_mosi));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(tx_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload1 (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_248 ();
endmodule
