module piso_register (clk,
    load,
    rst_n,
    serial_out,
    parallel_in);
 input clk;
 input load;
 input rst_n;
 output serial_out;
 input [7:0] parallel_in;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire \shift_reg[1] ;
 wire \shift_reg[2] ;
 wire \shift_reg[3] ;
 wire \shift_reg[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X2 _28_ (.A(rst_n),
    .Z(_11_));
 BUF_X4 _29_ (.A(load),
    .Z(_12_));
 MUX2_X1 _30_ (.A(_01_),
    .B(net6),
    .S(_12_),
    .Z(_13_));
 AND2_X1 _31_ (.A1(_11_),
    .A2(_13_),
    .ZN(_03_));
 MUX2_X1 _32_ (.A(_02_),
    .B(net7),
    .S(_12_),
    .Z(_14_));
 AND2_X1 _33_ (.A1(_11_),
    .A2(_14_),
    .ZN(_04_));
 AND3_X1 _34_ (.A1(_11_),
    .A2(_12_),
    .A3(net8),
    .ZN(_05_));
 MUX2_X1 _35_ (.A(\shift_reg[1] ),
    .B(net1),
    .S(_12_),
    .Z(_15_));
 AND2_X1 _36_ (.A1(_11_),
    .A2(_15_),
    .ZN(_06_));
 MUX2_X1 _37_ (.A(\shift_reg[2] ),
    .B(net2),
    .S(_12_),
    .Z(_16_));
 AND2_X1 _38_ (.A1(_11_),
    .A2(_16_),
    .ZN(_07_));
 MUX2_X1 _39_ (.A(\shift_reg[3] ),
    .B(net3),
    .S(_12_),
    .Z(_17_));
 AND2_X1 _40_ (.A1(_11_),
    .A2(_17_),
    .ZN(_08_));
 MUX2_X1 _41_ (.A(\shift_reg[4] ),
    .B(net4),
    .S(_12_),
    .Z(_18_));
 AND2_X1 _42_ (.A1(_11_),
    .A2(_18_),
    .ZN(_09_));
 MUX2_X1 _43_ (.A(_00_),
    .B(net5),
    .S(_12_),
    .Z(_19_));
 AND2_X1 _44_ (.A1(_11_),
    .A2(_19_),
    .ZN(_10_));
 DFF_X1 _45_ (.D(_03_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_00_),
    .QN(_27_));
 DFF_X1 _46_ (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_01_),
    .QN(_26_));
 DFF_X1 _47_ (.D(_05_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_02_),
    .QN(_25_));
 DFF_X1 \serial_out$_SDFF_PN0_  (.D(_06_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net9),
    .QN(_24_));
 DFF_X1 \shift_reg[1]$_SDFF_PN0_  (.D(_07_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[1] ),
    .QN(_23_));
 DFF_X1 \shift_reg[2]$_SDFF_PN0_  (.D(_08_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[2] ),
    .QN(_22_));
 DFF_X1 \shift_reg[3]$_SDFF_PN0_  (.D(_09_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[3] ),
    .QN(_21_));
 DFF_X1 \shift_reg[4]$_SDFF_PN0_  (.D(_10_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[4] ),
    .QN(_20_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_49 ();
 BUF_X1 input1 (.A(parallel_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(parallel_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(parallel_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(parallel_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(parallel_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(parallel_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(parallel_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(parallel_in[7]),
    .Z(net8));
 BUF_X1 output9 (.A(net9),
    .Z(serial_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_84 ();
 FILLCELL_X32 FILLER_0_116 ();
 FILLCELL_X32 FILLER_0_148 ();
 FILLCELL_X4 FILLER_0_180 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X16 FILLER_1_161 ();
 FILLCELL_X4 FILLER_1_177 ();
 FILLCELL_X2 FILLER_1_181 ();
 FILLCELL_X1 FILLER_1_183 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X16 FILLER_2_161 ();
 FILLCELL_X4 FILLER_2_177 ();
 FILLCELL_X2 FILLER_2_181 ();
 FILLCELL_X1 FILLER_2_183 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X16 FILLER_3_161 ();
 FILLCELL_X4 FILLER_3_177 ();
 FILLCELL_X2 FILLER_3_181 ();
 FILLCELL_X1 FILLER_3_183 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X16 FILLER_4_161 ();
 FILLCELL_X4 FILLER_4_177 ();
 FILLCELL_X2 FILLER_4_181 ();
 FILLCELL_X1 FILLER_4_183 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X16 FILLER_5_161 ();
 FILLCELL_X4 FILLER_5_177 ();
 FILLCELL_X2 FILLER_5_181 ();
 FILLCELL_X1 FILLER_5_183 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X4 FILLER_6_177 ();
 FILLCELL_X2 FILLER_6_181 ();
 FILLCELL_X1 FILLER_6_183 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X16 FILLER_7_161 ();
 FILLCELL_X4 FILLER_7_177 ();
 FILLCELL_X2 FILLER_7_181 ();
 FILLCELL_X1 FILLER_7_183 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X16 FILLER_8_161 ();
 FILLCELL_X4 FILLER_8_177 ();
 FILLCELL_X2 FILLER_8_181 ();
 FILLCELL_X1 FILLER_8_183 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X16 FILLER_9_161 ();
 FILLCELL_X4 FILLER_9_177 ();
 FILLCELL_X2 FILLER_9_181 ();
 FILLCELL_X1 FILLER_9_183 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_14 ();
 FILLCELL_X32 FILLER_10_46 ();
 FILLCELL_X32 FILLER_10_78 ();
 FILLCELL_X32 FILLER_10_110 ();
 FILLCELL_X4 FILLER_10_142 ();
 FILLCELL_X32 FILLER_10_149 ();
 FILLCELL_X2 FILLER_10_181 ();
 FILLCELL_X1 FILLER_10_183 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_9 ();
 FILLCELL_X2 FILLER_11_16 ();
 FILLCELL_X1 FILLER_11_18 ();
 FILLCELL_X4 FILLER_11_22 ();
 FILLCELL_X2 FILLER_11_43 ();
 FILLCELL_X4 FILLER_11_52 ();
 FILLCELL_X1 FILLER_11_60 ();
 FILLCELL_X2 FILLER_11_85 ();
 FILLCELL_X2 FILLER_11_108 ();
 FILLCELL_X32 FILLER_11_117 ();
 FILLCELL_X32 FILLER_11_149 ();
 FILLCELL_X2 FILLER_11_181 ();
 FILLCELL_X1 FILLER_11_183 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_6 ();
 FILLCELL_X2 FILLER_12_25 ();
 FILLCELL_X32 FILLER_12_31 ();
 FILLCELL_X32 FILLER_12_63 ();
 FILLCELL_X2 FILLER_12_95 ();
 FILLCELL_X1 FILLER_12_97 ();
 FILLCELL_X4 FILLER_12_102 ();
 FILLCELL_X2 FILLER_12_106 ();
 FILLCELL_X1 FILLER_12_108 ();
 FILLCELL_X32 FILLER_12_113 ();
 FILLCELL_X32 FILLER_12_145 ();
 FILLCELL_X4 FILLER_12_177 ();
 FILLCELL_X2 FILLER_12_181 ();
 FILLCELL_X1 FILLER_12_183 ();
 FILLCELL_X2 FILLER_13_4 ();
 FILLCELL_X1 FILLER_13_16 ();
 FILLCELL_X1 FILLER_13_21 ();
 FILLCELL_X8 FILLER_13_29 ();
 FILLCELL_X4 FILLER_13_37 ();
 FILLCELL_X2 FILLER_13_41 ();
 FILLCELL_X16 FILLER_13_48 ();
 FILLCELL_X8 FILLER_13_64 ();
 FILLCELL_X4 FILLER_13_72 ();
 FILLCELL_X1 FILLER_13_76 ();
 FILLCELL_X8 FILLER_13_82 ();
 FILLCELL_X4 FILLER_13_90 ();
 FILLCELL_X1 FILLER_13_94 ();
 FILLCELL_X1 FILLER_13_128 ();
 FILLCELL_X8 FILLER_13_146 ();
 FILLCELL_X4 FILLER_13_154 ();
 FILLCELL_X2 FILLER_13_158 ();
 FILLCELL_X16 FILLER_13_163 ();
 FILLCELL_X4 FILLER_13_179 ();
 FILLCELL_X1 FILLER_13_183 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X2 FILLER_14_13 ();
 FILLCELL_X32 FILLER_14_32 ();
 FILLCELL_X32 FILLER_14_64 ();
 FILLCELL_X8 FILLER_14_96 ();
 FILLCELL_X2 FILLER_14_104 ();
 FILLCELL_X16 FILLER_14_130 ();
 FILLCELL_X4 FILLER_14_146 ();
 FILLCELL_X1 FILLER_14_150 ();
 FILLCELL_X4 FILLER_14_154 ();
 FILLCELL_X2 FILLER_14_158 ();
 FILLCELL_X1 FILLER_14_160 ();
 FILLCELL_X16 FILLER_14_164 ();
 FILLCELL_X4 FILLER_14_180 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X16 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_177 ();
 FILLCELL_X2 FILLER_15_181 ();
 FILLCELL_X1 FILLER_15_183 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X16 FILLER_16_161 ();
 FILLCELL_X4 FILLER_16_177 ();
 FILLCELL_X2 FILLER_16_181 ();
 FILLCELL_X1 FILLER_16_183 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X16 FILLER_17_161 ();
 FILLCELL_X4 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_181 ();
 FILLCELL_X1 FILLER_17_183 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X16 FILLER_18_161 ();
 FILLCELL_X4 FILLER_18_177 ();
 FILLCELL_X2 FILLER_18_181 ();
 FILLCELL_X1 FILLER_18_183 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_177 ();
 FILLCELL_X2 FILLER_19_181 ();
 FILLCELL_X1 FILLER_19_183 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X16 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_177 ();
 FILLCELL_X2 FILLER_20_181 ();
 FILLCELL_X1 FILLER_20_183 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_177 ();
 FILLCELL_X2 FILLER_21_181 ();
 FILLCELL_X1 FILLER_21_183 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X4 FILLER_22_177 ();
 FILLCELL_X2 FILLER_22_181 ();
 FILLCELL_X1 FILLER_22_183 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X16 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_177 ();
 FILLCELL_X2 FILLER_23_181 ();
 FILLCELL_X1 FILLER_23_183 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X16 FILLER_24_161 ();
 FILLCELL_X4 FILLER_24_177 ();
 FILLCELL_X2 FILLER_24_181 ();
 FILLCELL_X1 FILLER_24_183 ();
endmodule
