module uart (clk,
    m_axis_tready,
    m_axis_tvalid,
    rst,
    rx_busy,
    rx_frame_error,
    rx_overrun_error,
    rxd,
    s_axis_tready,
    s_axis_tvalid,
    tx_busy,
    txd,
    m_axis_tdata,
    prescale,
    s_axis_tdata);
 input clk;
 input m_axis_tready;
 output m_axis_tvalid;
 input rst;
 output rx_busy;
 output rx_frame_error;
 output rx_overrun_error;
 input rxd;
 output s_axis_tready;
 input s_axis_tvalid;
 output tx_busy;
 output txd;
 output [7:0] m_axis_tdata;
 input [15:0] prescale;
 input [7:0] s_axis_tdata;

 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire \uart_tx_inst/_000_ ;
 wire \uart_tx_inst/_001_ ;
 wire \uart_tx_inst/_002_ ;
 wire \uart_tx_inst/_003_ ;
 wire \uart_tx_inst/_004_ ;
 wire \uart_tx_inst/_005_ ;
 wire \uart_tx_inst/_006_ ;
 wire \uart_tx_inst/_007_ ;
 wire \uart_tx_inst/_008_ ;
 wire \uart_tx_inst/_009_ ;
 wire \uart_tx_inst/_010_ ;
 wire \uart_tx_inst/_011_ ;
 wire \uart_tx_inst/_012_ ;
 wire \uart_tx_inst/_013_ ;
 wire \uart_tx_inst/_014_ ;
 wire \uart_tx_inst/_015_ ;
 wire \uart_tx_inst/_016_ ;
 wire \uart_tx_inst/_017_ ;
 wire \uart_tx_inst/_018_ ;
 wire \uart_tx_inst/_019_ ;
 wire \uart_tx_inst/_020_ ;
 wire \uart_tx_inst/_021_ ;
 wire \uart_tx_inst/_022_ ;
 wire \uart_tx_inst/_023_ ;
 wire \uart_tx_inst/_024_ ;
 wire \uart_tx_inst/_025_ ;
 wire \uart_tx_inst/_026_ ;
 wire \uart_tx_inst/_027_ ;
 wire \uart_tx_inst/_028_ ;
 wire \uart_tx_inst/_029_ ;
 wire \uart_tx_inst/_030_ ;
 wire \uart_tx_inst/_031_ ;
 wire \uart_tx_inst/_032_ ;
 wire \uart_tx_inst/_033_ ;
 wire \uart_tx_inst/_034_ ;
 wire \uart_tx_inst/_035_ ;
 wire \uart_tx_inst/_036_ ;
 wire net5;
 wire \uart_tx_inst/_038_ ;
 wire \uart_tx_inst/_039_ ;
 wire \uart_tx_inst/_040_ ;
 wire \uart_tx_inst/_041_ ;
 wire \uart_tx_inst/_042_ ;
 wire \uart_tx_inst/_043_ ;
 wire \uart_tx_inst/_044_ ;
 wire \uart_tx_inst/_045_ ;
 wire \uart_tx_inst/_046_ ;
 wire \uart_tx_inst/_047_ ;
 wire \uart_tx_inst/_048_ ;
 wire \uart_tx_inst/_049_ ;
 wire \uart_tx_inst/_050_ ;
 wire \uart_tx_inst/_051_ ;
 wire \uart_tx_inst/_052_ ;
 wire net4;
 wire \uart_tx_inst/_054_ ;
 wire \uart_tx_inst/_055_ ;
 wire \uart_tx_inst/_056_ ;
 wire \uart_tx_inst/_057_ ;
 wire \uart_tx_inst/_058_ ;
 wire \uart_tx_inst/_059_ ;
 wire \uart_tx_inst/_060_ ;
 wire net3;
 wire \uart_tx_inst/_062_ ;
 wire \uart_tx_inst/_063_ ;
 wire \uart_tx_inst/_064_ ;
 wire \uart_tx_inst/_065_ ;
 wire \uart_tx_inst/_066_ ;
 wire \uart_tx_inst/_067_ ;
 wire net2;
 wire \uart_tx_inst/_069_ ;
 wire \uart_tx_inst/_070_ ;
 wire \uart_tx_inst/_071_ ;
 wire \uart_tx_inst/_072_ ;
 wire \uart_tx_inst/_073_ ;
 wire \uart_tx_inst/_074_ ;
 wire \uart_tx_inst/_075_ ;
 wire \uart_tx_inst/_076_ ;
 wire \uart_tx_inst/_077_ ;
 wire \uart_tx_inst/_078_ ;
 wire \uart_tx_inst/_079_ ;
 wire \uart_tx_inst/_080_ ;
 wire \uart_tx_inst/_081_ ;
 wire \uart_tx_inst/_082_ ;
 wire \uart_tx_inst/_083_ ;
 wire \uart_tx_inst/_084_ ;
 wire \uart_tx_inst/_085_ ;
 wire \uart_tx_inst/_086_ ;
 wire net1;
 wire \uart_tx_inst/_088_ ;
 wire \uart_tx_inst/_089_ ;
 wire \uart_tx_inst/_090_ ;
 wire \uart_tx_inst/_091_ ;
 wire \uart_tx_inst/_092_ ;
 wire \uart_tx_inst/_093_ ;
 wire \uart_tx_inst/_094_ ;
 wire \uart_tx_inst/_095_ ;
 wire \uart_tx_inst/_096_ ;
 wire \uart_tx_inst/_097_ ;
 wire \uart_tx_inst/_098_ ;
 wire \uart_tx_inst/_099_ ;
 wire \uart_tx_inst/_100_ ;
 wire \uart_tx_inst/_101_ ;
 wire \uart_tx_inst/_102_ ;
 wire \uart_tx_inst/_103_ ;
 wire \uart_tx_inst/_104_ ;
 wire \uart_tx_inst/_105_ ;
 wire \uart_tx_inst/_106_ ;
 wire \uart_tx_inst/_107_ ;
 wire \uart_tx_inst/_108_ ;
 wire \uart_tx_inst/_109_ ;
 wire \uart_tx_inst/_110_ ;
 wire \uart_tx_inst/_111_ ;
 wire \uart_tx_inst/_112_ ;
 wire \uart_tx_inst/_113_ ;
 wire \uart_tx_inst/_114_ ;
 wire \uart_tx_inst/_115_ ;
 wire \uart_tx_inst/_116_ ;
 wire \uart_tx_inst/_117_ ;
 wire \uart_tx_inst/_118_ ;
 wire \uart_tx_inst/_119_ ;
 wire \uart_tx_inst/_120_ ;
 wire \uart_tx_inst/_121_ ;
 wire \uart_tx_inst/_122_ ;
 wire \uart_tx_inst/_123_ ;
 wire \uart_tx_inst/_124_ ;
 wire \uart_tx_inst/_125_ ;
 wire \uart_tx_inst/_126_ ;
 wire \uart_tx_inst/_127_ ;
 wire \uart_tx_inst/_128_ ;
 wire \uart_tx_inst/_129_ ;
 wire \uart_tx_inst/_130_ ;
 wire \uart_tx_inst/_131_ ;
 wire \uart_tx_inst/_132_ ;
 wire \uart_tx_inst/_133_ ;
 wire \uart_tx_inst/_134_ ;
 wire \uart_tx_inst/_135_ ;
 wire \uart_tx_inst/_136_ ;
 wire \uart_tx_inst/_137_ ;
 wire \uart_tx_inst/_138_ ;
 wire \uart_tx_inst/_139_ ;
 wire \uart_tx_inst/_140_ ;
 wire \uart_tx_inst/_141_ ;
 wire \uart_tx_inst/_142_ ;
 wire \uart_tx_inst/_143_ ;
 wire \uart_tx_inst/_144_ ;
 wire \uart_tx_inst/_145_ ;
 wire \uart_tx_inst/_146_ ;
 wire \uart_tx_inst/_147_ ;
 wire \uart_tx_inst/_148_ ;
 wire \uart_tx_inst/_149_ ;
 wire \uart_tx_inst/_150_ ;
 wire \uart_tx_inst/_151_ ;
 wire \uart_tx_inst/_152_ ;
 wire \uart_tx_inst/_153_ ;
 wire \uart_tx_inst/_154_ ;
 wire \uart_tx_inst/_155_ ;
 wire \uart_tx_inst/_156_ ;
 wire \uart_tx_inst/_157_ ;
 wire \uart_tx_inst/_158_ ;
 wire \uart_tx_inst/_159_ ;
 wire \uart_tx_inst/_160_ ;
 wire \uart_tx_inst/_161_ ;
 wire \uart_tx_inst/_162_ ;
 wire \uart_tx_inst/_163_ ;
 wire \uart_tx_inst/_164_ ;
 wire \uart_tx_inst/_165_ ;
 wire \uart_tx_inst/_166_ ;
 wire \uart_tx_inst/_167_ ;
 wire \uart_tx_inst/_168_ ;
 wire \uart_tx_inst/_169_ ;
 wire \uart_tx_inst/_170_ ;
 wire \uart_tx_inst/_171_ ;
 wire \uart_tx_inst/_172_ ;
 wire \uart_tx_inst/_173_ ;
 wire \uart_tx_inst/_174_ ;
 wire \uart_tx_inst/_175_ ;
 wire \uart_tx_inst/_176_ ;
 wire \uart_tx_inst/_177_ ;
 wire \uart_tx_inst/_178_ ;
 wire \uart_tx_inst/_179_ ;
 wire \uart_tx_inst/_180_ ;
 wire \uart_tx_inst/_181_ ;
 wire \uart_tx_inst/_182_ ;
 wire \uart_tx_inst/_183_ ;
 wire \uart_tx_inst/_184_ ;
 wire \uart_tx_inst/_185_ ;
 wire \uart_tx_inst/_186_ ;
 wire \uart_tx_inst/_187_ ;
 wire \uart_tx_inst/_188_ ;
 wire \uart_tx_inst/_189_ ;
 wire \uart_tx_inst/_190_ ;
 wire \uart_tx_inst/_191_ ;
 wire \uart_tx_inst/_192_ ;
 wire \uart_tx_inst/bit_cnt[0] ;
 wire \uart_tx_inst/bit_cnt[1] ;
 wire \uart_tx_inst/bit_cnt[2] ;
 wire \uart_tx_inst/bit_cnt[3] ;
 wire \uart_tx_inst/data_reg[0] ;
 wire \uart_tx_inst/data_reg[1] ;
 wire \uart_tx_inst/data_reg[2] ;
 wire \uart_tx_inst/data_reg[3] ;
 wire \uart_tx_inst/data_reg[4] ;
 wire \uart_tx_inst/data_reg[5] ;
 wire \uart_tx_inst/data_reg[6] ;
 wire \uart_tx_inst/data_reg[7] ;
 wire \uart_tx_inst/data_reg[8] ;
 wire \uart_tx_inst/prescale_reg[0] ;
 wire \uart_tx_inst/prescale_reg[10] ;
 wire \uart_tx_inst/prescale_reg[11] ;
 wire \uart_tx_inst/prescale_reg[12] ;
 wire \uart_tx_inst/prescale_reg[13] ;
 wire \uart_tx_inst/prescale_reg[14] ;
 wire \uart_tx_inst/prescale_reg[15] ;
 wire \uart_tx_inst/prescale_reg[16] ;
 wire \uart_tx_inst/prescale_reg[17] ;
 wire \uart_tx_inst/prescale_reg[18] ;
 wire \uart_tx_inst/prescale_reg[1] ;
 wire \uart_tx_inst/prescale_reg[2] ;
 wire \uart_tx_inst/prescale_reg[3] ;
 wire \uart_tx_inst/prescale_reg[4] ;
 wire \uart_tx_inst/prescale_reg[5] ;
 wire \uart_tx_inst/prescale_reg[6] ;
 wire \uart_tx_inst/prescale_reg[7] ;
 wire \uart_tx_inst/prescale_reg[8] ;
 wire \uart_tx_inst/prescale_reg[9] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire clk_regs;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_2_0__leaf_clk_regs;
 wire clknet_2_1__leaf_clk_regs;
 wire clknet_2_2__leaf_clk_regs;
 wire clknet_2_3__leaf_clk_regs;
 wire delaynet_0_clk;
 wire [0:0] \uart_tx_inst/_193_ ;
 wire [0:0] \uart_tx_inst/_194_ ;
 wire [0:0] \uart_tx_inst/_195_ ;
 wire [0:0] \uart_tx_inst/_196_ ;
 wire [0:0] \uart_tx_inst/_197_ ;
 wire [0:0] \uart_tx_inst/_198_ ;
 wire [0:0] \uart_tx_inst/_199_ ;
 wire [0:0] \uart_tx_inst/_200_ ;
 wire [0:0] \uart_tx_inst/_201_ ;
 wire [0:0] \uart_tx_inst/_202_ ;
 wire [0:0] \uart_tx_inst/_203_ ;
 wire [0:0] \uart_tx_inst/_204_ ;
 wire [0:0] \uart_tx_inst/_205_ ;
 wire [0:0] \uart_tx_inst/_206_ ;

 uart_rx uart_rx_inst (.busy(net38),
    .clk(clknet_1_0__leaf_clk),
    .frame_error(net39),
    .m_axis_tready(net1),
    .m_axis_tvalid(net37),
    .overrun_error(net40),
    .rst(net18),
    .rxd(net19),
    .m_axis_tdata({net36,
    net35,
    net34,
    net33,
    net32,
    net31,
    net30,
    net29}),
    .prescale({net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net17,
    net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9,
    net2}));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_207_  (.I(\uart_tx_inst/prescale_reg[0] ),
    .ZN(\uart_tx_inst/_193_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_208_  (.I(net2),
    .ZN(\uart_tx_inst/_197_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 \uart_tx_inst/_209_  (.I(\uart_tx_inst/bit_cnt[0] ),
    .ZN(\uart_tx_inst/_201_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_210_  (.I(\uart_tx_inst/prescale_reg[1] ),
    .ZN(\uart_tx_inst/_194_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_211_  (.I(net9),
    .ZN(\uart_tx_inst/_198_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_212_  (.I(\uart_tx_inst/bit_cnt[1] ),
    .ZN(\uart_tx_inst/_202_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 \uart_tx_inst/_213_  (.A1(\uart_tx_inst/bit_cnt[3] ),
    .A2(\uart_tx_inst/bit_cnt[2] ),
    .ZN(\uart_tx_inst/_035_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 \uart_tx_inst/_214_  (.A1(\uart_tx_inst/_203_ [0]),
    .A2(\uart_tx_inst/_035_ ),
    .Z(\uart_tx_inst/_036_ ));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input5 (.I(prescale[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_216_  (.I0(\uart_tx_inst/data_reg[1] ),
    .I1(net20),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_038_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 \uart_tx_inst/_217_  (.I(net18),
    .ZN(\uart_tx_inst/_039_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 \uart_tx_inst/_218_  (.A1(\uart_tx_inst/prescale_reg[0] ),
    .A2(\uart_tx_inst/prescale_reg[1] ),
    .Z(\uart_tx_inst/_040_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_219_  (.A1(\uart_tx_inst/prescale_reg[3] ),
    .A2(\uart_tx_inst/prescale_reg[2] ),
    .A3(\uart_tx_inst/prescale_reg[5] ),
    .A4(\uart_tx_inst/prescale_reg[4] ),
    .Z(\uart_tx_inst/_041_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 \uart_tx_inst/_220_  (.A1(\uart_tx_inst/prescale_reg[7] ),
    .A2(\uart_tx_inst/prescale_reg[6] ),
    .A3(\uart_tx_inst/prescale_reg[9] ),
    .A4(\uart_tx_inst/prescale_reg[8] ),
    .Z(\uart_tx_inst/_042_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 \uart_tx_inst/_221_  (.A1(\uart_tx_inst/prescale_reg[10] ),
    .A2(\uart_tx_inst/_040_ ),
    .A3(\uart_tx_inst/_041_ ),
    .A4(\uart_tx_inst/_042_ ),
    .Z(\uart_tx_inst/_043_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 \uart_tx_inst/_222_  (.A1(\uart_tx_inst/prescale_reg[15] ),
    .A2(\uart_tx_inst/prescale_reg[16] ),
    .Z(\uart_tx_inst/_044_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 \uart_tx_inst/_223_  (.A1(\uart_tx_inst/prescale_reg[14] ),
    .A2(\uart_tx_inst/prescale_reg[13] ),
    .A3(\uart_tx_inst/prescale_reg[12] ),
    .A4(\uart_tx_inst/prescale_reg[11] ),
    .Z(\uart_tx_inst/_045_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 \uart_tx_inst/_224_  (.A1(\uart_tx_inst/_043_ ),
    .A2(\uart_tx_inst/_044_ ),
    .A3(\uart_tx_inst/_045_ ),
    .ZN(\uart_tx_inst/_046_ ));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 \uart_tx_inst/_225_  (.I(net28),
    .ZN(\uart_tx_inst/_047_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_226_  (.I(\uart_tx_inst/_203_ [0]),
    .ZN(\uart_tx_inst/_048_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_227_  (.I0(\uart_tx_inst/_047_ ),
    .I1(\uart_tx_inst/_205_ [0]),
    .S(\uart_tx_inst/_048_ ),
    .Z(\uart_tx_inst/_049_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_228_  (.A1(\uart_tx_inst/_035_ ),
    .A2(\uart_tx_inst/_049_ ),
    .ZN(\uart_tx_inst/_050_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 \uart_tx_inst/_229_  (.A1(\uart_tx_inst/prescale_reg[17] ),
    .A2(\uart_tx_inst/prescale_reg[18] ),
    .ZN(\uart_tx_inst/_051_ ));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 \uart_tx_inst/_230_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_046_ ),
    .A3(\uart_tx_inst/_050_ ),
    .A4(\uart_tx_inst/_051_ ),
    .Z(\uart_tx_inst/_052_ ));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input4 (.I(prescale[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_232_  (.I0(\uart_tx_inst/data_reg[0] ),
    .I1(\uart_tx_inst/_038_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_005_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_233_  (.I0(\uart_tx_inst/data_reg[2] ),
    .I1(net21),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_054_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_234_  (.I0(\uart_tx_inst/data_reg[1] ),
    .I1(\uart_tx_inst/_054_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_006_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_235_  (.I0(\uart_tx_inst/data_reg[3] ),
    .I1(net22),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_055_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_236_  (.I0(\uart_tx_inst/data_reg[2] ),
    .I1(\uart_tx_inst/_055_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_007_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_237_  (.I0(\uart_tx_inst/data_reg[4] ),
    .I1(net23),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_056_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_238_  (.I0(\uart_tx_inst/data_reg[3] ),
    .I1(\uart_tx_inst/_056_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_008_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_239_  (.I0(\uart_tx_inst/data_reg[5] ),
    .I1(net24),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_057_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_240_  (.I0(\uart_tx_inst/data_reg[4] ),
    .I1(\uart_tx_inst/_057_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_009_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_241_  (.I0(\uart_tx_inst/data_reg[6] ),
    .I1(net25),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_058_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_242_  (.I0(\uart_tx_inst/data_reg[5] ),
    .I1(\uart_tx_inst/_058_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_010_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_243_  (.I0(\uart_tx_inst/data_reg[7] ),
    .I1(net26),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_059_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_244_  (.I0(\uart_tx_inst/data_reg[6] ),
    .I1(\uart_tx_inst/_059_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_011_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_245_  (.I0(\uart_tx_inst/data_reg[8] ),
    .I1(net27),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_060_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_246_  (.I0(\uart_tx_inst/data_reg[7] ),
    .I1(\uart_tx_inst/_060_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_012_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_247_  (.I0(\uart_tx_inst/data_reg[8] ),
    .I1(\uart_tx_inst/_036_ ),
    .S(\uart_tx_inst/_052_ ),
    .Z(\uart_tx_inst/_013_ ));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input3 (.I(prescale[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_249_  (.A1(\uart_tx_inst/_203_ [0]),
    .A2(\uart_tx_inst/_035_ ),
    .ZN(\uart_tx_inst/_062_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 \uart_tx_inst/_250_  (.A1(\uart_tx_inst/prescale_reg[10] ),
    .A2(\uart_tx_inst/_042_ ),
    .ZN(\uart_tx_inst/_063_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 \uart_tx_inst/_251_  (.A1(\uart_tx_inst/_044_ ),
    .A2(\uart_tx_inst/_045_ ),
    .ZN(\uart_tx_inst/_064_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 \uart_tx_inst/_252_  (.A1(\uart_tx_inst/prescale_reg[3] ),
    .A2(\uart_tx_inst/prescale_reg[2] ),
    .A3(\uart_tx_inst/prescale_reg[5] ),
    .A4(\uart_tx_inst/prescale_reg[4] ),
    .ZN(\uart_tx_inst/_065_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 \uart_tx_inst/_253_  (.A1(\uart_tx_inst/_195_ [0]),
    .A2(\uart_tx_inst/_065_ ),
    .Z(\uart_tx_inst/_066_ ));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 \uart_tx_inst/_254_  (.A1(\uart_tx_inst/_063_ ),
    .A2(\uart_tx_inst/_064_ ),
    .A3(\uart_tx_inst/_051_ ),
    .A4(\uart_tx_inst/_066_ ),
    .Z(\uart_tx_inst/_067_ ));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(prescale[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_256_  (.A1(\uart_tx_inst/_062_ ),
    .A2(\uart_tx_inst/_067_ ),
    .Z(\uart_tx_inst/_069_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 \uart_tx_inst/_257_  (.A1(\uart_tx_inst/_047_ ),
    .A2(\uart_tx_inst/_036_ ),
    .ZN(\uart_tx_inst/_070_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_258_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_070_ ),
    .ZN(\uart_tx_inst/_071_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_259_  (.I0(\uart_tx_inst/_069_ ),
    .I1(\uart_tx_inst/_071_ ),
    .S(\uart_tx_inst/_201_ [0]),
    .Z(\uart_tx_inst/_072_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_260_  (.A1(net18),
    .A2(\uart_tx_inst/_072_ ),
    .ZN(\uart_tx_inst/_000_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_261_  (.A1(\uart_tx_inst/bit_cnt[1] ),
    .A2(\uart_tx_inst/_071_ ),
    .ZN(\uart_tx_inst/_073_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 \uart_tx_inst/_262_  (.A1(\uart_tx_inst/_063_ ),
    .A2(\uart_tx_inst/_064_ ),
    .A3(\uart_tx_inst/_051_ ),
    .A4(\uart_tx_inst/_066_ ),
    .ZN(\uart_tx_inst/_074_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_263_  (.A1(\uart_tx_inst/_204_ [0]),
    .A2(\uart_tx_inst/_036_ ),
    .A3(\uart_tx_inst/_074_ ),
    .Z(\uart_tx_inst/_075_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 \uart_tx_inst/_264_  (.A1(\uart_tx_inst/_073_ ),
    .A2(\uart_tx_inst/_075_ ),
    .B(net18),
    .ZN(\uart_tx_inst/_001_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_265_  (.I(\uart_tx_inst/bit_cnt[2] ),
    .ZN(\uart_tx_inst/_076_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_266_  (.A1(\uart_tx_inst/bit_cnt[3] ),
    .A2(\uart_tx_inst/_076_ ),
    .Z(\uart_tx_inst/_077_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_267_  (.A1(\uart_tx_inst/_203_ [0]),
    .A2(\uart_tx_inst/_067_ ),
    .Z(\uart_tx_inst/_078_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_268_  (.I0(\uart_tx_inst/bit_cnt[2] ),
    .I1(\uart_tx_inst/_077_ ),
    .S(\uart_tx_inst/_078_ ),
    .Z(\uart_tx_inst/_079_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_269_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_079_ ),
    .Z(\uart_tx_inst/_002_ ));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 \uart_tx_inst/_270_  (.A1(\uart_tx_inst/_076_ ),
    .A2(\uart_tx_inst/_201_ [0]),
    .A3(\uart_tx_inst/_202_ [0]),
    .A4(\uart_tx_inst/_067_ ),
    .Z(\uart_tx_inst/_080_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 \uart_tx_inst/_271_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_070_ ),
    .Z(\uart_tx_inst/_081_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 \uart_tx_inst/_272_  (.A1(\uart_tx_inst/bit_cnt[2] ),
    .A2(\uart_tx_inst/bit_cnt[0] ),
    .A3(\uart_tx_inst/bit_cnt[1] ),
    .B(\uart_tx_inst/_062_ ),
    .ZN(\uart_tx_inst/_082_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 \uart_tx_inst/_273_  (.A1(\uart_tx_inst/_081_ ),
    .A2(\uart_tx_inst/_082_ ),
    .B(\uart_tx_inst/bit_cnt[3] ),
    .ZN(\uart_tx_inst/_083_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_274_  (.A1(\uart_tx_inst/bit_cnt[3] ),
    .A2(\uart_tx_inst/_080_ ),
    .B(\uart_tx_inst/_083_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_003_ ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 \uart_tx_inst/_275_  (.A1(\uart_tx_inst/_046_ ),
    .A2(\uart_tx_inst/_051_ ),
    .A3(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_084_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_276_  (.I0(net42),
    .I1(net28),
    .S(\uart_tx_inst/_084_ ),
    .Z(\uart_tx_inst/_085_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_277_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_085_ ),
    .Z(\uart_tx_inst/_004_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_278_  (.A1(\uart_tx_inst/prescale_reg[0] ),
    .A2(\uart_tx_inst/_074_ ),
    .ZN(\uart_tx_inst/_086_ ));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(m_axis_tready),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 \uart_tx_inst/_280_  (.A1(\uart_tx_inst/_035_ ),
    .A2(\uart_tx_inst/_049_ ),
    .Z(\uart_tx_inst/_088_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 \uart_tx_inst/_281_  (.A1(\uart_tx_inst/_193_ [0]),
    .A2(\uart_tx_inst/_070_ ),
    .B(\uart_tx_inst/_067_ ),
    .C(\uart_tx_inst/_088_ ),
    .ZN(\uart_tx_inst/_089_ ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 \uart_tx_inst/_282_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_086_ ),
    .A3(\uart_tx_inst/_089_ ),
    .Z(\uart_tx_inst/_014_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 \uart_tx_inst/_283_  (.A1(net9),
    .A2(net10),
    .A3(net2),
    .A4(net11),
    .Z(\uart_tx_inst/_090_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_284_  (.I(\uart_tx_inst/_205_ [0]),
    .ZN(\uart_tx_inst/_091_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 \uart_tx_inst/_285_  (.A1(\uart_tx_inst/bit_cnt[3] ),
    .A2(\uart_tx_inst/bit_cnt[2] ),
    .Z(\uart_tx_inst/_092_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_286_  (.A1(net12),
    .A2(net13),
    .ZN(\uart_tx_inst/_093_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 \uart_tx_inst/_287_  (.A1(\uart_tx_inst/_203_ [0]),
    .A2(\uart_tx_inst/_091_ ),
    .A3(\uart_tx_inst/_092_ ),
    .B(\uart_tx_inst/_093_ ),
    .ZN(\uart_tx_inst/_094_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_288_  (.A1(net14),
    .A2(\uart_tx_inst/_090_ ),
    .A3(\uart_tx_inst/_094_ ),
    .Z(\uart_tx_inst/_095_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_289_  (.A1(net15),
    .A2(\uart_tx_inst/_095_ ),
    .ZN(\uart_tx_inst/_096_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_290_  (.A1(\uart_tx_inst/_070_ ),
    .A2(\uart_tx_inst/_096_ ),
    .ZN(\uart_tx_inst/_097_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_291_  (.A1(\uart_tx_inst/_195_ [0]),
    .A2(\uart_tx_inst/_065_ ),
    .ZN(\uart_tx_inst/_098_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_292_  (.A1(\uart_tx_inst/_042_ ),
    .A2(\uart_tx_inst/_098_ ),
    .ZN(\uart_tx_inst/_099_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_293_  (.A1(\uart_tx_inst/prescale_reg[10] ),
    .A2(\uart_tx_inst/_099_ ),
    .ZN(\uart_tx_inst/_100_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_294_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_097_ ),
    .B(\uart_tx_inst/_100_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_015_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \uart_tx_inst/_295_  (.A1(net14),
    .A2(net15),
    .Z(\uart_tx_inst/_101_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_296_  (.I(\uart_tx_inst/_199_ [0]),
    .ZN(\uart_tx_inst/_102_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_297_  (.A1(net10),
    .A2(net11),
    .A3(\uart_tx_inst/_102_ ),
    .Z(\uart_tx_inst/_103_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 \uart_tx_inst/_298_  (.A1(\uart_tx_inst/_094_ ),
    .A2(\uart_tx_inst/_103_ ),
    .Z(\uart_tx_inst/_104_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \uart_tx_inst/_299_  (.A1(\uart_tx_inst/_101_ ),
    .A2(\uart_tx_inst/_104_ ),
    .Z(\uart_tx_inst/_105_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_300_  (.A1(net16),
    .A2(\uart_tx_inst/_105_ ),
    .Z(\uart_tx_inst/_106_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_301_  (.A1(\uart_tx_inst/prescale_reg[11] ),
    .A2(\uart_tx_inst/_043_ ),
    .Z(\uart_tx_inst/_107_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_302_  (.A1(\uart_tx_inst/_074_ ),
    .A2(\uart_tx_inst/_107_ ),
    .Z(\uart_tx_inst/_108_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_303_  (.A1(\uart_tx_inst/_047_ ),
    .A2(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_109_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_304_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_109_ ),
    .ZN(\uart_tx_inst/_110_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 \uart_tx_inst/_305_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_110_ ),
    .ZN(\uart_tx_inst/_111_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_306_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_106_ ),
    .B(\uart_tx_inst/_108_ ),
    .C(\uart_tx_inst/_111_ ),
    .ZN(\uart_tx_inst/_016_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_307_  (.A1(net16),
    .A2(\uart_tx_inst/_090_ ),
    .A3(\uart_tx_inst/_094_ ),
    .A4(\uart_tx_inst/_101_ ),
    .Z(\uart_tx_inst/_112_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_308_  (.A1(net17),
    .A2(\uart_tx_inst/_112_ ),
    .Z(\uart_tx_inst/_113_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_309_  (.A1(\uart_tx_inst/_063_ ),
    .A2(\uart_tx_inst/_066_ ),
    .ZN(\uart_tx_inst/_114_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_310_  (.A1(\uart_tx_inst/prescale_reg[11] ),
    .A2(\uart_tx_inst/_114_ ),
    .ZN(\uart_tx_inst/_115_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_311_  (.A1(\uart_tx_inst/prescale_reg[12] ),
    .A2(\uart_tx_inst/_115_ ),
    .ZN(\uart_tx_inst/_116_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_312_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_113_ ),
    .B(\uart_tx_inst/_116_ ),
    .C(\uart_tx_inst/_111_ ),
    .ZN(\uart_tx_inst/_017_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 \uart_tx_inst/_313_  (.A1(\uart_tx_inst/prescale_reg[13] ),
    .A2(\uart_tx_inst/prescale_reg[12] ),
    .A3(\uart_tx_inst/prescale_reg[11] ),
    .A4(\uart_tx_inst/_043_ ),
    .ZN(\uart_tx_inst/_117_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 \uart_tx_inst/_314_  (.A1(\uart_tx_inst/_064_ ),
    .A2(\uart_tx_inst/_051_ ),
    .A3(\uart_tx_inst/_066_ ),
    .ZN(\uart_tx_inst/_118_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_315_  (.A1(\uart_tx_inst/prescale_reg[12] ),
    .A2(\uart_tx_inst/prescale_reg[11] ),
    .A3(\uart_tx_inst/_043_ ),
    .Z(\uart_tx_inst/_119_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 \uart_tx_inst/_316_  (.A1(\uart_tx_inst/_117_ ),
    .A2(\uart_tx_inst/_118_ ),
    .B1(\uart_tx_inst/_119_ ),
    .B2(\uart_tx_inst/prescale_reg[13] ),
    .ZN(\uart_tx_inst/_120_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 \uart_tx_inst/_317_  (.A1(net14),
    .A2(net15),
    .A3(net16),
    .A4(net17),
    .Z(\uart_tx_inst/_121_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \uart_tx_inst/_318_  (.A1(\uart_tx_inst/_104_ ),
    .A2(\uart_tx_inst/_121_ ),
    .Z(\uart_tx_inst/_122_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_319_  (.A1(net3),
    .A2(\uart_tx_inst/_122_ ),
    .Z(\uart_tx_inst/_123_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_320_  (.A1(\uart_tx_inst/_063_ ),
    .A2(\uart_tx_inst/_064_ ),
    .Z(\uart_tx_inst/_124_ ));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 \uart_tx_inst/_321_  (.A1(\uart_tx_inst/_051_ ),
    .A2(\uart_tx_inst/_066_ ),
    .A3(\uart_tx_inst/_070_ ),
    .A4(\uart_tx_inst/_124_ ),
    .Z(\uart_tx_inst/_125_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_322_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_125_ ),
    .ZN(\uart_tx_inst/_126_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 \uart_tx_inst/_323_  (.A1(net18),
    .A2(\uart_tx_inst/_120_ ),
    .B1(\uart_tx_inst/_123_ ),
    .B2(\uart_tx_inst/_126_ ),
    .ZN(\uart_tx_inst/_018_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_324_  (.A1(\uart_tx_inst/prescale_reg[13] ),
    .A2(\uart_tx_inst/prescale_reg[12] ),
    .A3(\uart_tx_inst/prescale_reg[11] ),
    .A4(\uart_tx_inst/_114_ ),
    .Z(\uart_tx_inst/_127_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_325_  (.A1(\uart_tx_inst/prescale_reg[14] ),
    .A2(\uart_tx_inst/_127_ ),
    .ZN(\uart_tx_inst/_128_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \uart_tx_inst/_326_  (.A1(\uart_tx_inst/prescale_reg[17] ),
    .A2(\uart_tx_inst/prescale_reg[18] ),
    .Z(\uart_tx_inst/_129_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_327_  (.A1(net3),
    .A2(\uart_tx_inst/_090_ ),
    .A3(\uart_tx_inst/_094_ ),
    .A4(\uart_tx_inst/_121_ ),
    .Z(\uart_tx_inst/_130_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_328_  (.A1(net4),
    .A2(\uart_tx_inst/_130_ ),
    .ZN(\uart_tx_inst/_131_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_329_  (.A1(\uart_tx_inst/prescale_reg[14] ),
    .A2(\uart_tx_inst/_044_ ),
    .A3(\uart_tx_inst/_129_ ),
    .A4(\uart_tx_inst/_131_ ),
    .Z(\uart_tx_inst/_132_ ));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 \uart_tx_inst/_330_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_110_ ),
    .A3(\uart_tx_inst/_128_ ),
    .A4(\uart_tx_inst/_132_ ),
    .Z(\uart_tx_inst/_019_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_331_  (.A1(net3),
    .A2(net4),
    .A3(\uart_tx_inst/_104_ ),
    .A4(\uart_tx_inst/_121_ ),
    .Z(\uart_tx_inst/_133_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_332_  (.A1(net5),
    .A2(\uart_tx_inst/_133_ ),
    .Z(\uart_tx_inst/_134_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_333_  (.A1(\uart_tx_inst/_043_ ),
    .A2(\uart_tx_inst/_045_ ),
    .ZN(\uart_tx_inst/_135_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_334_  (.A1(\uart_tx_inst/prescale_reg[15] ),
    .A2(\uart_tx_inst/_135_ ),
    .ZN(\uart_tx_inst/_136_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_335_  (.A1(\uart_tx_inst/_074_ ),
    .A2(\uart_tx_inst/_136_ ),
    .Z(\uart_tx_inst/_137_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_336_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_134_ ),
    .B(\uart_tx_inst/_137_ ),
    .C(\uart_tx_inst/_111_ ),
    .ZN(\uart_tx_inst/_020_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 \uart_tx_inst/_337_  (.A1(\uart_tx_inst/prescale_reg[15] ),
    .A2(\uart_tx_inst/_045_ ),
    .A3(\uart_tx_inst/_114_ ),
    .ZN(\uart_tx_inst/_138_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_338_  (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(\uart_tx_inst/_121_ ),
    .Z(\uart_tx_inst/_139_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_339_  (.A1(\uart_tx_inst/_090_ ),
    .A2(\uart_tx_inst/_094_ ),
    .A3(\uart_tx_inst/_139_ ),
    .Z(\uart_tx_inst/_140_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_340_  (.A1(net6),
    .A2(\uart_tx_inst/_140_ ),
    .ZN(\uart_tx_inst/_141_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 \uart_tx_inst/_341_  (.A1(\uart_tx_inst/_081_ ),
    .A2(\uart_tx_inst/_141_ ),
    .B1(\uart_tx_inst/_138_ ),
    .B2(\uart_tx_inst/_129_ ),
    .C(\uart_tx_inst/prescale_reg[16] ),
    .ZN(\uart_tx_inst/_142_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_342_  (.A1(\uart_tx_inst/prescale_reg[16] ),
    .A2(\uart_tx_inst/_138_ ),
    .B(\uart_tx_inst/_142_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_021_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 \uart_tx_inst/_343_  (.A1(\uart_tx_inst/prescale_reg[18] ),
    .A2(\uart_tx_inst/_098_ ),
    .B(\uart_tx_inst/_046_ ),
    .ZN(\uart_tx_inst/_143_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_344_  (.I0(\uart_tx_inst/_143_ ),
    .I1(\uart_tx_inst/_046_ ),
    .S(\uart_tx_inst/prescale_reg[17] ),
    .Z(\uart_tx_inst/_144_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_345_  (.A1(net6),
    .A2(\uart_tx_inst/_104_ ),
    .A3(\uart_tx_inst/_139_ ),
    .Z(\uart_tx_inst/_145_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_346_  (.A1(net7),
    .A2(\uart_tx_inst/_145_ ),
    .Z(\uart_tx_inst/_146_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 \uart_tx_inst/_347_  (.A1(net18),
    .A2(\uart_tx_inst/_144_ ),
    .B1(\uart_tx_inst/_146_ ),
    .B2(\uart_tx_inst/_126_ ),
    .ZN(\uart_tx_inst/_022_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_348_  (.A1(\uart_tx_inst/prescale_reg[17] ),
    .A2(\uart_tx_inst/_044_ ),
    .A3(\uart_tx_inst/_045_ ),
    .A4(\uart_tx_inst/_114_ ),
    .Z(\uart_tx_inst/_147_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 \uart_tx_inst/_349_  (.A1(\uart_tx_inst/prescale_reg[18] ),
    .A2(\uart_tx_inst/_039_ ),
    .A3(\uart_tx_inst/_147_ ),
    .ZN(\uart_tx_inst/_148_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_350_  (.A1(net6),
    .A2(net7),
    .A3(\uart_tx_inst/_140_ ),
    .Z(\uart_tx_inst/_149_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_351_  (.A1(net8),
    .A2(\uart_tx_inst/_149_ ),
    .Z(\uart_tx_inst/_150_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 \uart_tx_inst/_352_  (.A1(\uart_tx_inst/_126_ ),
    .A2(\uart_tx_inst/_148_ ),
    .B1(\uart_tx_inst/_150_ ),
    .B2(\uart_tx_inst/_067_ ),
    .ZN(\uart_tx_inst/_023_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 \uart_tx_inst/_353_  (.A1(\uart_tx_inst/_203_ [0]),
    .A2(\uart_tx_inst/_091_ ),
    .A3(\uart_tx_inst/_092_ ),
    .Z(\uart_tx_inst/_151_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 \uart_tx_inst/_354_  (.A1(\uart_tx_inst/prescale_reg[1] ),
    .A2(\uart_tx_inst/_070_ ),
    .B(\uart_tx_inst/_151_ ),
    .ZN(\uart_tx_inst/_152_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_355_  (.I0(\uart_tx_inst/_196_ [0]),
    .I1(\uart_tx_inst/_152_ ),
    .S(\uart_tx_inst/_067_ ),
    .Z(\uart_tx_inst/_153_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_356_  (.A1(net18),
    .A2(\uart_tx_inst/_153_ ),
    .ZN(\uart_tx_inst/_024_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_357_  (.A1(\uart_tx_inst/prescale_reg[2] ),
    .A2(\uart_tx_inst/_195_ [0]),
    .ZN(\uart_tx_inst/_154_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_358_  (.A1(\uart_tx_inst/_088_ ),
    .A2(\uart_tx_inst/_067_ ),
    .B(\uart_tx_inst/_154_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_025_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_359_  (.A1(\uart_tx_inst/prescale_reg[2] ),
    .A2(\uart_tx_inst/_040_ ),
    .A3(\uart_tx_inst/_067_ ),
    .Z(\uart_tx_inst/_155_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_360_  (.A1(\uart_tx_inst/prescale_reg[3] ),
    .A2(\uart_tx_inst/_155_ ),
    .Z(\uart_tx_inst/_156_ ));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 \uart_tx_inst/_361_  (.A1(\uart_tx_inst/_048_ ),
    .A2(\uart_tx_inst/_205_ [0]),
    .A3(\uart_tx_inst/_035_ ),
    .Z(\uart_tx_inst/_157_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_362_  (.A1(\uart_tx_inst/_197_ [0]),
    .A2(\uart_tx_inst/_157_ ),
    .ZN(\uart_tx_inst/_158_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_363_  (.A1(net18),
    .A2(\uart_tx_inst/_071_ ),
    .A3(\uart_tx_inst/_158_ ),
    .Z(\uart_tx_inst/_159_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 \uart_tx_inst/_364_  (.A1(net18),
    .A2(\uart_tx_inst/_156_ ),
    .B(\uart_tx_inst/_159_ ),
    .ZN(\uart_tx_inst/_026_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_365_  (.I(\uart_tx_inst/_195_ [0]),
    .ZN(\uart_tx_inst/_160_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 \uart_tx_inst/_366_  (.A1(\uart_tx_inst/prescale_reg[3] ),
    .A2(\uart_tx_inst/prescale_reg[2] ),
    .A3(\uart_tx_inst/_160_ ),
    .A4(\uart_tx_inst/_067_ ),
    .ZN(\uart_tx_inst/_161_ ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \uart_tx_inst/_367_  (.I(\uart_tx_inst/_200_ [0]),
    .ZN(\uart_tx_inst/_162_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_368_  (.I0(net9),
    .I1(\uart_tx_inst/_162_ ),
    .S(\uart_tx_inst/_151_ ),
    .Z(\uart_tx_inst/_163_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_369_  (.A1(\uart_tx_inst/_125_ ),
    .A2(\uart_tx_inst/_163_ ),
    .B(\uart_tx_inst/_161_ ),
    .C(\uart_tx_inst/prescale_reg[4] ),
    .ZN(\uart_tx_inst/_164_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_370_  (.A1(\uart_tx_inst/prescale_reg[4] ),
    .A2(\uart_tx_inst/_161_ ),
    .B(\uart_tx_inst/_164_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_027_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_371_  (.A1(\uart_tx_inst/prescale_reg[3] ),
    .A2(\uart_tx_inst/prescale_reg[2] ),
    .A3(\uart_tx_inst/prescale_reg[4] ),
    .A4(\uart_tx_inst/_040_ ),
    .Z(\uart_tx_inst/_165_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_372_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_165_ ),
    .ZN(\uart_tx_inst/_166_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_373_  (.A1(\uart_tx_inst/_199_ [0]),
    .A2(\uart_tx_inst/_151_ ),
    .ZN(\uart_tx_inst/_167_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_374_  (.A1(net10),
    .A2(\uart_tx_inst/_167_ ),
    .ZN(\uart_tx_inst/_168_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_375_  (.A1(\uart_tx_inst/_081_ ),
    .A2(\uart_tx_inst/_168_ ),
    .B(\uart_tx_inst/_166_ ),
    .C(\uart_tx_inst/prescale_reg[5] ),
    .ZN(\uart_tx_inst/_169_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_376_  (.A1(\uart_tx_inst/prescale_reg[5] ),
    .A2(\uart_tx_inst/_166_ ),
    .B(\uart_tx_inst/_169_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_028_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 \uart_tx_inst/_377_  (.A1(net9),
    .A2(net10),
    .A3(net2),
    .A4(\uart_tx_inst/_157_ ),
    .ZN(\uart_tx_inst/_170_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_378_  (.A1(net11),
    .A2(\uart_tx_inst/_170_ ),
    .Z(\uart_tx_inst/_171_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_379_  (.A1(\uart_tx_inst/_070_ ),
    .A2(\uart_tx_inst/_171_ ),
    .ZN(\uart_tx_inst/_172_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_380_  (.A1(\uart_tx_inst/prescale_reg[6] ),
    .A2(\uart_tx_inst/_066_ ),
    .ZN(\uart_tx_inst/_173_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_381_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_172_ ),
    .B(\uart_tx_inst/_173_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_029_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \uart_tx_inst/_382_  (.A1(\uart_tx_inst/_040_ ),
    .A2(\uart_tx_inst/_041_ ),
    .Z(\uart_tx_inst/_174_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 \uart_tx_inst/_383_  (.A1(\uart_tx_inst/prescale_reg[6] ),
    .A2(\uart_tx_inst/_174_ ),
    .A3(\uart_tx_inst/_067_ ),
    .ZN(\uart_tx_inst/_175_ ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \uart_tx_inst/_384_  (.A1(\uart_tx_inst/_157_ ),
    .A2(\uart_tx_inst/_103_ ),
    .Z(\uart_tx_inst/_176_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_385_  (.A1(net12),
    .A2(\uart_tx_inst/_176_ ),
    .ZN(\uart_tx_inst/_177_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_386_  (.A1(\uart_tx_inst/_125_ ),
    .A2(\uart_tx_inst/_177_ ),
    .B(\uart_tx_inst/_175_ ),
    .C(\uart_tx_inst/prescale_reg[7] ),
    .ZN(\uart_tx_inst/_178_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_387_  (.A1(\uart_tx_inst/prescale_reg[7] ),
    .A2(\uart_tx_inst/_175_ ),
    .B(\uart_tx_inst/_178_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_030_ ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \uart_tx_inst/_388_  (.A1(net12),
    .A2(\uart_tx_inst/_090_ ),
    .A3(\uart_tx_inst/_157_ ),
    .Z(\uart_tx_inst/_179_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_389_  (.A1(net13),
    .A2(\uart_tx_inst/_179_ ),
    .ZN(\uart_tx_inst/_180_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_390_  (.A1(\uart_tx_inst/_070_ ),
    .A2(\uart_tx_inst/_180_ ),
    .ZN(\uart_tx_inst/_181_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 \uart_tx_inst/_391_  (.A1(\uart_tx_inst/prescale_reg[7] ),
    .A2(\uart_tx_inst/prescale_reg[6] ),
    .A3(\uart_tx_inst/_098_ ),
    .ZN(\uart_tx_inst/_182_ ));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \uart_tx_inst/_392_  (.A1(\uart_tx_inst/prescale_reg[8] ),
    .A2(\uart_tx_inst/_182_ ),
    .ZN(\uart_tx_inst/_183_ ));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \uart_tx_inst/_393_  (.A1(\uart_tx_inst/_067_ ),
    .A2(\uart_tx_inst/_181_ ),
    .B(\uart_tx_inst/_183_ ),
    .C(net18),
    .ZN(\uart_tx_inst/_031_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_394_  (.A1(net14),
    .A2(\uart_tx_inst/_104_ ),
    .Z(\uart_tx_inst/_184_ ));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \uart_tx_inst/_395_  (.A1(\uart_tx_inst/prescale_reg[7] ),
    .A2(\uart_tx_inst/prescale_reg[6] ),
    .A3(\uart_tx_inst/prescale_reg[8] ),
    .A4(\uart_tx_inst/_174_ ),
    .Z(\uart_tx_inst/_185_ ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \uart_tx_inst/_396_  (.A1(\uart_tx_inst/prescale_reg[9] ),
    .A2(\uart_tx_inst/_185_ ),
    .Z(\uart_tx_inst/_186_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_397_  (.I0(\uart_tx_inst/_184_ ),
    .I1(\uart_tx_inst/_186_ ),
    .S(\uart_tx_inst/_074_ ),
    .Z(\uart_tx_inst/_187_ ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \uart_tx_inst/_398_  (.A1(\uart_tx_inst/_111_ ),
    .A2(\uart_tx_inst/_187_ ),
    .ZN(\uart_tx_inst/_032_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_399_  (.A1(net28),
    .A2(net41),
    .ZN(\uart_tx_inst/_188_ ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \uart_tx_inst/_400_  (.I0(net41),
    .I1(\uart_tx_inst/_188_ ),
    .S(\uart_tx_inst/_036_ ),
    .Z(\uart_tx_inst/_189_ ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 \uart_tx_inst/_401_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_067_ ),
    .A3(\uart_tx_inst/_189_ ),
    .Z(\uart_tx_inst/_033_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \uart_tx_inst/_402_  (.A1(net43),
    .A2(\uart_tx_inst/_071_ ),
    .ZN(\uart_tx_inst/_190_ ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \uart_tx_inst/_403_  (.A1(\uart_tx_inst/_205_ [0]),
    .A2(\uart_tx_inst/_035_ ),
    .Z(\uart_tx_inst/_191_ ));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 \uart_tx_inst/_404_  (.A1(\uart_tx_inst/data_reg[0] ),
    .A2(\uart_tx_inst/_191_ ),
    .B(\uart_tx_inst/_069_ ),
    .ZN(\uart_tx_inst/_192_ ));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 \uart_tx_inst/_405_  (.A1(\uart_tx_inst/_039_ ),
    .A2(\uart_tx_inst/_190_ ),
    .A3(\uart_tx_inst/_192_ ),
    .ZN(\uart_tx_inst/_034_ ));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 \uart_tx_inst/_406_  (.A(\uart_tx_inst/_193_ [0]),
    .B(\uart_tx_inst/_194_ [0]),
    .CO(\uart_tx_inst/_195_ [0]),
    .S(\uart_tx_inst/_196_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 \uart_tx_inst/_407_  (.A(\uart_tx_inst/_197_ [0]),
    .B(\uart_tx_inst/_198_ [0]),
    .CO(\uart_tx_inst/_199_ [0]),
    .S(\uart_tx_inst/_200_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 \uart_tx_inst/_408_  (.A(\uart_tx_inst/_201_ [0]),
    .B(\uart_tx_inst/_202_ [0]),
    .CO(\uart_tx_inst/_203_ [0]),
    .S(\uart_tx_inst/_204_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 \uart_tx_inst/_409_  (.A(\uart_tx_inst/bit_cnt[0] ),
    .B(\uart_tx_inst/_202_ [0]),
    .CO(\uart_tx_inst/_205_ [0]),
    .S(\uart_tx_inst/_206_ [0]));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/bit_cnt[0]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_000_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/bit_cnt[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/bit_cnt[1]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_001_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/bit_cnt[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/bit_cnt[2]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_002_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/bit_cnt[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/bit_cnt[3]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_003_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/bit_cnt[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/busy_reg$_SDFFE_PP0P_  (.D(\uart_tx_inst/_004_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[0]$_DFFE_PP_  (.D(\uart_tx_inst/_005_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[1]$_DFFE_PP_  (.D(\uart_tx_inst/_006_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[2]$_DFFE_PP_  (.D(\uart_tx_inst/_007_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[3]$_DFFE_PP_  (.D(\uart_tx_inst/_008_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[4]$_DFFE_PP_  (.D(\uart_tx_inst/_009_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[5]$_DFFE_PP_  (.D(\uart_tx_inst/_010_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[6]$_DFFE_PP_  (.D(\uart_tx_inst/_011_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[7]$_DFFE_PP_  (.D(\uart_tx_inst/_012_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/data_reg[8]$_DFFE_PP_  (.D(\uart_tx_inst/_013_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(\uart_tx_inst/data_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[0]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_014_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[10]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_015_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[11]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_016_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[12]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_017_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[13]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_018_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[14]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_019_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[15]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_020_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[16]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_021_ ),
    .CLK(clknet_2_3__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[17]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_022_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[18]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_023_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[1]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_024_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[2]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_025_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[3]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_026_ ),
    .CLK(clknet_2_0__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[4]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_027_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[5]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_028_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[6]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_029_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[7]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_030_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[8]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_031_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/prescale_reg[9]$_SDFFE_PP0P_  (.D(\uart_tx_inst/_032_ ),
    .CLK(clknet_2_1__leaf_clk_regs),
    .Q(\uart_tx_inst/prescale_reg[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/s_axis_tready_reg$_SDFFE_PP0P_  (.D(\uart_tx_inst/_033_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \uart_tx_inst/txd_reg$_SDFFE_PP1P_  (.D(\uart_tx_inst/_034_ ),
    .CLK(clknet_2_2__leaf_clk_regs),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_2_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_2_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_2_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_2_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_2_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_2_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_2_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_2_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_2_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_2_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_2_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_2_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_2_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_2_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_2_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_2_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_2_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_2_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_2_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_2_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_2_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_2_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_2_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_2_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_2_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_2_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_2_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_2_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_2_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_2_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_2_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_2_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_2_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_2_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_2_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_2_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_2_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_2_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_2_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_2_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_2_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_2_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_2_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_2_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_2_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_2_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_2_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_2_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_2_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_2_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_2_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_1_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_1_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_1_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_1_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_1_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_1_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_1_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_1_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_1_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_1_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_1_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_1_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_1_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_1_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_1_Left_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_1_Left_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_1_Left_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_1_Left_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_1_Left_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_1_Left_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_1_Left_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_1_Left_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_1_Left_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_1_Left_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_1_Left_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_1_Left_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_1_Left_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_1_Left_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_1_Left_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_1_Left_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_1_Left_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_1_Left_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_1_Left_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_1_Left_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_1_Left_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_1_Left_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_1_Left_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_1_Left_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_1_Left_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_1_Left_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_1_Left_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_1_Left_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_1_Left_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_1_Left_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_1_Left_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_1_Left_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_1_Left_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_1_Left_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_1_Left_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_1_Left_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_1_Left_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_2_Left_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_2_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_2_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_2_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_2_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_2_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_2_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_2_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_2_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_2_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_2_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_2_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_2_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_2_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_2_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_2_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_2_Left_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_2_Left_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_2_Left_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_2_Left_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_2_Left_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_2_Left_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_2_Left_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_2_Left_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_2_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_2_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_2_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_2_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_2_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_2_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_2_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_2_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_2_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_2_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_2_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_2_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_2_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_2_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_2_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_2_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_2_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_2_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_2_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_2_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_2_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_2_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_2_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_2_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_2_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_2_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_2_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_1_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_1_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_1_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_1_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_1_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_1_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_1_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_1_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_1_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_1_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_1_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_1_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_1_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_1_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_1_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_1_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_1_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_1_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_1_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_1_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_1_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_1_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_1_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_1_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_1_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_1_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_1_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_1_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_1_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_1_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_1_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_1_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_1_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_1_Right_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_1_Right_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_1_Right_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_1_Right_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_1_Right_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_1_Right_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_1_Right_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_1_Right_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_1_Right_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_1_Right_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_1_Right_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_1_Right_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_1_Right_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_1_Right_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_1_Right_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_1_Right_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_1_Right_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_1_Right_263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1_268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1_269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1_270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1_271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1_272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1_273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1_274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1_275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1_276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1_277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1_278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1_279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1_280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1_281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1_282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1_283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1_284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1_285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1_286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1_287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1_288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1_289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1_290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1_291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1_292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_354 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input6 (.I(prescale[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(prescale[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(prescale[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(prescale[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input10 (.I(prescale[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input11 (.I(prescale[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(prescale[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input13 (.I(prescale[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(prescale[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input15 (.I(prescale[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input16 (.I(prescale[8]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input17 (.I(prescale[9]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 input18 (.I(rst),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(rxd),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(s_axis_tdata[0]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input21 (.I(s_axis_tdata[1]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(s_axis_tdata[2]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input23 (.I(s_axis_tdata[3]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input24 (.I(s_axis_tdata[4]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input25 (.I(s_axis_tdata[5]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input26 (.I(s_axis_tdata[6]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input27 (.I(s_axis_tdata[7]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input28 (.I(s_axis_tvalid),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output29 (.I(net29),
    .Z(m_axis_tdata[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output30 (.I(net30),
    .Z(m_axis_tdata[1]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output31 (.I(net31),
    .Z(m_axis_tdata[2]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output32 (.I(net32),
    .Z(m_axis_tdata[3]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output33 (.I(net33),
    .Z(m_axis_tdata[4]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output34 (.I(net34),
    .Z(m_axis_tdata[5]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output35 (.I(net35),
    .Z(m_axis_tdata[6]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output36 (.I(net36),
    .Z(m_axis_tdata[7]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output37 (.I(net37),
    .Z(m_axis_tvalid));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output38 (.I(net38),
    .Z(rx_busy));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output39 (.I(net39),
    .Z(rx_frame_error));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output40 (.I(net40),
    .Z(rx_overrun_error));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output41 (.I(net41),
    .Z(s_axis_tready));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output42 (.I(net42),
    .Z(tx_busy));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output43 (.I(net43),
    .Z(txd));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_regs_0_clk (.I(clk),
    .Z(delaynet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk_regs (.I(clk_regs),
    .Z(clknet_0_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_2_0__f_clk_regs (.I(clknet_0_clk_regs),
    .Z(clknet_2_0__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_2_1__f_clk_regs (.I(clknet_0_clk_regs),
    .Z(clknet_2_1__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_2_2__f_clk_regs (.I(clknet_0_clk_regs),
    .Z(clknet_2_2__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_2_3__f_clk_regs (.I(clknet_0_clk_regs),
    .Z(clknet_2_3__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_2_0__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_2_1__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload2 (.I(clknet_2_3__leaf_clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 delaybuf_0_clk (.I(delaynet_0_clk),
    .Z(clk_regs));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_11 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_714 ();
endmodule
