module smart_fifo (almost_empty,
    almost_full,
    clear_errors,
    clk,
    empty,
    error_detected,
    full,
    overflow_detected,
    rd_en,
    rd_valid,
    rst_n,
    underflow_detected,
    wr_en,
    wr_ready,
    data_count,
    error_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clear_errors;
 input clk;
 output empty;
 output error_detected;
 output full;
 output overflow_detected;
 input rd_en;
 output rd_valid;
 input rst_n;
 output underflow_detected;
 input wr_en;
 output wr_ready;
 output [4:0] data_count;
 output [15:0] error_count;
 output [31:0] rd_data;
 input [31:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire \last_valid_data[0] ;
 wire \last_valid_data[10] ;
 wire \last_valid_data[11] ;
 wire \last_valid_data[12] ;
 wire \last_valid_data[13] ;
 wire \last_valid_data[14] ;
 wire \last_valid_data[15] ;
 wire \last_valid_data[16] ;
 wire \last_valid_data[17] ;
 wire \last_valid_data[18] ;
 wire \last_valid_data[19] ;
 wire \last_valid_data[1] ;
 wire \last_valid_data[20] ;
 wire \last_valid_data[21] ;
 wire \last_valid_data[22] ;
 wire \last_valid_data[23] ;
 wire \last_valid_data[24] ;
 wire \last_valid_data[25] ;
 wire \last_valid_data[26] ;
 wire \last_valid_data[27] ;
 wire \last_valid_data[28] ;
 wire \last_valid_data[29] ;
 wire \last_valid_data[2] ;
 wire \last_valid_data[30] ;
 wire \last_valid_data[31] ;
 wire \last_valid_data[3] ;
 wire \last_valid_data[4] ;
 wire \last_valid_data[5] ;
 wire \last_valid_data[6] ;
 wire \last_valid_data[7] ;
 wire \last_valid_data[8] ;
 wire \last_valid_data[9] ;
 wire last_valid_data_available;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;

 INV_X1 _2322_ (.A(_2321_),
    .ZN(net4));
 BUF_X4 _2323_ (.A(_2309_),
    .Z(_0583_));
 XOR2_X2 _2324_ (.A(_0583_),
    .B(_2301_),
    .Z(net6));
 AOI21_X1 _2325_ (.A(_2308_),
    .B1(_2305_),
    .B2(_0583_),
    .ZN(_0584_));
 NAND2_X1 _2326_ (.A1(_0583_),
    .A2(_2306_),
    .ZN(_0585_));
 OAI21_X2 _2327_ (.A(_0584_),
    .B1(_0585_),
    .B2(net64),
    .ZN(_0586_));
 XNOR2_X1 _2328_ (.A(_2304_),
    .B(_0586_),
    .ZN(_0587_));
 INV_X1 _2329_ (.A(_0587_),
    .ZN(net7));
 INV_X1 _2330_ (.A(_2303_),
    .ZN(_0588_));
 AOI21_X1 _2331_ (.A(_2308_),
    .B1(_2301_),
    .B2(_0583_),
    .ZN(_0589_));
 INV_X1 _2332_ (.A(_2304_),
    .ZN(_0590_));
 OAI21_X1 _2333_ (.A(_0588_),
    .B1(_0589_),
    .B2(_0590_),
    .ZN(_0591_));
 XOR2_X2 _2334_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Z(_0592_));
 XOR2_X2 _2335_ (.A(_0591_),
    .B(_0592_),
    .Z(_0593_));
 INV_X1 _2336_ (.A(_0593_),
    .ZN(_0594_));
 BUF_X4 _2337_ (.A(_0594_),
    .Z(_0595_));
 BUF_X4 _2338_ (.A(_0595_),
    .Z(_0596_));
 CLKBUF_X3 _2339_ (.A(_0596_),
    .Z(net8));
 BUF_X4 _2340_ (.A(_0595_),
    .Z(_0597_));
 BUF_X1 _2341_ (.A(net5),
    .Z(_0598_));
 NOR4_X1 _2342_ (.A1(_2304_),
    .A2(net4),
    .A3(_0598_),
    .A4(net6),
    .ZN(_0599_));
 NOR4_X1 _2343_ (.A1(_0590_),
    .A2(net4),
    .A3(_0598_),
    .A4(net6),
    .ZN(_0600_));
 MUX2_X2 _2344_ (.A(_0599_),
    .B(_0600_),
    .S(_0586_),
    .Z(_0601_));
 CLKBUF_X3 _2345_ (.A(_0601_),
    .Z(_0602_));
 NAND2_X1 _2346_ (.A1(_0597_),
    .A2(_0602_),
    .ZN(net63));
 INV_X1 _2347_ (.A(net63),
    .ZN(net27));
 OR4_X2 _2348_ (.A1(_2304_),
    .A2(net6),
    .A3(_0598_),
    .A4(net4),
    .ZN(_0603_));
 OR4_X2 _2349_ (.A1(net6),
    .A2(net4),
    .A3(_0598_),
    .A4(_0590_),
    .ZN(_0604_));
 MUX2_X2 _2350_ (.A(_0603_),
    .B(_0604_),
    .S(_0586_),
    .Z(_0605_));
 NOR2_X4 _2351_ (.A1(_0594_),
    .A2(_0605_),
    .ZN(net9));
 INV_X8 _2352_ (.A(net9),
    .ZN(_0606_));
 BUF_X32 _2353_ (.A(_0606_),
    .Z(_0607_));
 BUF_X4 _2354_ (.A(_0607_),
    .Z(net61));
 CLKBUF_X3 _2355_ (.A(rd_en),
    .Z(_0608_));
 NAND3_X2 _2356_ (.A1(_0608_),
    .A2(_0593_),
    .A3(_0601_),
    .ZN(_0609_));
 INV_X1 _2357_ (.A(_0609_),
    .ZN(net62));
 INV_X1 _2358_ (.A(_2320_),
    .ZN(_2300_));
 CLKBUF_X2 _2359_ (.A(wr_data[0]),
    .Z(_0610_));
 BUF_X2 _2360_ (.A(_0610_),
    .Z(_0611_));
 BUF_X2 _2361_ (.A(_2313_),
    .Z(_0612_));
 BUF_X1 _2362_ (.A(wr_en),
    .Z(_0613_));
 INV_X2 _2363_ (.A(_0613_),
    .ZN(_0614_));
 BUF_X2 _2364_ (.A(\wr_ptr[3] ),
    .Z(_0615_));
 CLKBUF_X2 _2365_ (.A(\wr_ptr[2] ),
    .Z(_0616_));
 NOR3_X2 _2366_ (.A1(_0614_),
    .A2(_0615_),
    .A3(_0616_),
    .ZN(_0617_));
 AND2_X1 _2367_ (.A1(_0612_),
    .A2(_0617_),
    .ZN(_0618_));
 CLKBUF_X3 _2368_ (.A(_0618_),
    .Z(_0619_));
 BUF_X4 _2369_ (.A(_0619_),
    .Z(_0620_));
 MUX2_X1 _2370_ (.A(\mem[0][0] ),
    .B(_0611_),
    .S(_0620_),
    .Z(_0064_));
 BUF_X1 _2371_ (.A(wr_data[10]),
    .Z(_0621_));
 CLKBUF_X2 _2372_ (.A(_0621_),
    .Z(_0622_));
 MUX2_X1 _2373_ (.A(\mem[0][10] ),
    .B(_0622_),
    .S(_0620_),
    .Z(_0065_));
 CLKBUF_X2 _2374_ (.A(wr_data[11]),
    .Z(_0623_));
 BUF_X2 _2375_ (.A(_0623_),
    .Z(_0624_));
 MUX2_X1 _2376_ (.A(\mem[0][11] ),
    .B(_0624_),
    .S(_0620_),
    .Z(_0066_));
 CLKBUF_X2 _2377_ (.A(wr_data[12]),
    .Z(_0625_));
 BUF_X2 _2378_ (.A(_0625_),
    .Z(_0626_));
 MUX2_X1 _2379_ (.A(\mem[0][12] ),
    .B(_0626_),
    .S(_0620_),
    .Z(_0067_));
 BUF_X1 _2380_ (.A(wr_data[13]),
    .Z(_0627_));
 BUF_X2 _2381_ (.A(_0627_),
    .Z(_0628_));
 MUX2_X1 _2382_ (.A(\mem[0][13] ),
    .B(_0628_),
    .S(_0620_),
    .Z(_0068_));
 CLKBUF_X2 _2383_ (.A(wr_data[14]),
    .Z(_0629_));
 BUF_X2 _2384_ (.A(_0629_),
    .Z(_0630_));
 MUX2_X1 _2385_ (.A(\mem[0][14] ),
    .B(_0630_),
    .S(_0620_),
    .Z(_0069_));
 CLKBUF_X2 _2386_ (.A(wr_data[15]),
    .Z(_0631_));
 BUF_X2 _2387_ (.A(_0631_),
    .Z(_0632_));
 MUX2_X1 _2388_ (.A(\mem[0][15] ),
    .B(_0632_),
    .S(_0620_),
    .Z(_0070_));
 CLKBUF_X2 _2389_ (.A(wr_data[16]),
    .Z(_0633_));
 CLKBUF_X2 _2390_ (.A(_0633_),
    .Z(_0634_));
 MUX2_X1 _2391_ (.A(\mem[0][16] ),
    .B(_0634_),
    .S(_0620_),
    .Z(_0071_));
 BUF_X2 _2392_ (.A(wr_data[17]),
    .Z(_0635_));
 BUF_X2 _2393_ (.A(_0635_),
    .Z(_0636_));
 MUX2_X1 _2394_ (.A(\mem[0][17] ),
    .B(_0636_),
    .S(_0620_),
    .Z(_0072_));
 BUF_X2 _2395_ (.A(wr_data[18]),
    .Z(_0637_));
 CLKBUF_X2 _2396_ (.A(_0637_),
    .Z(_0638_));
 MUX2_X1 _2397_ (.A(\mem[0][18] ),
    .B(_0638_),
    .S(_0620_),
    .Z(_0073_));
 BUF_X2 _2398_ (.A(wr_data[19]),
    .Z(_0639_));
 CLKBUF_X2 _2399_ (.A(_0639_),
    .Z(_0640_));
 BUF_X4 _2400_ (.A(_0619_),
    .Z(_0641_));
 MUX2_X1 _2401_ (.A(\mem[0][19] ),
    .B(_0640_),
    .S(_0641_),
    .Z(_0074_));
 BUF_X1 _2402_ (.A(wr_data[1]),
    .Z(_0642_));
 BUF_X2 _2403_ (.A(_0642_),
    .Z(_0643_));
 MUX2_X1 _2404_ (.A(\mem[0][1] ),
    .B(_0643_),
    .S(_0641_),
    .Z(_0075_));
 BUF_X1 _2405_ (.A(wr_data[20]),
    .Z(_0644_));
 BUF_X2 _2406_ (.A(_0644_),
    .Z(_0645_));
 MUX2_X1 _2407_ (.A(\mem[0][20] ),
    .B(_0645_),
    .S(_0641_),
    .Z(_0076_));
 BUF_X1 _2408_ (.A(wr_data[21]),
    .Z(_0646_));
 BUF_X2 _2409_ (.A(_0646_),
    .Z(_0647_));
 MUX2_X1 _2410_ (.A(\mem[0][21] ),
    .B(_0647_),
    .S(_0641_),
    .Z(_0077_));
 BUF_X1 _2411_ (.A(wr_data[22]),
    .Z(_0648_));
 BUF_X2 _2412_ (.A(_0648_),
    .Z(_0649_));
 MUX2_X1 _2413_ (.A(\mem[0][22] ),
    .B(_0649_),
    .S(_0641_),
    .Z(_0078_));
 BUF_X1 _2414_ (.A(wr_data[23]),
    .Z(_0650_));
 CLKBUF_X2 _2415_ (.A(_0650_),
    .Z(_0651_));
 MUX2_X1 _2416_ (.A(\mem[0][23] ),
    .B(_0651_),
    .S(_0641_),
    .Z(_0079_));
 BUF_X1 _2417_ (.A(wr_data[24]),
    .Z(_0652_));
 BUF_X2 _2418_ (.A(_0652_),
    .Z(_0653_));
 MUX2_X1 _2419_ (.A(\mem[0][24] ),
    .B(_0653_),
    .S(_0641_),
    .Z(_0080_));
 BUF_X1 _2420_ (.A(wr_data[25]),
    .Z(_0654_));
 BUF_X2 _2421_ (.A(_0654_),
    .Z(_0655_));
 MUX2_X1 _2422_ (.A(\mem[0][25] ),
    .B(_0655_),
    .S(_0641_),
    .Z(_0081_));
 BUF_X1 _2423_ (.A(wr_data[26]),
    .Z(_0656_));
 BUF_X2 _2424_ (.A(_0656_),
    .Z(_0657_));
 MUX2_X1 _2425_ (.A(\mem[0][26] ),
    .B(_0657_),
    .S(_0641_),
    .Z(_0082_));
 CLKBUF_X2 _2426_ (.A(wr_data[27]),
    .Z(_0658_));
 BUF_X2 _2427_ (.A(_0658_),
    .Z(_0659_));
 MUX2_X1 _2428_ (.A(\mem[0][27] ),
    .B(_0659_),
    .S(_0641_),
    .Z(_0083_));
 CLKBUF_X2 _2429_ (.A(wr_data[28]),
    .Z(_0660_));
 BUF_X2 _2430_ (.A(_0660_),
    .Z(_0661_));
 BUF_X4 _2431_ (.A(_0619_),
    .Z(_0662_));
 MUX2_X1 _2432_ (.A(\mem[0][28] ),
    .B(_0661_),
    .S(_0662_),
    .Z(_0084_));
 BUF_X2 _2433_ (.A(wr_data[29]),
    .Z(_0663_));
 BUF_X2 _2434_ (.A(_0663_),
    .Z(_0664_));
 MUX2_X1 _2435_ (.A(\mem[0][29] ),
    .B(_0664_),
    .S(_0662_),
    .Z(_0085_));
 CLKBUF_X2 _2436_ (.A(wr_data[2]),
    .Z(_0665_));
 BUF_X2 _2437_ (.A(_0665_),
    .Z(_0666_));
 MUX2_X1 _2438_ (.A(\mem[0][2] ),
    .B(_0666_),
    .S(_0662_),
    .Z(_0086_));
 CLKBUF_X2 _2439_ (.A(wr_data[30]),
    .Z(_0667_));
 BUF_X2 _2440_ (.A(_0667_),
    .Z(_0668_));
 MUX2_X1 _2441_ (.A(\mem[0][30] ),
    .B(_0668_),
    .S(_0662_),
    .Z(_0087_));
 CLKBUF_X2 _2442_ (.A(wr_data[31]),
    .Z(_0669_));
 BUF_X2 _2443_ (.A(_0669_),
    .Z(_0670_));
 MUX2_X1 _2444_ (.A(\mem[0][31] ),
    .B(_0670_),
    .S(_0662_),
    .Z(_0088_));
 BUF_X1 _2445_ (.A(wr_data[3]),
    .Z(_0671_));
 BUF_X2 _2446_ (.A(_0671_),
    .Z(_0672_));
 MUX2_X1 _2447_ (.A(\mem[0][3] ),
    .B(_0672_),
    .S(_0662_),
    .Z(_0089_));
 CLKBUF_X2 _2448_ (.A(wr_data[4]),
    .Z(_0673_));
 BUF_X2 _2449_ (.A(_0673_),
    .Z(_0674_));
 MUX2_X1 _2450_ (.A(\mem[0][4] ),
    .B(_0674_),
    .S(_0662_),
    .Z(_0090_));
 CLKBUF_X2 _2451_ (.A(wr_data[5]),
    .Z(_0675_));
 BUF_X2 _2452_ (.A(_0675_),
    .Z(_0676_));
 MUX2_X1 _2453_ (.A(\mem[0][5] ),
    .B(_0676_),
    .S(_0662_),
    .Z(_0091_));
 CLKBUF_X2 _2454_ (.A(wr_data[6]),
    .Z(_0677_));
 BUF_X2 _2455_ (.A(_0677_),
    .Z(_0678_));
 MUX2_X1 _2456_ (.A(\mem[0][6] ),
    .B(_0678_),
    .S(_0662_),
    .Z(_0092_));
 CLKBUF_X2 _2457_ (.A(wr_data[7]),
    .Z(_0679_));
 BUF_X2 _2458_ (.A(_0679_),
    .Z(_0680_));
 MUX2_X1 _2459_ (.A(\mem[0][7] ),
    .B(_0680_),
    .S(_0662_),
    .Z(_0093_));
 CLKBUF_X2 _2460_ (.A(wr_data[8]),
    .Z(_0681_));
 BUF_X2 _2461_ (.A(_0681_),
    .Z(_0682_));
 MUX2_X1 _2462_ (.A(\mem[0][8] ),
    .B(_0682_),
    .S(_0619_),
    .Z(_0094_));
 CLKBUF_X2 _2463_ (.A(wr_data[9]),
    .Z(_0683_));
 BUF_X2 _2464_ (.A(_0683_),
    .Z(_0684_));
 MUX2_X1 _2465_ (.A(\mem[0][9] ),
    .B(_0684_),
    .S(_0619_),
    .Z(_0095_));
 BUF_X1 _2466_ (.A(_2314_),
    .Z(_0685_));
 INV_X1 _2467_ (.A(_0616_),
    .ZN(_0686_));
 AND3_X1 _2468_ (.A1(_0613_),
    .A2(_0615_),
    .A3(_0686_),
    .ZN(_0687_));
 CLKBUF_X3 _2469_ (.A(_0687_),
    .Z(_0688_));
 NAND2_X2 _2470_ (.A1(_0685_),
    .A2(_0688_),
    .ZN(_0689_));
 BUF_X4 _2471_ (.A(_0689_),
    .Z(_0690_));
 MUX2_X1 _2472_ (.A(_0611_),
    .B(\mem[10][0] ),
    .S(_0690_),
    .Z(_0096_));
 MUX2_X1 _2473_ (.A(_0622_),
    .B(\mem[10][10] ),
    .S(_0690_),
    .Z(_0097_));
 MUX2_X1 _2474_ (.A(_0624_),
    .B(\mem[10][11] ),
    .S(_0690_),
    .Z(_0098_));
 MUX2_X1 _2475_ (.A(_0626_),
    .B(\mem[10][12] ),
    .S(_0690_),
    .Z(_0099_));
 MUX2_X1 _2476_ (.A(_0628_),
    .B(\mem[10][13] ),
    .S(_0690_),
    .Z(_0100_));
 MUX2_X1 _2477_ (.A(_0630_),
    .B(\mem[10][14] ),
    .S(_0690_),
    .Z(_0101_));
 MUX2_X1 _2478_ (.A(_0632_),
    .B(\mem[10][15] ),
    .S(_0690_),
    .Z(_0102_));
 MUX2_X1 _2479_ (.A(_0634_),
    .B(\mem[10][16] ),
    .S(_0690_),
    .Z(_0103_));
 MUX2_X1 _2480_ (.A(_0636_),
    .B(\mem[10][17] ),
    .S(_0690_),
    .Z(_0104_));
 MUX2_X1 _2481_ (.A(_0638_),
    .B(\mem[10][18] ),
    .S(_0690_),
    .Z(_0105_));
 BUF_X4 _2482_ (.A(_0689_),
    .Z(_0691_));
 MUX2_X1 _2483_ (.A(_0640_),
    .B(\mem[10][19] ),
    .S(_0691_),
    .Z(_0106_));
 MUX2_X1 _2484_ (.A(_0643_),
    .B(\mem[10][1] ),
    .S(_0691_),
    .Z(_0107_));
 MUX2_X1 _2485_ (.A(_0645_),
    .B(\mem[10][20] ),
    .S(_0691_),
    .Z(_0108_));
 MUX2_X1 _2486_ (.A(_0647_),
    .B(\mem[10][21] ),
    .S(_0691_),
    .Z(_0109_));
 MUX2_X1 _2487_ (.A(_0649_),
    .B(\mem[10][22] ),
    .S(_0691_),
    .Z(_0110_));
 MUX2_X1 _2488_ (.A(_0651_),
    .B(\mem[10][23] ),
    .S(_0691_),
    .Z(_0111_));
 MUX2_X1 _2489_ (.A(_0653_),
    .B(\mem[10][24] ),
    .S(_0691_),
    .Z(_0112_));
 MUX2_X1 _2490_ (.A(_0655_),
    .B(\mem[10][25] ),
    .S(_0691_),
    .Z(_0113_));
 MUX2_X1 _2491_ (.A(_0657_),
    .B(\mem[10][26] ),
    .S(_0691_),
    .Z(_0114_));
 MUX2_X1 _2492_ (.A(_0659_),
    .B(\mem[10][27] ),
    .S(_0691_),
    .Z(_0115_));
 CLKBUF_X3 _2493_ (.A(_0689_),
    .Z(_0692_));
 MUX2_X1 _2494_ (.A(_0661_),
    .B(\mem[10][28] ),
    .S(_0692_),
    .Z(_0116_));
 MUX2_X1 _2495_ (.A(_0664_),
    .B(\mem[10][29] ),
    .S(_0692_),
    .Z(_0117_));
 MUX2_X1 _2496_ (.A(_0666_),
    .B(\mem[10][2] ),
    .S(_0692_),
    .Z(_0118_));
 MUX2_X1 _2497_ (.A(_0668_),
    .B(\mem[10][30] ),
    .S(_0692_),
    .Z(_0119_));
 MUX2_X1 _2498_ (.A(_0670_),
    .B(\mem[10][31] ),
    .S(_0692_),
    .Z(_0120_));
 MUX2_X1 _2499_ (.A(_0672_),
    .B(\mem[10][3] ),
    .S(_0692_),
    .Z(_0121_));
 MUX2_X1 _2500_ (.A(_0674_),
    .B(\mem[10][4] ),
    .S(_0692_),
    .Z(_0122_));
 MUX2_X1 _2501_ (.A(_0676_),
    .B(\mem[10][5] ),
    .S(_0692_),
    .Z(_0123_));
 MUX2_X1 _2502_ (.A(_0678_),
    .B(\mem[10][6] ),
    .S(_0692_),
    .Z(_0124_));
 MUX2_X1 _2503_ (.A(_0680_),
    .B(\mem[10][7] ),
    .S(_0692_),
    .Z(_0125_));
 MUX2_X1 _2504_ (.A(_0682_),
    .B(\mem[10][8] ),
    .S(_0689_),
    .Z(_0126_));
 MUX2_X1 _2505_ (.A(_0684_),
    .B(\mem[10][9] ),
    .S(_0689_),
    .Z(_0127_));
 BUF_X2 _2506_ (.A(_2318_),
    .Z(_0693_));
 NAND2_X2 _2507_ (.A1(_0693_),
    .A2(_0688_),
    .ZN(_0694_));
 BUF_X4 _2508_ (.A(_0694_),
    .Z(_0695_));
 MUX2_X1 _2509_ (.A(_0611_),
    .B(\mem[11][0] ),
    .S(_0695_),
    .Z(_0128_));
 MUX2_X1 _2510_ (.A(_0622_),
    .B(\mem[11][10] ),
    .S(_0695_),
    .Z(_0129_));
 MUX2_X1 _2511_ (.A(_0624_),
    .B(\mem[11][11] ),
    .S(_0695_),
    .Z(_0130_));
 MUX2_X1 _2512_ (.A(_0626_),
    .B(\mem[11][12] ),
    .S(_0695_),
    .Z(_0131_));
 MUX2_X1 _2513_ (.A(_0628_),
    .B(\mem[11][13] ),
    .S(_0695_),
    .Z(_0132_));
 MUX2_X1 _2514_ (.A(_0630_),
    .B(\mem[11][14] ),
    .S(_0695_),
    .Z(_0133_));
 MUX2_X1 _2515_ (.A(_0632_),
    .B(\mem[11][15] ),
    .S(_0695_),
    .Z(_0134_));
 MUX2_X1 _2516_ (.A(_0634_),
    .B(\mem[11][16] ),
    .S(_0695_),
    .Z(_0135_));
 MUX2_X1 _2517_ (.A(_0636_),
    .B(\mem[11][17] ),
    .S(_0695_),
    .Z(_0136_));
 MUX2_X1 _2518_ (.A(_0638_),
    .B(\mem[11][18] ),
    .S(_0695_),
    .Z(_0137_));
 BUF_X4 _2519_ (.A(_0694_),
    .Z(_0696_));
 MUX2_X1 _2520_ (.A(_0640_),
    .B(\mem[11][19] ),
    .S(_0696_),
    .Z(_0138_));
 MUX2_X1 _2521_ (.A(_0643_),
    .B(\mem[11][1] ),
    .S(_0696_),
    .Z(_0139_));
 MUX2_X1 _2522_ (.A(_0645_),
    .B(\mem[11][20] ),
    .S(_0696_),
    .Z(_0140_));
 MUX2_X1 _2523_ (.A(_0647_),
    .B(\mem[11][21] ),
    .S(_0696_),
    .Z(_0141_));
 MUX2_X1 _2524_ (.A(_0649_),
    .B(\mem[11][22] ),
    .S(_0696_),
    .Z(_0142_));
 MUX2_X1 _2525_ (.A(_0651_),
    .B(\mem[11][23] ),
    .S(_0696_),
    .Z(_0143_));
 MUX2_X1 _2526_ (.A(_0653_),
    .B(\mem[11][24] ),
    .S(_0696_),
    .Z(_0144_));
 MUX2_X1 _2527_ (.A(_0655_),
    .B(\mem[11][25] ),
    .S(_0696_),
    .Z(_0145_));
 MUX2_X1 _2528_ (.A(_0657_),
    .B(\mem[11][26] ),
    .S(_0696_),
    .Z(_0146_));
 MUX2_X1 _2529_ (.A(_0659_),
    .B(\mem[11][27] ),
    .S(_0696_),
    .Z(_0147_));
 CLKBUF_X3 _2530_ (.A(_0694_),
    .Z(_0697_));
 MUX2_X1 _2531_ (.A(_0661_),
    .B(\mem[11][28] ),
    .S(_0697_),
    .Z(_0148_));
 MUX2_X1 _2532_ (.A(_0664_),
    .B(\mem[11][29] ),
    .S(_0697_),
    .Z(_0149_));
 MUX2_X1 _2533_ (.A(_0666_),
    .B(\mem[11][2] ),
    .S(_0697_),
    .Z(_0150_));
 MUX2_X1 _2534_ (.A(_0668_),
    .B(\mem[11][30] ),
    .S(_0697_),
    .Z(_0151_));
 MUX2_X1 _2535_ (.A(_0670_),
    .B(\mem[11][31] ),
    .S(_0697_),
    .Z(_0152_));
 MUX2_X1 _2536_ (.A(_0672_),
    .B(\mem[11][3] ),
    .S(_0697_),
    .Z(_0153_));
 MUX2_X1 _2537_ (.A(_0674_),
    .B(\mem[11][4] ),
    .S(_0697_),
    .Z(_0154_));
 MUX2_X1 _2538_ (.A(_0676_),
    .B(\mem[11][5] ),
    .S(_0697_),
    .Z(_0155_));
 MUX2_X1 _2539_ (.A(_0678_),
    .B(\mem[11][6] ),
    .S(_0697_),
    .Z(_0156_));
 MUX2_X1 _2540_ (.A(_0680_),
    .B(\mem[11][7] ),
    .S(_0697_),
    .Z(_0157_));
 MUX2_X1 _2541_ (.A(_0682_),
    .B(\mem[11][8] ),
    .S(_0694_),
    .Z(_0158_));
 MUX2_X1 _2542_ (.A(_0684_),
    .B(\mem[11][9] ),
    .S(_0694_),
    .Z(_0159_));
 AND3_X1 _2543_ (.A1(_0613_),
    .A2(_0615_),
    .A3(_0616_),
    .ZN(_0698_));
 CLKBUF_X3 _2544_ (.A(_0698_),
    .Z(_0699_));
 NAND2_X4 _2545_ (.A1(_0612_),
    .A2(_0699_),
    .ZN(_0700_));
 BUF_X4 _2546_ (.A(_0700_),
    .Z(_0701_));
 MUX2_X1 _2547_ (.A(_0610_),
    .B(\mem[12][0] ),
    .S(_0701_),
    .Z(_0160_));
 MUX2_X1 _2548_ (.A(_0621_),
    .B(\mem[12][10] ),
    .S(_0701_),
    .Z(_0161_));
 MUX2_X1 _2549_ (.A(_0623_),
    .B(\mem[12][11] ),
    .S(_0701_),
    .Z(_0162_));
 MUX2_X1 _2550_ (.A(_0625_),
    .B(\mem[12][12] ),
    .S(_0701_),
    .Z(_0163_));
 MUX2_X1 _2551_ (.A(_0627_),
    .B(\mem[12][13] ),
    .S(_0701_),
    .Z(_0164_));
 MUX2_X1 _2552_ (.A(_0629_),
    .B(\mem[12][14] ),
    .S(_0701_),
    .Z(_0165_));
 MUX2_X1 _2553_ (.A(_0631_),
    .B(\mem[12][15] ),
    .S(_0701_),
    .Z(_0166_));
 MUX2_X1 _2554_ (.A(_0633_),
    .B(\mem[12][16] ),
    .S(_0701_),
    .Z(_0167_));
 MUX2_X1 _2555_ (.A(_0635_),
    .B(\mem[12][17] ),
    .S(_0701_),
    .Z(_0168_));
 MUX2_X1 _2556_ (.A(_0637_),
    .B(\mem[12][18] ),
    .S(_0701_),
    .Z(_0169_));
 BUF_X4 _2557_ (.A(_0700_),
    .Z(_0702_));
 MUX2_X1 _2558_ (.A(_0639_),
    .B(\mem[12][19] ),
    .S(_0702_),
    .Z(_0170_));
 MUX2_X1 _2559_ (.A(_0642_),
    .B(\mem[12][1] ),
    .S(_0702_),
    .Z(_0171_));
 MUX2_X1 _2560_ (.A(_0644_),
    .B(\mem[12][20] ),
    .S(_0702_),
    .Z(_0172_));
 MUX2_X1 _2561_ (.A(_0646_),
    .B(\mem[12][21] ),
    .S(_0702_),
    .Z(_0173_));
 MUX2_X1 _2562_ (.A(_0648_),
    .B(\mem[12][22] ),
    .S(_0702_),
    .Z(_0174_));
 MUX2_X1 _2563_ (.A(_0650_),
    .B(\mem[12][23] ),
    .S(_0702_),
    .Z(_0175_));
 MUX2_X1 _2564_ (.A(_0652_),
    .B(\mem[12][24] ),
    .S(_0702_),
    .Z(_0176_));
 MUX2_X1 _2565_ (.A(_0654_),
    .B(\mem[12][25] ),
    .S(_0702_),
    .Z(_0177_));
 MUX2_X1 _2566_ (.A(_0656_),
    .B(\mem[12][26] ),
    .S(_0702_),
    .Z(_0178_));
 MUX2_X1 _2567_ (.A(_0658_),
    .B(\mem[12][27] ),
    .S(_0702_),
    .Z(_0179_));
 CLKBUF_X3 _2568_ (.A(_0700_),
    .Z(_0703_));
 MUX2_X1 _2569_ (.A(_0660_),
    .B(\mem[12][28] ),
    .S(_0703_),
    .Z(_0180_));
 MUX2_X1 _2570_ (.A(_0663_),
    .B(\mem[12][29] ),
    .S(_0703_),
    .Z(_0181_));
 MUX2_X1 _2571_ (.A(_0665_),
    .B(\mem[12][2] ),
    .S(_0703_),
    .Z(_0182_));
 MUX2_X1 _2572_ (.A(_0667_),
    .B(\mem[12][30] ),
    .S(_0703_),
    .Z(_0183_));
 MUX2_X1 _2573_ (.A(_0669_),
    .B(\mem[12][31] ),
    .S(_0703_),
    .Z(_0184_));
 MUX2_X1 _2574_ (.A(_0671_),
    .B(\mem[12][3] ),
    .S(_0703_),
    .Z(_0185_));
 MUX2_X1 _2575_ (.A(_0673_),
    .B(\mem[12][4] ),
    .S(_0703_),
    .Z(_0186_));
 MUX2_X1 _2576_ (.A(_0675_),
    .B(\mem[12][5] ),
    .S(_0703_),
    .Z(_0187_));
 MUX2_X1 _2577_ (.A(_0677_),
    .B(\mem[12][6] ),
    .S(_0703_),
    .Z(_0188_));
 MUX2_X1 _2578_ (.A(_0679_),
    .B(\mem[12][7] ),
    .S(_0703_),
    .Z(_0189_));
 MUX2_X1 _2579_ (.A(_0681_),
    .B(\mem[12][8] ),
    .S(_0700_),
    .Z(_0190_));
 MUX2_X1 _2580_ (.A(_0683_),
    .B(\mem[12][9] ),
    .S(_0700_),
    .Z(_0191_));
 BUF_X2 _2581_ (.A(_2316_),
    .Z(_0704_));
 NAND2_X4 _2582_ (.A1(_0704_),
    .A2(_0699_),
    .ZN(_0705_));
 BUF_X4 _2583_ (.A(_0705_),
    .Z(_0706_));
 MUX2_X1 _2584_ (.A(_0610_),
    .B(\mem[13][0] ),
    .S(_0706_),
    .Z(_0192_));
 MUX2_X1 _2585_ (.A(_0621_),
    .B(\mem[13][10] ),
    .S(_0706_),
    .Z(_0193_));
 MUX2_X1 _2586_ (.A(_0623_),
    .B(\mem[13][11] ),
    .S(_0706_),
    .Z(_0194_));
 MUX2_X1 _2587_ (.A(_0625_),
    .B(\mem[13][12] ),
    .S(_0706_),
    .Z(_0195_));
 MUX2_X1 _2588_ (.A(_0627_),
    .B(\mem[13][13] ),
    .S(_0706_),
    .Z(_0196_));
 MUX2_X1 _2589_ (.A(_0629_),
    .B(\mem[13][14] ),
    .S(_0706_),
    .Z(_0197_));
 MUX2_X1 _2590_ (.A(_0631_),
    .B(\mem[13][15] ),
    .S(_0706_),
    .Z(_0198_));
 MUX2_X1 _2591_ (.A(_0633_),
    .B(\mem[13][16] ),
    .S(_0706_),
    .Z(_0199_));
 MUX2_X1 _2592_ (.A(_0635_),
    .B(\mem[13][17] ),
    .S(_0706_),
    .Z(_0200_));
 MUX2_X1 _2593_ (.A(_0637_),
    .B(\mem[13][18] ),
    .S(_0706_),
    .Z(_0201_));
 BUF_X4 _2594_ (.A(_0705_),
    .Z(_0707_));
 MUX2_X1 _2595_ (.A(_0639_),
    .B(\mem[13][19] ),
    .S(_0707_),
    .Z(_0202_));
 MUX2_X1 _2596_ (.A(_0642_),
    .B(\mem[13][1] ),
    .S(_0707_),
    .Z(_0203_));
 MUX2_X1 _2597_ (.A(_0644_),
    .B(\mem[13][20] ),
    .S(_0707_),
    .Z(_0204_));
 MUX2_X1 _2598_ (.A(_0646_),
    .B(\mem[13][21] ),
    .S(_0707_),
    .Z(_0205_));
 MUX2_X1 _2599_ (.A(_0648_),
    .B(\mem[13][22] ),
    .S(_0707_),
    .Z(_0206_));
 MUX2_X1 _2600_ (.A(_0650_),
    .B(\mem[13][23] ),
    .S(_0707_),
    .Z(_0207_));
 MUX2_X1 _2601_ (.A(_0652_),
    .B(\mem[13][24] ),
    .S(_0707_),
    .Z(_0208_));
 MUX2_X1 _2602_ (.A(_0654_),
    .B(\mem[13][25] ),
    .S(_0707_),
    .Z(_0209_));
 MUX2_X1 _2603_ (.A(_0656_),
    .B(\mem[13][26] ),
    .S(_0707_),
    .Z(_0210_));
 MUX2_X1 _2604_ (.A(_0658_),
    .B(\mem[13][27] ),
    .S(_0707_),
    .Z(_0211_));
 CLKBUF_X3 _2605_ (.A(_0705_),
    .Z(_0708_));
 MUX2_X1 _2606_ (.A(_0660_),
    .B(\mem[13][28] ),
    .S(_0708_),
    .Z(_0212_));
 MUX2_X1 _2607_ (.A(_0663_),
    .B(\mem[13][29] ),
    .S(_0708_),
    .Z(_0213_));
 MUX2_X1 _2608_ (.A(_0665_),
    .B(\mem[13][2] ),
    .S(_0708_),
    .Z(_0214_));
 MUX2_X1 _2609_ (.A(_0667_),
    .B(\mem[13][30] ),
    .S(_0708_),
    .Z(_0215_));
 MUX2_X1 _2610_ (.A(_0669_),
    .B(\mem[13][31] ),
    .S(_0708_),
    .Z(_0216_));
 MUX2_X1 _2611_ (.A(_0671_),
    .B(\mem[13][3] ),
    .S(_0708_),
    .Z(_0217_));
 MUX2_X1 _2612_ (.A(_0673_),
    .B(\mem[13][4] ),
    .S(_0708_),
    .Z(_0218_));
 MUX2_X1 _2613_ (.A(_0675_),
    .B(\mem[13][5] ),
    .S(_0708_),
    .Z(_0219_));
 MUX2_X1 _2614_ (.A(_0677_),
    .B(\mem[13][6] ),
    .S(_0708_),
    .Z(_0220_));
 MUX2_X1 _2615_ (.A(_0679_),
    .B(\mem[13][7] ),
    .S(_0708_),
    .Z(_0221_));
 MUX2_X1 _2616_ (.A(_0681_),
    .B(\mem[13][8] ),
    .S(_0705_),
    .Z(_0222_));
 MUX2_X1 _2617_ (.A(_0683_),
    .B(\mem[13][9] ),
    .S(_0705_),
    .Z(_0223_));
 NAND2_X2 _2618_ (.A1(_0685_),
    .A2(_0699_),
    .ZN(_0709_));
 BUF_X4 _2619_ (.A(_0709_),
    .Z(_0710_));
 MUX2_X1 _2620_ (.A(_0610_),
    .B(\mem[14][0] ),
    .S(_0710_),
    .Z(_0224_));
 MUX2_X1 _2621_ (.A(_0621_),
    .B(\mem[14][10] ),
    .S(_0710_),
    .Z(_0225_));
 MUX2_X1 _2622_ (.A(_0623_),
    .B(\mem[14][11] ),
    .S(_0710_),
    .Z(_0226_));
 MUX2_X1 _2623_ (.A(_0625_),
    .B(\mem[14][12] ),
    .S(_0710_),
    .Z(_0227_));
 MUX2_X1 _2624_ (.A(_0627_),
    .B(\mem[14][13] ),
    .S(_0710_),
    .Z(_0228_));
 MUX2_X1 _2625_ (.A(_0629_),
    .B(\mem[14][14] ),
    .S(_0710_),
    .Z(_0229_));
 MUX2_X1 _2626_ (.A(_0631_),
    .B(\mem[14][15] ),
    .S(_0710_),
    .Z(_0230_));
 MUX2_X1 _2627_ (.A(_0633_),
    .B(\mem[14][16] ),
    .S(_0710_),
    .Z(_0231_));
 MUX2_X1 _2628_ (.A(_0635_),
    .B(\mem[14][17] ),
    .S(_0710_),
    .Z(_0232_));
 MUX2_X1 _2629_ (.A(_0637_),
    .B(\mem[14][18] ),
    .S(_0710_),
    .Z(_0233_));
 BUF_X4 _2630_ (.A(_0709_),
    .Z(_0711_));
 MUX2_X1 _2631_ (.A(_0639_),
    .B(\mem[14][19] ),
    .S(_0711_),
    .Z(_0234_));
 MUX2_X1 _2632_ (.A(_0642_),
    .B(\mem[14][1] ),
    .S(_0711_),
    .Z(_0235_));
 MUX2_X1 _2633_ (.A(_0644_),
    .B(\mem[14][20] ),
    .S(_0711_),
    .Z(_0236_));
 MUX2_X1 _2634_ (.A(_0646_),
    .B(\mem[14][21] ),
    .S(_0711_),
    .Z(_0237_));
 MUX2_X1 _2635_ (.A(_0648_),
    .B(\mem[14][22] ),
    .S(_0711_),
    .Z(_0238_));
 MUX2_X1 _2636_ (.A(_0650_),
    .B(\mem[14][23] ),
    .S(_0711_),
    .Z(_0239_));
 MUX2_X1 _2637_ (.A(_0652_),
    .B(\mem[14][24] ),
    .S(_0711_),
    .Z(_0240_));
 MUX2_X1 _2638_ (.A(_0654_),
    .B(\mem[14][25] ),
    .S(_0711_),
    .Z(_0241_));
 MUX2_X1 _2639_ (.A(_0656_),
    .B(\mem[14][26] ),
    .S(_0711_),
    .Z(_0242_));
 MUX2_X1 _2640_ (.A(_0658_),
    .B(\mem[14][27] ),
    .S(_0711_),
    .Z(_0243_));
 CLKBUF_X3 _2641_ (.A(_0709_),
    .Z(_0712_));
 MUX2_X1 _2642_ (.A(_0660_),
    .B(\mem[14][28] ),
    .S(_0712_),
    .Z(_0244_));
 MUX2_X1 _2643_ (.A(_0663_),
    .B(\mem[14][29] ),
    .S(_0712_),
    .Z(_0245_));
 MUX2_X1 _2644_ (.A(_0665_),
    .B(\mem[14][2] ),
    .S(_0712_),
    .Z(_0246_));
 MUX2_X1 _2645_ (.A(_0667_),
    .B(\mem[14][30] ),
    .S(_0712_),
    .Z(_0247_));
 MUX2_X1 _2646_ (.A(_0669_),
    .B(\mem[14][31] ),
    .S(_0712_),
    .Z(_0248_));
 MUX2_X1 _2647_ (.A(_0671_),
    .B(\mem[14][3] ),
    .S(_0712_),
    .Z(_0249_));
 MUX2_X1 _2648_ (.A(_0673_),
    .B(\mem[14][4] ),
    .S(_0712_),
    .Z(_0250_));
 MUX2_X1 _2649_ (.A(_0675_),
    .B(\mem[14][5] ),
    .S(_0712_),
    .Z(_0251_));
 MUX2_X1 _2650_ (.A(_0677_),
    .B(\mem[14][6] ),
    .S(_0712_),
    .Z(_0252_));
 MUX2_X1 _2651_ (.A(_0679_),
    .B(\mem[14][7] ),
    .S(_0712_),
    .Z(_0253_));
 MUX2_X1 _2652_ (.A(_0681_),
    .B(\mem[14][8] ),
    .S(_0709_),
    .Z(_0254_));
 MUX2_X1 _2653_ (.A(_0683_),
    .B(\mem[14][9] ),
    .S(_0709_),
    .Z(_0255_));
 NAND2_X4 _2654_ (.A1(_0693_),
    .A2(_0699_),
    .ZN(_0713_));
 BUF_X4 _2655_ (.A(_0713_),
    .Z(_0714_));
 MUX2_X1 _2656_ (.A(_0610_),
    .B(\mem[15][0] ),
    .S(_0714_),
    .Z(_0256_));
 MUX2_X1 _2657_ (.A(_0621_),
    .B(\mem[15][10] ),
    .S(_0714_),
    .Z(_0257_));
 MUX2_X1 _2658_ (.A(_0623_),
    .B(\mem[15][11] ),
    .S(_0714_),
    .Z(_0258_));
 MUX2_X1 _2659_ (.A(_0625_),
    .B(\mem[15][12] ),
    .S(_0714_),
    .Z(_0259_));
 MUX2_X1 _2660_ (.A(_0627_),
    .B(\mem[15][13] ),
    .S(_0714_),
    .Z(_0260_));
 MUX2_X1 _2661_ (.A(_0629_),
    .B(\mem[15][14] ),
    .S(_0714_),
    .Z(_0261_));
 MUX2_X1 _2662_ (.A(_0631_),
    .B(\mem[15][15] ),
    .S(_0714_),
    .Z(_0262_));
 MUX2_X1 _2663_ (.A(_0633_),
    .B(\mem[15][16] ),
    .S(_0714_),
    .Z(_0263_));
 MUX2_X1 _2664_ (.A(_0635_),
    .B(\mem[15][17] ),
    .S(_0714_),
    .Z(_0264_));
 MUX2_X1 _2665_ (.A(_0637_),
    .B(\mem[15][18] ),
    .S(_0714_),
    .Z(_0265_));
 BUF_X4 _2666_ (.A(_0713_),
    .Z(_0715_));
 MUX2_X1 _2667_ (.A(_0639_),
    .B(\mem[15][19] ),
    .S(_0715_),
    .Z(_0266_));
 MUX2_X1 _2668_ (.A(_0642_),
    .B(\mem[15][1] ),
    .S(_0715_),
    .Z(_0267_));
 MUX2_X1 _2669_ (.A(_0644_),
    .B(\mem[15][20] ),
    .S(_0715_),
    .Z(_0268_));
 MUX2_X1 _2670_ (.A(_0646_),
    .B(\mem[15][21] ),
    .S(_0715_),
    .Z(_0269_));
 MUX2_X1 _2671_ (.A(_0648_),
    .B(\mem[15][22] ),
    .S(_0715_),
    .Z(_0270_));
 MUX2_X1 _2672_ (.A(_0650_),
    .B(\mem[15][23] ),
    .S(_0715_),
    .Z(_0271_));
 MUX2_X1 _2673_ (.A(_0652_),
    .B(\mem[15][24] ),
    .S(_0715_),
    .Z(_0272_));
 MUX2_X1 _2674_ (.A(_0654_),
    .B(\mem[15][25] ),
    .S(_0715_),
    .Z(_0273_));
 MUX2_X1 _2675_ (.A(_0656_),
    .B(\mem[15][26] ),
    .S(_0715_),
    .Z(_0274_));
 MUX2_X1 _2676_ (.A(_0658_),
    .B(\mem[15][27] ),
    .S(_0715_),
    .Z(_0275_));
 CLKBUF_X3 _2677_ (.A(_0713_),
    .Z(_0716_));
 MUX2_X1 _2678_ (.A(_0660_),
    .B(\mem[15][28] ),
    .S(_0716_),
    .Z(_0276_));
 MUX2_X1 _2679_ (.A(_0663_),
    .B(\mem[15][29] ),
    .S(_0716_),
    .Z(_0277_));
 MUX2_X1 _2680_ (.A(_0665_),
    .B(\mem[15][2] ),
    .S(_0716_),
    .Z(_0278_));
 MUX2_X1 _2681_ (.A(_0667_),
    .B(\mem[15][30] ),
    .S(_0716_),
    .Z(_0279_));
 MUX2_X1 _2682_ (.A(_0669_),
    .B(\mem[15][31] ),
    .S(_0716_),
    .Z(_0280_));
 MUX2_X1 _2683_ (.A(_0671_),
    .B(\mem[15][3] ),
    .S(_0716_),
    .Z(_0281_));
 MUX2_X1 _2684_ (.A(_0673_),
    .B(\mem[15][4] ),
    .S(_0716_),
    .Z(_0282_));
 MUX2_X1 _2685_ (.A(_0675_),
    .B(\mem[15][5] ),
    .S(_0716_),
    .Z(_0283_));
 MUX2_X1 _2686_ (.A(_0677_),
    .B(\mem[15][6] ),
    .S(_0716_),
    .Z(_0284_));
 MUX2_X1 _2687_ (.A(_0679_),
    .B(\mem[15][7] ),
    .S(_0716_),
    .Z(_0285_));
 MUX2_X1 _2688_ (.A(_0681_),
    .B(\mem[15][8] ),
    .S(_0713_),
    .Z(_0286_));
 MUX2_X1 _2689_ (.A(_0683_),
    .B(\mem[15][9] ),
    .S(_0713_),
    .Z(_0287_));
 AND2_X1 _2690_ (.A1(_0704_),
    .A2(_0617_),
    .ZN(_0717_));
 BUF_X2 _2691_ (.A(_0717_),
    .Z(_0718_));
 BUF_X4 _2692_ (.A(_0718_),
    .Z(_0719_));
 MUX2_X1 _2693_ (.A(\mem[1][0] ),
    .B(_0611_),
    .S(_0719_),
    .Z(_0288_));
 MUX2_X1 _2694_ (.A(\mem[1][10] ),
    .B(_0622_),
    .S(_0719_),
    .Z(_0289_));
 MUX2_X1 _2695_ (.A(\mem[1][11] ),
    .B(_0624_),
    .S(_0719_),
    .Z(_0290_));
 MUX2_X1 _2696_ (.A(\mem[1][12] ),
    .B(_0626_),
    .S(_0719_),
    .Z(_0291_));
 MUX2_X1 _2697_ (.A(\mem[1][13] ),
    .B(_0628_),
    .S(_0719_),
    .Z(_0292_));
 MUX2_X1 _2698_ (.A(\mem[1][14] ),
    .B(_0630_),
    .S(_0719_),
    .Z(_0293_));
 MUX2_X1 _2699_ (.A(\mem[1][15] ),
    .B(_0632_),
    .S(_0719_),
    .Z(_0294_));
 MUX2_X1 _2700_ (.A(\mem[1][16] ),
    .B(_0634_),
    .S(_0719_),
    .Z(_0295_));
 MUX2_X1 _2701_ (.A(\mem[1][17] ),
    .B(_0636_),
    .S(_0719_),
    .Z(_0296_));
 MUX2_X1 _2702_ (.A(\mem[1][18] ),
    .B(_0638_),
    .S(_0719_),
    .Z(_0297_));
 BUF_X4 _2703_ (.A(_0718_),
    .Z(_0720_));
 MUX2_X1 _2704_ (.A(\mem[1][19] ),
    .B(_0640_),
    .S(_0720_),
    .Z(_0298_));
 MUX2_X1 _2705_ (.A(\mem[1][1] ),
    .B(_0643_),
    .S(_0720_),
    .Z(_0299_));
 MUX2_X1 _2706_ (.A(\mem[1][20] ),
    .B(_0645_),
    .S(_0720_),
    .Z(_0300_));
 MUX2_X1 _2707_ (.A(\mem[1][21] ),
    .B(_0647_),
    .S(_0720_),
    .Z(_0301_));
 MUX2_X1 _2708_ (.A(\mem[1][22] ),
    .B(_0649_),
    .S(_0720_),
    .Z(_0302_));
 MUX2_X1 _2709_ (.A(\mem[1][23] ),
    .B(_0651_),
    .S(_0720_),
    .Z(_0303_));
 MUX2_X1 _2710_ (.A(\mem[1][24] ),
    .B(_0653_),
    .S(_0720_),
    .Z(_0304_));
 MUX2_X1 _2711_ (.A(\mem[1][25] ),
    .B(_0655_),
    .S(_0720_),
    .Z(_0305_));
 MUX2_X1 _2712_ (.A(\mem[1][26] ),
    .B(_0657_),
    .S(_0720_),
    .Z(_0306_));
 MUX2_X1 _2713_ (.A(\mem[1][27] ),
    .B(_0659_),
    .S(_0720_),
    .Z(_0307_));
 CLKBUF_X3 _2714_ (.A(_0718_),
    .Z(_0721_));
 MUX2_X1 _2715_ (.A(\mem[1][28] ),
    .B(_0661_),
    .S(_0721_),
    .Z(_0308_));
 MUX2_X1 _2716_ (.A(\mem[1][29] ),
    .B(_0664_),
    .S(_0721_),
    .Z(_0309_));
 MUX2_X1 _2717_ (.A(\mem[1][2] ),
    .B(_0666_),
    .S(_0721_),
    .Z(_0310_));
 MUX2_X1 _2718_ (.A(\mem[1][30] ),
    .B(_0668_),
    .S(_0721_),
    .Z(_0311_));
 MUX2_X1 _2719_ (.A(\mem[1][31] ),
    .B(_0670_),
    .S(_0721_),
    .Z(_0312_));
 MUX2_X1 _2720_ (.A(\mem[1][3] ),
    .B(_0672_),
    .S(_0721_),
    .Z(_0313_));
 MUX2_X1 _2721_ (.A(\mem[1][4] ),
    .B(_0674_),
    .S(_0721_),
    .Z(_0314_));
 MUX2_X1 _2722_ (.A(\mem[1][5] ),
    .B(_0676_),
    .S(_0721_),
    .Z(_0315_));
 MUX2_X1 _2723_ (.A(\mem[1][6] ),
    .B(_0678_),
    .S(_0721_),
    .Z(_0316_));
 MUX2_X1 _2724_ (.A(\mem[1][7] ),
    .B(_0680_),
    .S(_0721_),
    .Z(_0317_));
 MUX2_X1 _2725_ (.A(\mem[1][8] ),
    .B(_0682_),
    .S(_0718_),
    .Z(_0318_));
 MUX2_X1 _2726_ (.A(\mem[1][9] ),
    .B(_0684_),
    .S(_0718_),
    .Z(_0319_));
 AND2_X1 _2727_ (.A1(_0685_),
    .A2(_0617_),
    .ZN(_0722_));
 BUF_X2 _2728_ (.A(_0722_),
    .Z(_0723_));
 BUF_X4 _2729_ (.A(_0723_),
    .Z(_0724_));
 MUX2_X1 _2730_ (.A(\mem[2][0] ),
    .B(_0611_),
    .S(_0724_),
    .Z(_0320_));
 MUX2_X1 _2731_ (.A(\mem[2][10] ),
    .B(_0622_),
    .S(_0724_),
    .Z(_0321_));
 MUX2_X1 _2732_ (.A(\mem[2][11] ),
    .B(_0624_),
    .S(_0724_),
    .Z(_0322_));
 MUX2_X1 _2733_ (.A(\mem[2][12] ),
    .B(_0626_),
    .S(_0724_),
    .Z(_0323_));
 MUX2_X1 _2734_ (.A(\mem[2][13] ),
    .B(_0628_),
    .S(_0724_),
    .Z(_0324_));
 MUX2_X1 _2735_ (.A(\mem[2][14] ),
    .B(_0630_),
    .S(_0724_),
    .Z(_0325_));
 MUX2_X1 _2736_ (.A(\mem[2][15] ),
    .B(_0632_),
    .S(_0724_),
    .Z(_0326_));
 MUX2_X1 _2737_ (.A(\mem[2][16] ),
    .B(_0634_),
    .S(_0724_),
    .Z(_0327_));
 MUX2_X1 _2738_ (.A(\mem[2][17] ),
    .B(_0636_),
    .S(_0724_),
    .Z(_0328_));
 MUX2_X1 _2739_ (.A(\mem[2][18] ),
    .B(_0638_),
    .S(_0724_),
    .Z(_0329_));
 BUF_X4 _2740_ (.A(_0723_),
    .Z(_0725_));
 MUX2_X1 _2741_ (.A(\mem[2][19] ),
    .B(_0640_),
    .S(_0725_),
    .Z(_0330_));
 MUX2_X1 _2742_ (.A(\mem[2][1] ),
    .B(_0643_),
    .S(_0725_),
    .Z(_0331_));
 MUX2_X1 _2743_ (.A(\mem[2][20] ),
    .B(_0645_),
    .S(_0725_),
    .Z(_0332_));
 MUX2_X1 _2744_ (.A(\mem[2][21] ),
    .B(_0647_),
    .S(_0725_),
    .Z(_0333_));
 MUX2_X1 _2745_ (.A(\mem[2][22] ),
    .B(_0649_),
    .S(_0725_),
    .Z(_0334_));
 MUX2_X1 _2746_ (.A(\mem[2][23] ),
    .B(_0651_),
    .S(_0725_),
    .Z(_0335_));
 MUX2_X1 _2747_ (.A(\mem[2][24] ),
    .B(_0653_),
    .S(_0725_),
    .Z(_0336_));
 MUX2_X1 _2748_ (.A(\mem[2][25] ),
    .B(_0655_),
    .S(_0725_),
    .Z(_0337_));
 MUX2_X1 _2749_ (.A(\mem[2][26] ),
    .B(_0657_),
    .S(_0725_),
    .Z(_0338_));
 MUX2_X1 _2750_ (.A(\mem[2][27] ),
    .B(_0659_),
    .S(_0725_),
    .Z(_0339_));
 BUF_X4 _2751_ (.A(_0723_),
    .Z(_0726_));
 MUX2_X1 _2752_ (.A(\mem[2][28] ),
    .B(_0661_),
    .S(_0726_),
    .Z(_0340_));
 MUX2_X1 _2753_ (.A(\mem[2][29] ),
    .B(_0664_),
    .S(_0726_),
    .Z(_0341_));
 MUX2_X1 _2754_ (.A(\mem[2][2] ),
    .B(_0666_),
    .S(_0726_),
    .Z(_0342_));
 MUX2_X1 _2755_ (.A(\mem[2][30] ),
    .B(_0668_),
    .S(_0726_),
    .Z(_0343_));
 MUX2_X1 _2756_ (.A(\mem[2][31] ),
    .B(_0670_),
    .S(_0726_),
    .Z(_0344_));
 MUX2_X1 _2757_ (.A(\mem[2][3] ),
    .B(_0672_),
    .S(_0726_),
    .Z(_0345_));
 MUX2_X1 _2758_ (.A(\mem[2][4] ),
    .B(_0674_),
    .S(_0726_),
    .Z(_0346_));
 MUX2_X1 _2759_ (.A(\mem[2][5] ),
    .B(_0676_),
    .S(_0726_),
    .Z(_0347_));
 MUX2_X1 _2760_ (.A(\mem[2][6] ),
    .B(_0678_),
    .S(_0726_),
    .Z(_0348_));
 MUX2_X1 _2761_ (.A(\mem[2][7] ),
    .B(_0680_),
    .S(_0726_),
    .Z(_0349_));
 MUX2_X1 _2762_ (.A(\mem[2][8] ),
    .B(_0682_),
    .S(_0723_),
    .Z(_0350_));
 MUX2_X1 _2763_ (.A(\mem[2][9] ),
    .B(_0684_),
    .S(_0723_),
    .Z(_0351_));
 AND2_X1 _2764_ (.A1(_0693_),
    .A2(_0617_),
    .ZN(_0727_));
 BUF_X2 _2765_ (.A(_0727_),
    .Z(_0728_));
 BUF_X4 _2766_ (.A(_0728_),
    .Z(_0729_));
 MUX2_X1 _2767_ (.A(\mem[3][0] ),
    .B(_0611_),
    .S(_0729_),
    .Z(_0352_));
 MUX2_X1 _2768_ (.A(\mem[3][10] ),
    .B(_0622_),
    .S(_0729_),
    .Z(_0353_));
 MUX2_X1 _2769_ (.A(\mem[3][11] ),
    .B(_0624_),
    .S(_0729_),
    .Z(_0354_));
 MUX2_X1 _2770_ (.A(\mem[3][12] ),
    .B(_0626_),
    .S(_0729_),
    .Z(_0355_));
 MUX2_X1 _2771_ (.A(\mem[3][13] ),
    .B(_0628_),
    .S(_0729_),
    .Z(_0356_));
 MUX2_X1 _2772_ (.A(\mem[3][14] ),
    .B(_0630_),
    .S(_0729_),
    .Z(_0357_));
 MUX2_X1 _2773_ (.A(\mem[3][15] ),
    .B(_0632_),
    .S(_0729_),
    .Z(_0358_));
 MUX2_X1 _2774_ (.A(\mem[3][16] ),
    .B(_0634_),
    .S(_0729_),
    .Z(_0359_));
 MUX2_X1 _2775_ (.A(\mem[3][17] ),
    .B(_0636_),
    .S(_0729_),
    .Z(_0360_));
 MUX2_X1 _2776_ (.A(\mem[3][18] ),
    .B(_0638_),
    .S(_0729_),
    .Z(_0361_));
 BUF_X4 _2777_ (.A(_0728_),
    .Z(_0730_));
 MUX2_X1 _2778_ (.A(\mem[3][19] ),
    .B(_0640_),
    .S(_0730_),
    .Z(_0362_));
 MUX2_X1 _2779_ (.A(\mem[3][1] ),
    .B(_0643_),
    .S(_0730_),
    .Z(_0363_));
 MUX2_X1 _2780_ (.A(\mem[3][20] ),
    .B(_0645_),
    .S(_0730_),
    .Z(_0364_));
 MUX2_X1 _2781_ (.A(\mem[3][21] ),
    .B(_0647_),
    .S(_0730_),
    .Z(_0365_));
 MUX2_X1 _2782_ (.A(\mem[3][22] ),
    .B(_0649_),
    .S(_0730_),
    .Z(_0366_));
 MUX2_X1 _2783_ (.A(\mem[3][23] ),
    .B(_0651_),
    .S(_0730_),
    .Z(_0367_));
 MUX2_X1 _2784_ (.A(\mem[3][24] ),
    .B(_0653_),
    .S(_0730_),
    .Z(_0368_));
 MUX2_X1 _2785_ (.A(\mem[3][25] ),
    .B(_0655_),
    .S(_0730_),
    .Z(_0369_));
 MUX2_X1 _2786_ (.A(\mem[3][26] ),
    .B(_0657_),
    .S(_0730_),
    .Z(_0370_));
 MUX2_X1 _2787_ (.A(\mem[3][27] ),
    .B(_0659_),
    .S(_0730_),
    .Z(_0371_));
 BUF_X4 _2788_ (.A(_0728_),
    .Z(_0731_));
 MUX2_X1 _2789_ (.A(\mem[3][28] ),
    .B(_0661_),
    .S(_0731_),
    .Z(_0372_));
 MUX2_X1 _2790_ (.A(\mem[3][29] ),
    .B(_0664_),
    .S(_0731_),
    .Z(_0373_));
 MUX2_X1 _2791_ (.A(\mem[3][2] ),
    .B(_0666_),
    .S(_0731_),
    .Z(_0374_));
 MUX2_X1 _2792_ (.A(\mem[3][30] ),
    .B(_0668_),
    .S(_0731_),
    .Z(_0375_));
 MUX2_X1 _2793_ (.A(\mem[3][31] ),
    .B(_0670_),
    .S(_0731_),
    .Z(_0376_));
 MUX2_X1 _2794_ (.A(\mem[3][3] ),
    .B(_0672_),
    .S(_0731_),
    .Z(_0377_));
 MUX2_X1 _2795_ (.A(\mem[3][4] ),
    .B(_0674_),
    .S(_0731_),
    .Z(_0378_));
 MUX2_X1 _2796_ (.A(\mem[3][5] ),
    .B(_0676_),
    .S(_0731_),
    .Z(_0379_));
 MUX2_X1 _2797_ (.A(\mem[3][6] ),
    .B(_0678_),
    .S(_0731_),
    .Z(_0380_));
 MUX2_X1 _2798_ (.A(\mem[3][7] ),
    .B(_0680_),
    .S(_0731_),
    .Z(_0381_));
 MUX2_X1 _2799_ (.A(\mem[3][8] ),
    .B(_0682_),
    .S(_0728_),
    .Z(_0382_));
 MUX2_X1 _2800_ (.A(\mem[3][9] ),
    .B(_0684_),
    .S(_0728_),
    .Z(_0383_));
 NOR3_X2 _2801_ (.A1(_0614_),
    .A2(_0615_),
    .A3(_0686_),
    .ZN(_0732_));
 AND2_X1 _2802_ (.A1(_0612_),
    .A2(_0732_),
    .ZN(_0733_));
 CLKBUF_X3 _2803_ (.A(_0733_),
    .Z(_0734_));
 BUF_X4 _2804_ (.A(_0734_),
    .Z(_0735_));
 MUX2_X1 _2805_ (.A(\mem[4][0] ),
    .B(_0611_),
    .S(_0735_),
    .Z(_0384_));
 MUX2_X1 _2806_ (.A(\mem[4][10] ),
    .B(_0622_),
    .S(_0735_),
    .Z(_0385_));
 MUX2_X1 _2807_ (.A(\mem[4][11] ),
    .B(_0624_),
    .S(_0735_),
    .Z(_0386_));
 MUX2_X1 _2808_ (.A(\mem[4][12] ),
    .B(_0626_),
    .S(_0735_),
    .Z(_0387_));
 MUX2_X1 _2809_ (.A(\mem[4][13] ),
    .B(_0628_),
    .S(_0735_),
    .Z(_0388_));
 MUX2_X1 _2810_ (.A(\mem[4][14] ),
    .B(_0630_),
    .S(_0735_),
    .Z(_0389_));
 MUX2_X1 _2811_ (.A(\mem[4][15] ),
    .B(_0632_),
    .S(_0735_),
    .Z(_0390_));
 MUX2_X1 _2812_ (.A(\mem[4][16] ),
    .B(_0634_),
    .S(_0735_),
    .Z(_0391_));
 MUX2_X1 _2813_ (.A(\mem[4][17] ),
    .B(_0636_),
    .S(_0735_),
    .Z(_0392_));
 MUX2_X1 _2814_ (.A(\mem[4][18] ),
    .B(_0638_),
    .S(_0735_),
    .Z(_0393_));
 BUF_X4 _2815_ (.A(_0734_),
    .Z(_0736_));
 MUX2_X1 _2816_ (.A(\mem[4][19] ),
    .B(_0640_),
    .S(_0736_),
    .Z(_0394_));
 MUX2_X1 _2817_ (.A(\mem[4][1] ),
    .B(_0643_),
    .S(_0736_),
    .Z(_0395_));
 MUX2_X1 _2818_ (.A(\mem[4][20] ),
    .B(_0645_),
    .S(_0736_),
    .Z(_0396_));
 MUX2_X1 _2819_ (.A(\mem[4][21] ),
    .B(_0647_),
    .S(_0736_),
    .Z(_0397_));
 MUX2_X1 _2820_ (.A(\mem[4][22] ),
    .B(_0649_),
    .S(_0736_),
    .Z(_0398_));
 MUX2_X1 _2821_ (.A(\mem[4][23] ),
    .B(_0651_),
    .S(_0736_),
    .Z(_0399_));
 MUX2_X1 _2822_ (.A(\mem[4][24] ),
    .B(_0653_),
    .S(_0736_),
    .Z(_0400_));
 MUX2_X1 _2823_ (.A(\mem[4][25] ),
    .B(_0655_),
    .S(_0736_),
    .Z(_0401_));
 MUX2_X1 _2824_ (.A(\mem[4][26] ),
    .B(_0657_),
    .S(_0736_),
    .Z(_0402_));
 MUX2_X1 _2825_ (.A(\mem[4][27] ),
    .B(_0659_),
    .S(_0736_),
    .Z(_0403_));
 BUF_X4 _2826_ (.A(_0734_),
    .Z(_0737_));
 MUX2_X1 _2827_ (.A(\mem[4][28] ),
    .B(_0661_),
    .S(_0737_),
    .Z(_0404_));
 MUX2_X1 _2828_ (.A(\mem[4][29] ),
    .B(_0664_),
    .S(_0737_),
    .Z(_0405_));
 MUX2_X1 _2829_ (.A(\mem[4][2] ),
    .B(_0666_),
    .S(_0737_),
    .Z(_0406_));
 MUX2_X1 _2830_ (.A(\mem[4][30] ),
    .B(_0668_),
    .S(_0737_),
    .Z(_0407_));
 MUX2_X1 _2831_ (.A(\mem[4][31] ),
    .B(_0670_),
    .S(_0737_),
    .Z(_0408_));
 MUX2_X1 _2832_ (.A(\mem[4][3] ),
    .B(_0672_),
    .S(_0737_),
    .Z(_0409_));
 MUX2_X1 _2833_ (.A(\mem[4][4] ),
    .B(_0674_),
    .S(_0737_),
    .Z(_0410_));
 MUX2_X1 _2834_ (.A(\mem[4][5] ),
    .B(_0676_),
    .S(_0737_),
    .Z(_0411_));
 MUX2_X1 _2835_ (.A(\mem[4][6] ),
    .B(_0678_),
    .S(_0737_),
    .Z(_0412_));
 MUX2_X1 _2836_ (.A(\mem[4][7] ),
    .B(_0680_),
    .S(_0737_),
    .Z(_0413_));
 MUX2_X1 _2837_ (.A(\mem[4][8] ),
    .B(_0682_),
    .S(_0734_),
    .Z(_0414_));
 MUX2_X1 _2838_ (.A(\mem[4][9] ),
    .B(_0684_),
    .S(_0734_),
    .Z(_0415_));
 AND2_X1 _2839_ (.A1(_0704_),
    .A2(_0732_),
    .ZN(_0738_));
 BUF_X2 _2840_ (.A(_0738_),
    .Z(_0739_));
 BUF_X4 _2841_ (.A(_0739_),
    .Z(_0740_));
 MUX2_X1 _2842_ (.A(\mem[5][0] ),
    .B(_0611_),
    .S(_0740_),
    .Z(_0416_));
 MUX2_X1 _2843_ (.A(\mem[5][10] ),
    .B(_0622_),
    .S(_0740_),
    .Z(_0417_));
 MUX2_X1 _2844_ (.A(\mem[5][11] ),
    .B(_0624_),
    .S(_0740_),
    .Z(_0418_));
 MUX2_X1 _2845_ (.A(\mem[5][12] ),
    .B(_0626_),
    .S(_0740_),
    .Z(_0419_));
 MUX2_X1 _2846_ (.A(\mem[5][13] ),
    .B(_0628_),
    .S(_0740_),
    .Z(_0420_));
 MUX2_X1 _2847_ (.A(\mem[5][14] ),
    .B(_0630_),
    .S(_0740_),
    .Z(_0421_));
 MUX2_X1 _2848_ (.A(\mem[5][15] ),
    .B(_0632_),
    .S(_0740_),
    .Z(_0422_));
 MUX2_X1 _2849_ (.A(\mem[5][16] ),
    .B(_0634_),
    .S(_0740_),
    .Z(_0423_));
 MUX2_X1 _2850_ (.A(\mem[5][17] ),
    .B(_0636_),
    .S(_0740_),
    .Z(_0424_));
 MUX2_X1 _2851_ (.A(\mem[5][18] ),
    .B(_0638_),
    .S(_0740_),
    .Z(_0425_));
 BUF_X4 _2852_ (.A(_0739_),
    .Z(_0741_));
 MUX2_X1 _2853_ (.A(\mem[5][19] ),
    .B(_0640_),
    .S(_0741_),
    .Z(_0426_));
 MUX2_X1 _2854_ (.A(\mem[5][1] ),
    .B(_0643_),
    .S(_0741_),
    .Z(_0427_));
 MUX2_X1 _2855_ (.A(\mem[5][20] ),
    .B(_0645_),
    .S(_0741_),
    .Z(_0428_));
 MUX2_X1 _2856_ (.A(\mem[5][21] ),
    .B(_0647_),
    .S(_0741_),
    .Z(_0429_));
 MUX2_X1 _2857_ (.A(\mem[5][22] ),
    .B(_0649_),
    .S(_0741_),
    .Z(_0430_));
 MUX2_X1 _2858_ (.A(\mem[5][23] ),
    .B(_0651_),
    .S(_0741_),
    .Z(_0431_));
 MUX2_X1 _2859_ (.A(\mem[5][24] ),
    .B(_0653_),
    .S(_0741_),
    .Z(_0432_));
 MUX2_X1 _2860_ (.A(\mem[5][25] ),
    .B(_0655_),
    .S(_0741_),
    .Z(_0433_));
 MUX2_X1 _2861_ (.A(\mem[5][26] ),
    .B(_0657_),
    .S(_0741_),
    .Z(_0434_));
 MUX2_X1 _2862_ (.A(\mem[5][27] ),
    .B(_0659_),
    .S(_0741_),
    .Z(_0435_));
 CLKBUF_X3 _2863_ (.A(_0739_),
    .Z(_0742_));
 MUX2_X1 _2864_ (.A(\mem[5][28] ),
    .B(_0661_),
    .S(_0742_),
    .Z(_0436_));
 MUX2_X1 _2865_ (.A(\mem[5][29] ),
    .B(_0664_),
    .S(_0742_),
    .Z(_0437_));
 MUX2_X1 _2866_ (.A(\mem[5][2] ),
    .B(_0666_),
    .S(_0742_),
    .Z(_0438_));
 MUX2_X1 _2867_ (.A(\mem[5][30] ),
    .B(_0668_),
    .S(_0742_),
    .Z(_0439_));
 MUX2_X1 _2868_ (.A(\mem[5][31] ),
    .B(_0670_),
    .S(_0742_),
    .Z(_0440_));
 MUX2_X1 _2869_ (.A(\mem[5][3] ),
    .B(_0672_),
    .S(_0742_),
    .Z(_0441_));
 MUX2_X1 _2870_ (.A(\mem[5][4] ),
    .B(_0674_),
    .S(_0742_),
    .Z(_0442_));
 MUX2_X1 _2871_ (.A(\mem[5][5] ),
    .B(_0676_),
    .S(_0742_),
    .Z(_0443_));
 MUX2_X1 _2872_ (.A(\mem[5][6] ),
    .B(_0678_),
    .S(_0742_),
    .Z(_0444_));
 MUX2_X1 _2873_ (.A(\mem[5][7] ),
    .B(_0680_),
    .S(_0742_),
    .Z(_0445_));
 MUX2_X1 _2874_ (.A(\mem[5][8] ),
    .B(_0682_),
    .S(_0739_),
    .Z(_0446_));
 MUX2_X1 _2875_ (.A(\mem[5][9] ),
    .B(_0684_),
    .S(_0739_),
    .Z(_0447_));
 AND2_X1 _2876_ (.A1(_0685_),
    .A2(_0732_),
    .ZN(_0743_));
 BUF_X2 _2877_ (.A(_0743_),
    .Z(_0744_));
 BUF_X4 _2878_ (.A(_0744_),
    .Z(_0745_));
 MUX2_X1 _2879_ (.A(\mem[6][0] ),
    .B(_0611_),
    .S(_0745_),
    .Z(_0448_));
 MUX2_X1 _2880_ (.A(\mem[6][10] ),
    .B(_0622_),
    .S(_0745_),
    .Z(_0449_));
 MUX2_X1 _2881_ (.A(\mem[6][11] ),
    .B(_0624_),
    .S(_0745_),
    .Z(_0450_));
 MUX2_X1 _2882_ (.A(\mem[6][12] ),
    .B(_0626_),
    .S(_0745_),
    .Z(_0451_));
 MUX2_X1 _2883_ (.A(\mem[6][13] ),
    .B(_0628_),
    .S(_0745_),
    .Z(_0452_));
 MUX2_X1 _2884_ (.A(\mem[6][14] ),
    .B(_0630_),
    .S(_0745_),
    .Z(_0453_));
 MUX2_X1 _2885_ (.A(\mem[6][15] ),
    .B(_0632_),
    .S(_0745_),
    .Z(_0454_));
 MUX2_X1 _2886_ (.A(\mem[6][16] ),
    .B(_0634_),
    .S(_0745_),
    .Z(_0455_));
 MUX2_X1 _2887_ (.A(\mem[6][17] ),
    .B(_0636_),
    .S(_0745_),
    .Z(_0456_));
 MUX2_X1 _2888_ (.A(\mem[6][18] ),
    .B(_0638_),
    .S(_0745_),
    .Z(_0457_));
 BUF_X4 _2889_ (.A(_0744_),
    .Z(_0746_));
 MUX2_X1 _2890_ (.A(\mem[6][19] ),
    .B(_0640_),
    .S(_0746_),
    .Z(_0458_));
 MUX2_X1 _2891_ (.A(\mem[6][1] ),
    .B(_0643_),
    .S(_0746_),
    .Z(_0459_));
 MUX2_X1 _2892_ (.A(\mem[6][20] ),
    .B(_0645_),
    .S(_0746_),
    .Z(_0460_));
 MUX2_X1 _2893_ (.A(\mem[6][21] ),
    .B(_0647_),
    .S(_0746_),
    .Z(_0461_));
 MUX2_X1 _2894_ (.A(\mem[6][22] ),
    .B(_0649_),
    .S(_0746_),
    .Z(_0462_));
 MUX2_X1 _2895_ (.A(\mem[6][23] ),
    .B(_0651_),
    .S(_0746_),
    .Z(_0463_));
 MUX2_X1 _2896_ (.A(\mem[6][24] ),
    .B(_0653_),
    .S(_0746_),
    .Z(_0464_));
 MUX2_X1 _2897_ (.A(\mem[6][25] ),
    .B(_0655_),
    .S(_0746_),
    .Z(_0465_));
 MUX2_X1 _2898_ (.A(\mem[6][26] ),
    .B(_0657_),
    .S(_0746_),
    .Z(_0466_));
 MUX2_X1 _2899_ (.A(\mem[6][27] ),
    .B(_0659_),
    .S(_0746_),
    .Z(_0467_));
 BUF_X4 _2900_ (.A(_0744_),
    .Z(_0747_));
 MUX2_X1 _2901_ (.A(\mem[6][28] ),
    .B(_0661_),
    .S(_0747_),
    .Z(_0468_));
 MUX2_X1 _2902_ (.A(\mem[6][29] ),
    .B(_0664_),
    .S(_0747_),
    .Z(_0469_));
 MUX2_X1 _2903_ (.A(\mem[6][2] ),
    .B(_0666_),
    .S(_0747_),
    .Z(_0470_));
 MUX2_X1 _2904_ (.A(\mem[6][30] ),
    .B(_0668_),
    .S(_0747_),
    .Z(_0471_));
 MUX2_X1 _2905_ (.A(\mem[6][31] ),
    .B(_0670_),
    .S(_0747_),
    .Z(_0472_));
 MUX2_X1 _2906_ (.A(\mem[6][3] ),
    .B(_0672_),
    .S(_0747_),
    .Z(_0473_));
 MUX2_X1 _2907_ (.A(\mem[6][4] ),
    .B(_0674_),
    .S(_0747_),
    .Z(_0474_));
 MUX2_X1 _2908_ (.A(\mem[6][5] ),
    .B(_0676_),
    .S(_0747_),
    .Z(_0475_));
 MUX2_X1 _2909_ (.A(\mem[6][6] ),
    .B(_0678_),
    .S(_0747_),
    .Z(_0476_));
 MUX2_X1 _2910_ (.A(\mem[6][7] ),
    .B(_0680_),
    .S(_0747_),
    .Z(_0477_));
 MUX2_X1 _2911_ (.A(\mem[6][8] ),
    .B(_0682_),
    .S(_0744_),
    .Z(_0478_));
 MUX2_X1 _2912_ (.A(\mem[6][9] ),
    .B(_0684_),
    .S(_0744_),
    .Z(_0479_));
 AND2_X1 _2913_ (.A1(_0693_),
    .A2(_0732_),
    .ZN(_0748_));
 BUF_X2 _2914_ (.A(_0748_),
    .Z(_0749_));
 BUF_X4 _2915_ (.A(_0749_),
    .Z(_0750_));
 MUX2_X1 _2916_ (.A(\mem[7][0] ),
    .B(_0611_),
    .S(_0750_),
    .Z(_0480_));
 MUX2_X1 _2917_ (.A(\mem[7][10] ),
    .B(_0622_),
    .S(_0750_),
    .Z(_0481_));
 MUX2_X1 _2918_ (.A(\mem[7][11] ),
    .B(_0624_),
    .S(_0750_),
    .Z(_0482_));
 MUX2_X1 _2919_ (.A(\mem[7][12] ),
    .B(_0626_),
    .S(_0750_),
    .Z(_0483_));
 MUX2_X1 _2920_ (.A(\mem[7][13] ),
    .B(_0628_),
    .S(_0750_),
    .Z(_0484_));
 MUX2_X1 _2921_ (.A(\mem[7][14] ),
    .B(_0630_),
    .S(_0750_),
    .Z(_0485_));
 MUX2_X1 _2922_ (.A(\mem[7][15] ),
    .B(_0632_),
    .S(_0750_),
    .Z(_0486_));
 MUX2_X1 _2923_ (.A(\mem[7][16] ),
    .B(_0634_),
    .S(_0750_),
    .Z(_0487_));
 MUX2_X1 _2924_ (.A(\mem[7][17] ),
    .B(_0636_),
    .S(_0750_),
    .Z(_0488_));
 MUX2_X1 _2925_ (.A(\mem[7][18] ),
    .B(_0638_),
    .S(_0750_),
    .Z(_0489_));
 BUF_X4 _2926_ (.A(_0749_),
    .Z(_0751_));
 MUX2_X1 _2927_ (.A(\mem[7][19] ),
    .B(_0640_),
    .S(_0751_),
    .Z(_0490_));
 MUX2_X1 _2928_ (.A(\mem[7][1] ),
    .B(_0643_),
    .S(_0751_),
    .Z(_0491_));
 MUX2_X1 _2929_ (.A(\mem[7][20] ),
    .B(_0645_),
    .S(_0751_),
    .Z(_0492_));
 MUX2_X1 _2930_ (.A(\mem[7][21] ),
    .B(_0647_),
    .S(_0751_),
    .Z(_0493_));
 MUX2_X1 _2931_ (.A(\mem[7][22] ),
    .B(_0649_),
    .S(_0751_),
    .Z(_0494_));
 MUX2_X1 _2932_ (.A(\mem[7][23] ),
    .B(_0651_),
    .S(_0751_),
    .Z(_0495_));
 MUX2_X1 _2933_ (.A(\mem[7][24] ),
    .B(_0653_),
    .S(_0751_),
    .Z(_0496_));
 MUX2_X1 _2934_ (.A(\mem[7][25] ),
    .B(_0655_),
    .S(_0751_),
    .Z(_0497_));
 MUX2_X1 _2935_ (.A(\mem[7][26] ),
    .B(_0657_),
    .S(_0751_),
    .Z(_0498_));
 MUX2_X1 _2936_ (.A(\mem[7][27] ),
    .B(_0659_),
    .S(_0751_),
    .Z(_0499_));
 BUF_X4 _2937_ (.A(_0749_),
    .Z(_0752_));
 MUX2_X1 _2938_ (.A(\mem[7][28] ),
    .B(_0661_),
    .S(_0752_),
    .Z(_0500_));
 MUX2_X1 _2939_ (.A(\mem[7][29] ),
    .B(_0664_),
    .S(_0752_),
    .Z(_0501_));
 MUX2_X1 _2940_ (.A(\mem[7][2] ),
    .B(_0666_),
    .S(_0752_),
    .Z(_0502_));
 MUX2_X1 _2941_ (.A(\mem[7][30] ),
    .B(_0668_),
    .S(_0752_),
    .Z(_0503_));
 MUX2_X1 _2942_ (.A(\mem[7][31] ),
    .B(_0670_),
    .S(_0752_),
    .Z(_0504_));
 MUX2_X1 _2943_ (.A(\mem[7][3] ),
    .B(_0672_),
    .S(_0752_),
    .Z(_0505_));
 MUX2_X1 _2944_ (.A(\mem[7][4] ),
    .B(_0674_),
    .S(_0752_),
    .Z(_0506_));
 MUX2_X1 _2945_ (.A(\mem[7][5] ),
    .B(_0676_),
    .S(_0752_),
    .Z(_0507_));
 MUX2_X1 _2946_ (.A(\mem[7][6] ),
    .B(_0678_),
    .S(_0752_),
    .Z(_0508_));
 MUX2_X1 _2947_ (.A(\mem[7][7] ),
    .B(_0680_),
    .S(_0752_),
    .Z(_0509_));
 MUX2_X1 _2948_ (.A(\mem[7][8] ),
    .B(_0682_),
    .S(_0749_),
    .Z(_0510_));
 MUX2_X1 _2949_ (.A(\mem[7][9] ),
    .B(_0684_),
    .S(_0749_),
    .Z(_0511_));
 NAND2_X4 _2950_ (.A1(_0612_),
    .A2(_0688_),
    .ZN(_0753_));
 BUF_X4 _2951_ (.A(_0753_),
    .Z(_0754_));
 MUX2_X1 _2952_ (.A(_0610_),
    .B(\mem[8][0] ),
    .S(_0754_),
    .Z(_0512_));
 MUX2_X1 _2953_ (.A(_0621_),
    .B(\mem[8][10] ),
    .S(_0754_),
    .Z(_0513_));
 MUX2_X1 _2954_ (.A(_0623_),
    .B(\mem[8][11] ),
    .S(_0754_),
    .Z(_0514_));
 MUX2_X1 _2955_ (.A(_0625_),
    .B(\mem[8][12] ),
    .S(_0754_),
    .Z(_0515_));
 MUX2_X1 _2956_ (.A(_0627_),
    .B(\mem[8][13] ),
    .S(_0754_),
    .Z(_0516_));
 MUX2_X1 _2957_ (.A(_0629_),
    .B(\mem[8][14] ),
    .S(_0754_),
    .Z(_0517_));
 MUX2_X1 _2958_ (.A(_0631_),
    .B(\mem[8][15] ),
    .S(_0754_),
    .Z(_0518_));
 MUX2_X1 _2959_ (.A(_0633_),
    .B(\mem[8][16] ),
    .S(_0754_),
    .Z(_0519_));
 MUX2_X1 _2960_ (.A(_0635_),
    .B(\mem[8][17] ),
    .S(_0754_),
    .Z(_0520_));
 MUX2_X1 _2961_ (.A(_0637_),
    .B(\mem[8][18] ),
    .S(_0754_),
    .Z(_0521_));
 BUF_X4 _2962_ (.A(_0753_),
    .Z(_0755_));
 MUX2_X1 _2963_ (.A(_0639_),
    .B(\mem[8][19] ),
    .S(_0755_),
    .Z(_0522_));
 MUX2_X1 _2964_ (.A(_0642_),
    .B(\mem[8][1] ),
    .S(_0755_),
    .Z(_0523_));
 MUX2_X1 _2965_ (.A(_0644_),
    .B(\mem[8][20] ),
    .S(_0755_),
    .Z(_0524_));
 MUX2_X1 _2966_ (.A(_0646_),
    .B(\mem[8][21] ),
    .S(_0755_),
    .Z(_0525_));
 MUX2_X1 _2967_ (.A(_0648_),
    .B(\mem[8][22] ),
    .S(_0755_),
    .Z(_0526_));
 MUX2_X1 _2968_ (.A(_0650_),
    .B(\mem[8][23] ),
    .S(_0755_),
    .Z(_0527_));
 MUX2_X1 _2969_ (.A(_0652_),
    .B(\mem[8][24] ),
    .S(_0755_),
    .Z(_0528_));
 MUX2_X1 _2970_ (.A(_0654_),
    .B(\mem[8][25] ),
    .S(_0755_),
    .Z(_0529_));
 MUX2_X1 _2971_ (.A(_0656_),
    .B(\mem[8][26] ),
    .S(_0755_),
    .Z(_0530_));
 MUX2_X1 _2972_ (.A(_0658_),
    .B(\mem[8][27] ),
    .S(_0755_),
    .Z(_0531_));
 CLKBUF_X3 _2973_ (.A(_0753_),
    .Z(_0756_));
 MUX2_X1 _2974_ (.A(_0660_),
    .B(\mem[8][28] ),
    .S(_0756_),
    .Z(_0532_));
 MUX2_X1 _2975_ (.A(_0663_),
    .B(\mem[8][29] ),
    .S(_0756_),
    .Z(_0533_));
 MUX2_X1 _2976_ (.A(_0665_),
    .B(\mem[8][2] ),
    .S(_0756_),
    .Z(_0534_));
 MUX2_X1 _2977_ (.A(_0667_),
    .B(\mem[8][30] ),
    .S(_0756_),
    .Z(_0535_));
 MUX2_X1 _2978_ (.A(_0669_),
    .B(\mem[8][31] ),
    .S(_0756_),
    .Z(_0536_));
 MUX2_X1 _2979_ (.A(_0671_),
    .B(\mem[8][3] ),
    .S(_0756_),
    .Z(_0537_));
 MUX2_X1 _2980_ (.A(_0673_),
    .B(\mem[8][4] ),
    .S(_0756_),
    .Z(_0538_));
 MUX2_X1 _2981_ (.A(_0675_),
    .B(\mem[8][5] ),
    .S(_0756_),
    .Z(_0539_));
 MUX2_X1 _2982_ (.A(_0677_),
    .B(\mem[8][6] ),
    .S(_0756_),
    .Z(_0540_));
 MUX2_X1 _2983_ (.A(_0679_),
    .B(\mem[8][7] ),
    .S(_0756_),
    .Z(_0541_));
 MUX2_X1 _2984_ (.A(_0681_),
    .B(\mem[8][8] ),
    .S(_0753_),
    .Z(_0542_));
 MUX2_X1 _2985_ (.A(_0683_),
    .B(\mem[8][9] ),
    .S(_0753_),
    .Z(_0543_));
 NAND2_X4 _2986_ (.A1(_0704_),
    .A2(_0688_),
    .ZN(_0757_));
 BUF_X4 _2987_ (.A(_0757_),
    .Z(_0758_));
 MUX2_X1 _2988_ (.A(_0610_),
    .B(\mem[9][0] ),
    .S(_0758_),
    .Z(_0544_));
 MUX2_X1 _2989_ (.A(_0621_),
    .B(\mem[9][10] ),
    .S(_0758_),
    .Z(_0545_));
 MUX2_X1 _2990_ (.A(_0623_),
    .B(\mem[9][11] ),
    .S(_0758_),
    .Z(_0546_));
 MUX2_X1 _2991_ (.A(_0625_),
    .B(\mem[9][12] ),
    .S(_0758_),
    .Z(_0547_));
 MUX2_X1 _2992_ (.A(_0627_),
    .B(\mem[9][13] ),
    .S(_0758_),
    .Z(_0548_));
 MUX2_X1 _2993_ (.A(_0629_),
    .B(\mem[9][14] ),
    .S(_0758_),
    .Z(_0549_));
 MUX2_X1 _2994_ (.A(_0631_),
    .B(\mem[9][15] ),
    .S(_0758_),
    .Z(_0550_));
 MUX2_X1 _2995_ (.A(_0633_),
    .B(\mem[9][16] ),
    .S(_0758_),
    .Z(_0551_));
 MUX2_X1 _2996_ (.A(_0635_),
    .B(\mem[9][17] ),
    .S(_0758_),
    .Z(_0552_));
 MUX2_X1 _2997_ (.A(_0637_),
    .B(\mem[9][18] ),
    .S(_0758_),
    .Z(_0553_));
 BUF_X4 _2998_ (.A(_0757_),
    .Z(_0759_));
 MUX2_X1 _2999_ (.A(_0639_),
    .B(\mem[9][19] ),
    .S(_0759_),
    .Z(_0554_));
 MUX2_X1 _3000_ (.A(_0642_),
    .B(\mem[9][1] ),
    .S(_0759_),
    .Z(_0555_));
 MUX2_X1 _3001_ (.A(_0644_),
    .B(\mem[9][20] ),
    .S(_0759_),
    .Z(_0556_));
 MUX2_X1 _3002_ (.A(_0646_),
    .B(\mem[9][21] ),
    .S(_0759_),
    .Z(_0557_));
 MUX2_X1 _3003_ (.A(_0648_),
    .B(\mem[9][22] ),
    .S(_0759_),
    .Z(_0558_));
 MUX2_X1 _3004_ (.A(_0650_),
    .B(\mem[9][23] ),
    .S(_0759_),
    .Z(_0559_));
 MUX2_X1 _3005_ (.A(_0652_),
    .B(\mem[9][24] ),
    .S(_0759_),
    .Z(_0560_));
 MUX2_X1 _3006_ (.A(_0654_),
    .B(\mem[9][25] ),
    .S(_0759_),
    .Z(_0561_));
 MUX2_X1 _3007_ (.A(_0656_),
    .B(\mem[9][26] ),
    .S(_0759_),
    .Z(_0562_));
 MUX2_X1 _3008_ (.A(_0658_),
    .B(\mem[9][27] ),
    .S(_0759_),
    .Z(_0563_));
 CLKBUF_X3 _3009_ (.A(_0757_),
    .Z(_0760_));
 MUX2_X1 _3010_ (.A(_0660_),
    .B(\mem[9][28] ),
    .S(_0760_),
    .Z(_0564_));
 MUX2_X1 _3011_ (.A(_0663_),
    .B(\mem[9][29] ),
    .S(_0760_),
    .Z(_0565_));
 MUX2_X1 _3012_ (.A(_0665_),
    .B(\mem[9][2] ),
    .S(_0760_),
    .Z(_0566_));
 MUX2_X1 _3013_ (.A(_0667_),
    .B(\mem[9][30] ),
    .S(_0760_),
    .Z(_0567_));
 MUX2_X1 _3014_ (.A(_0669_),
    .B(\mem[9][31] ),
    .S(_0760_),
    .Z(_0568_));
 MUX2_X1 _3015_ (.A(_0671_),
    .B(\mem[9][3] ),
    .S(_0760_),
    .Z(_0569_));
 MUX2_X1 _3016_ (.A(_0673_),
    .B(\mem[9][4] ),
    .S(_0760_),
    .Z(_0570_));
 MUX2_X1 _3017_ (.A(_0675_),
    .B(\mem[9][5] ),
    .S(_0760_),
    .Z(_0571_));
 MUX2_X1 _3018_ (.A(_0677_),
    .B(\mem[9][6] ),
    .S(_0760_),
    .Z(_0572_));
 MUX2_X1 _3019_ (.A(_0679_),
    .B(\mem[9][7] ),
    .S(_0760_),
    .Z(_0573_));
 MUX2_X1 _3020_ (.A(_0681_),
    .B(\mem[9][8] ),
    .S(_0757_),
    .Z(_0574_));
 MUX2_X1 _3021_ (.A(_0683_),
    .B(\mem[9][9] ),
    .S(_0757_),
    .Z(_0575_));
 CLKBUF_X3 _3022_ (.A(rst_n),
    .Z(_0761_));
 INV_X2 _3023_ (.A(_0761_),
    .ZN(_0762_));
 CLKBUF_X3 _3024_ (.A(_0762_),
    .Z(_0763_));
 NOR2_X1 _3025_ (.A1(\rd_ptr[0] ),
    .A2(_0763_),
    .ZN(_0764_));
 AND2_X1 _3026_ (.A1(\rd_ptr[0] ),
    .A2(_0761_),
    .ZN(_0765_));
 OAI21_X2 _3027_ (.A(_0608_),
    .B1(_0595_),
    .B2(_0605_),
    .ZN(_0766_));
 MUX2_X1 _3028_ (.A(_0764_),
    .B(_0765_),
    .S(_0766_),
    .Z(_0010_));
 BUF_X2 _3029_ (.A(_0761_),
    .Z(_0767_));
 AND2_X1 _3030_ (.A1(_0007_),
    .A2(_0767_),
    .ZN(_0768_));
 CLKBUF_X3 _3031_ (.A(_0761_),
    .Z(_0769_));
 AND2_X1 _3032_ (.A1(\rd_ptr[1] ),
    .A2(_0769_),
    .ZN(_0770_));
 MUX2_X1 _3033_ (.A(_0768_),
    .B(_0770_),
    .S(_0766_),
    .Z(_0011_));
 AND2_X1 _3034_ (.A1(\rd_ptr[2] ),
    .A2(_0767_),
    .ZN(_0771_));
 BUF_X4 _3035_ (.A(_0762_),
    .Z(_0772_));
 NOR2_X1 _3036_ (.A1(\rd_ptr[2] ),
    .A2(_0772_),
    .ZN(_0773_));
 NAND2_X1 _3037_ (.A1(_0608_),
    .A2(_2310_),
    .ZN(_0774_));
 AOI21_X1 _3038_ (.A(_0774_),
    .B1(_0602_),
    .B2(_0593_),
    .ZN(_0775_));
 MUX2_X1 _3039_ (.A(_0771_),
    .B(_0773_),
    .S(_0775_),
    .Z(_0012_));
 AND2_X1 _3040_ (.A1(\rd_ptr[3] ),
    .A2(_0767_),
    .ZN(_0776_));
 NOR2_X1 _3041_ (.A1(\rd_ptr[3] ),
    .A2(_0772_),
    .ZN(_0777_));
 NAND4_X1 _3042_ (.A1(_0608_),
    .A2(\rd_ptr[0] ),
    .A3(\rd_ptr[2] ),
    .A4(\rd_ptr[1] ),
    .ZN(_0778_));
 AOI21_X1 _3043_ (.A(_0778_),
    .B1(_0602_),
    .B2(_0593_),
    .ZN(_0779_));
 MUX2_X1 _3044_ (.A(_0776_),
    .B(_0777_),
    .S(_0779_),
    .Z(_0013_));
 AND2_X1 _3045_ (.A1(_0008_),
    .A2(_0767_),
    .ZN(_0780_));
 AND2_X1 _3046_ (.A1(net10),
    .A2(_0769_),
    .ZN(_0781_));
 MUX2_X1 _3047_ (.A(_0780_),
    .B(_0781_),
    .S(_0609_),
    .Z(_0014_));
 BUF_X1 _3048_ (.A(net11),
    .Z(_0782_));
 NOR2_X1 _3049_ (.A1(_0782_),
    .A2(_0763_),
    .ZN(_0783_));
 AND2_X1 _3050_ (.A1(_0782_),
    .A2(_0769_),
    .ZN(_0784_));
 INV_X1 _3051_ (.A(net25),
    .ZN(_0785_));
 CLKBUF_X2 _3052_ (.A(net21),
    .Z(_0786_));
 BUF_X1 _3053_ (.A(net22),
    .Z(_0787_));
 NAND4_X2 _3054_ (.A1(_0786_),
    .A2(_0787_),
    .A3(net23),
    .A4(net24),
    .ZN(_0788_));
 NOR2_X1 _3055_ (.A1(_0785_),
    .A2(_0788_),
    .ZN(_0789_));
 AND2_X1 _3056_ (.A1(_0608_),
    .A2(net18),
    .ZN(_0790_));
 BUF_X2 _3057_ (.A(_0790_),
    .Z(_0791_));
 AND3_X1 _3058_ (.A1(_2311_),
    .A2(net19),
    .A3(net20),
    .ZN(_0792_));
 AND2_X1 _3059_ (.A1(_0791_),
    .A2(_0792_),
    .ZN(_0793_));
 NAND4_X1 _3060_ (.A1(_0593_),
    .A2(_0602_),
    .A3(_0789_),
    .A4(_0793_),
    .ZN(_0794_));
 MUX2_X1 _3061_ (.A(_0783_),
    .B(_0784_),
    .S(_0794_),
    .Z(_0015_));
 AND2_X1 _3062_ (.A1(net12),
    .A2(_0767_),
    .ZN(_0795_));
 NOR2_X1 _3063_ (.A1(net12),
    .A2(_0772_),
    .ZN(_0796_));
 BUF_X4 _3064_ (.A(_0595_),
    .Z(_0797_));
 BUF_X8 _3065_ (.A(_0605_),
    .Z(_0798_));
 AND4_X1 _3066_ (.A1(net17),
    .A2(net10),
    .A3(net19),
    .A4(net20),
    .ZN(_0799_));
 NAND4_X1 _3067_ (.A1(_0782_),
    .A2(_0789_),
    .A3(_0791_),
    .A4(_0799_),
    .ZN(_0800_));
 NOR3_X1 _3068_ (.A1(_0797_),
    .A2(_0798_),
    .A3(_0800_),
    .ZN(_0801_));
 MUX2_X1 _3069_ (.A(_0795_),
    .B(_0796_),
    .S(_0801_),
    .Z(_0016_));
 AND2_X1 _3070_ (.A1(net13),
    .A2(_0767_),
    .ZN(_0802_));
 NOR2_X1 _3071_ (.A1(net13),
    .A2(_0772_),
    .ZN(_0803_));
 NAND4_X1 _3072_ (.A1(_0782_),
    .A2(net12),
    .A3(_0789_),
    .A4(_0793_),
    .ZN(_0804_));
 NOR3_X1 _3073_ (.A1(_0797_),
    .A2(_0798_),
    .A3(_0804_),
    .ZN(_0805_));
 MUX2_X1 _3074_ (.A(_0802_),
    .B(_0803_),
    .S(_0805_),
    .Z(_0017_));
 NOR2_X1 _3075_ (.A1(net14),
    .A2(_0763_),
    .ZN(_0806_));
 AND2_X1 _3076_ (.A1(net14),
    .A2(_0769_),
    .ZN(_0807_));
 NAND2_X1 _3077_ (.A1(_0791_),
    .A2(_0799_),
    .ZN(_0808_));
 INV_X1 _3078_ (.A(_0808_),
    .ZN(_0809_));
 NAND4_X1 _3079_ (.A1(net25),
    .A2(_0782_),
    .A3(net12),
    .A4(net13),
    .ZN(_0810_));
 NOR2_X1 _3080_ (.A1(_0788_),
    .A2(_0810_),
    .ZN(_0811_));
 NAND4_X1 _3081_ (.A1(_0593_),
    .A2(_0602_),
    .A3(_0809_),
    .A4(_0811_),
    .ZN(_0812_));
 MUX2_X1 _3082_ (.A(_0806_),
    .B(_0807_),
    .S(_0812_),
    .Z(_0018_));
 AND2_X1 _3083_ (.A1(net15),
    .A2(_0767_),
    .ZN(_0813_));
 NOR2_X1 _3084_ (.A1(net15),
    .A2(_0772_),
    .ZN(_0814_));
 BUF_X4 _3085_ (.A(_0605_),
    .Z(_0815_));
 NAND3_X1 _3086_ (.A1(net14),
    .A2(_0793_),
    .A3(_0811_),
    .ZN(_0816_));
 NOR3_X1 _3087_ (.A1(_0797_),
    .A2(_0815_),
    .A3(_0816_),
    .ZN(_0817_));
 MUX2_X1 _3088_ (.A(_0813_),
    .B(_0814_),
    .S(_0817_),
    .Z(_0019_));
 AND2_X1 _3089_ (.A1(net16),
    .A2(_0767_),
    .ZN(_0818_));
 NOR2_X1 _3090_ (.A1(net16),
    .A2(_0772_),
    .ZN(_0819_));
 AND3_X1 _3091_ (.A1(net15),
    .A2(_0791_),
    .A3(_0799_),
    .ZN(_0820_));
 NAND3_X1 _3092_ (.A1(net14),
    .A2(_0811_),
    .A3(_0820_),
    .ZN(_0821_));
 NOR3_X1 _3093_ (.A1(_0797_),
    .A2(_0815_),
    .A3(_0821_),
    .ZN(_0822_));
 MUX2_X1 _3094_ (.A(_0818_),
    .B(_0819_),
    .S(_0822_),
    .Z(_0020_));
 AND2_X1 _3095_ (.A1(_0009_),
    .A2(_0767_),
    .ZN(_0823_));
 AND2_X1 _3096_ (.A1(net17),
    .A2(_0769_),
    .ZN(_0824_));
 MUX2_X1 _3097_ (.A(_0823_),
    .B(_0824_),
    .S(_0609_),
    .Z(_0021_));
 NOR2_X1 _3098_ (.A1(net18),
    .A2(_0763_),
    .ZN(_0825_));
 AND2_X1 _3099_ (.A1(net18),
    .A2(_0769_),
    .ZN(_0826_));
 NAND4_X1 _3100_ (.A1(_0608_),
    .A2(_2311_),
    .A3(_0593_),
    .A4(_0601_),
    .ZN(_0827_));
 MUX2_X1 _3101_ (.A(_0825_),
    .B(_0826_),
    .S(_0827_),
    .Z(_0022_));
 BUF_X2 _3102_ (.A(_0761_),
    .Z(_0828_));
 AND2_X1 _3103_ (.A1(net19),
    .A2(_0828_),
    .ZN(_0829_));
 CLKBUF_X3 _3104_ (.A(_0762_),
    .Z(_0830_));
 NOR2_X1 _3105_ (.A1(net19),
    .A2(_0830_),
    .ZN(_0831_));
 NAND3_X1 _3106_ (.A1(net17),
    .A2(net10),
    .A3(_0791_),
    .ZN(_0832_));
 NOR3_X1 _3107_ (.A1(_0797_),
    .A2(_0815_),
    .A3(_0832_),
    .ZN(_0833_));
 MUX2_X1 _3108_ (.A(_0829_),
    .B(_0831_),
    .S(_0833_),
    .Z(_0023_));
 AND2_X1 _3109_ (.A1(net20),
    .A2(_0828_),
    .ZN(_0834_));
 NOR2_X1 _3110_ (.A1(net20),
    .A2(_0830_),
    .ZN(_0835_));
 NAND3_X1 _3111_ (.A1(_2311_),
    .A2(net19),
    .A3(_0791_),
    .ZN(_0836_));
 NOR3_X1 _3112_ (.A1(_0797_),
    .A2(_0815_),
    .A3(_0836_),
    .ZN(_0837_));
 MUX2_X1 _3113_ (.A(_0834_),
    .B(_0835_),
    .S(_0837_),
    .Z(_0024_));
 AND2_X1 _3114_ (.A1(_0786_),
    .A2(_0828_),
    .ZN(_0838_));
 NOR2_X1 _3115_ (.A1(_0786_),
    .A2(_0830_),
    .ZN(_0839_));
 NOR3_X1 _3116_ (.A1(_0797_),
    .A2(_0798_),
    .A3(_0808_),
    .ZN(_0840_));
 MUX2_X1 _3117_ (.A(_0838_),
    .B(_0839_),
    .S(_0840_),
    .Z(_0025_));
 AND2_X1 _3118_ (.A1(_0787_),
    .A2(_0828_),
    .ZN(_0841_));
 NOR2_X1 _3119_ (.A1(_0787_),
    .A2(_0830_),
    .ZN(_0842_));
 NAND3_X1 _3120_ (.A1(_0786_),
    .A2(_0791_),
    .A3(_0792_),
    .ZN(_0843_));
 NOR3_X1 _3121_ (.A1(_0797_),
    .A2(_0815_),
    .A3(_0843_),
    .ZN(_0844_));
 MUX2_X1 _3122_ (.A(_0841_),
    .B(_0842_),
    .S(_0844_),
    .Z(_0026_));
 AND2_X1 _3123_ (.A1(net23),
    .A2(_0828_),
    .ZN(_0845_));
 NOR2_X1 _3124_ (.A1(net23),
    .A2(_0830_),
    .ZN(_0846_));
 NAND4_X1 _3125_ (.A1(_0786_),
    .A2(_0787_),
    .A3(_0791_),
    .A4(_0799_),
    .ZN(_0847_));
 NOR3_X1 _3126_ (.A1(_0797_),
    .A2(_0815_),
    .A3(_0847_),
    .ZN(_0848_));
 MUX2_X1 _3127_ (.A(_0845_),
    .B(_0846_),
    .S(_0848_),
    .Z(_0027_));
 NOR2_X1 _3128_ (.A1(net24),
    .A2(_0763_),
    .ZN(_0849_));
 AND2_X1 _3129_ (.A1(net24),
    .A2(_0769_),
    .ZN(_0850_));
 AND3_X1 _3130_ (.A1(_0786_),
    .A2(_0787_),
    .A3(net23),
    .ZN(_0851_));
 NAND4_X1 _3131_ (.A1(_0593_),
    .A2(_0602_),
    .A3(_0851_),
    .A4(_0793_),
    .ZN(_0852_));
 MUX2_X1 _3132_ (.A(_0849_),
    .B(_0850_),
    .S(_0852_),
    .Z(_0028_));
 NOR2_X1 _3133_ (.A1(_0785_),
    .A2(_0763_),
    .ZN(_0853_));
 NOR2_X1 _3134_ (.A1(net25),
    .A2(_0830_),
    .ZN(_0854_));
 NOR4_X1 _3135_ (.A1(_0595_),
    .A2(_0815_),
    .A3(_0788_),
    .A4(_0808_),
    .ZN(_0855_));
 MUX2_X1 _3136_ (.A(_0853_),
    .B(_0854_),
    .S(_0855_),
    .Z(_0029_));
 CLKBUF_X3 _3137_ (.A(_0763_),
    .Z(_0856_));
 INV_X1 _3138_ (.A(net1),
    .ZN(_0857_));
 NAND2_X1 _3139_ (.A1(net26),
    .A2(_0857_),
    .ZN(_0858_));
 AOI21_X1 _3140_ (.A(_0856_),
    .B1(_0609_),
    .B2(_0858_),
    .ZN(_0030_));
 INV_X2 _3141_ (.A(_0608_),
    .ZN(_0859_));
 NOR2_X4 _3142_ (.A1(_0859_),
    .A2(_0762_),
    .ZN(_0860_));
 CLKBUF_X3 _3143_ (.A(_0860_),
    .Z(_0861_));
 CLKBUF_X2 _3144_ (.A(_0000_),
    .Z(_0862_));
 BUF_X4 _3145_ (.A(_0862_),
    .Z(_0863_));
 CLKBUF_X3 _3146_ (.A(_0863_),
    .Z(_0864_));
 BUF_X2 _3147_ (.A(_0002_),
    .Z(_0865_));
 BUF_X4 _3148_ (.A(_0865_),
    .Z(_0866_));
 BUF_X4 _3149_ (.A(_0866_),
    .Z(_0867_));
 MUX2_X1 _3150_ (.A(\mem[2][0] ),
    .B(\mem[6][0] ),
    .S(_0867_),
    .Z(_0868_));
 NOR2_X1 _3151_ (.A1(_0864_),
    .A2(_0868_),
    .ZN(_0869_));
 INV_X1 _3152_ (.A(_0862_),
    .ZN(_0870_));
 BUF_X4 _3153_ (.A(_0870_),
    .Z(_0871_));
 BUF_X4 _3154_ (.A(_0871_),
    .Z(_0872_));
 BUF_X4 _3155_ (.A(_0866_),
    .Z(_0873_));
 MUX2_X1 _3156_ (.A(\mem[3][0] ),
    .B(\mem[7][0] ),
    .S(_0873_),
    .Z(_0874_));
 NOR2_X1 _3157_ (.A1(_0872_),
    .A2(_0874_),
    .ZN(_0875_));
 INV_X1 _3158_ (.A(_0001_),
    .ZN(_0876_));
 BUF_X2 _3159_ (.A(_0003_),
    .Z(_0877_));
 OR2_X1 _3160_ (.A1(_0876_),
    .A2(_0877_),
    .ZN(_0878_));
 CLKBUF_X2 _3161_ (.A(_0878_),
    .Z(_0879_));
 CLKBUF_X3 _3162_ (.A(_0879_),
    .Z(_0880_));
 NAND2_X2 _3163_ (.A1(_0001_),
    .A2(_0877_),
    .ZN(_0881_));
 BUF_X4 _3164_ (.A(_0865_),
    .Z(_0882_));
 BUF_X4 _3165_ (.A(_0882_),
    .Z(_0883_));
 MUX2_X1 _3166_ (.A(\mem[10][0] ),
    .B(\mem[14][0] ),
    .S(_0883_),
    .Z(_0884_));
 NOR2_X1 _3167_ (.A1(_0863_),
    .A2(_0884_),
    .ZN(_0885_));
 BUF_X4 _3168_ (.A(_0870_),
    .Z(_0886_));
 CLKBUF_X3 _3169_ (.A(_0886_),
    .Z(_0887_));
 MUX2_X1 _3170_ (.A(\mem[11][0] ),
    .B(\mem[15][0] ),
    .S(_0883_),
    .Z(_0888_));
 NOR2_X1 _3171_ (.A1(_0887_),
    .A2(_0888_),
    .ZN(_0889_));
 OAI33_X1 _3172_ (.A1(_0869_),
    .A2(_0875_),
    .A3(_0880_),
    .B1(_0881_),
    .B2(_0885_),
    .B3(_0889_),
    .ZN(_0890_));
 MUX2_X1 _3173_ (.A(\mem[0][0] ),
    .B(\mem[4][0] ),
    .S(_0867_),
    .Z(_0891_));
 NOR2_X1 _3174_ (.A1(_0864_),
    .A2(_0891_),
    .ZN(_0892_));
 BUF_X4 _3175_ (.A(_0886_),
    .Z(_0893_));
 BUF_X4 _3176_ (.A(_0865_),
    .Z(_0894_));
 BUF_X4 _3177_ (.A(_0894_),
    .Z(_0895_));
 MUX2_X1 _3178_ (.A(\mem[1][0] ),
    .B(\mem[5][0] ),
    .S(_0895_),
    .Z(_0896_));
 NOR2_X1 _3179_ (.A1(_0893_),
    .A2(_0896_),
    .ZN(_0897_));
 OR2_X1 _3180_ (.A1(_0001_),
    .A2(_0877_),
    .ZN(_0898_));
 BUF_X2 _3181_ (.A(_0898_),
    .Z(_0899_));
 BUF_X4 _3182_ (.A(_0899_),
    .Z(_0900_));
 NAND2_X4 _3183_ (.A1(_0876_),
    .A2(_0877_),
    .ZN(_0901_));
 MUX2_X1 _3184_ (.A(\mem[8][0] ),
    .B(\mem[12][0] ),
    .S(_0883_),
    .Z(_0902_));
 NOR2_X1 _3185_ (.A1(_0863_),
    .A2(_0902_),
    .ZN(_0903_));
 MUX2_X1 _3186_ (.A(\mem[9][0] ),
    .B(\mem[13][0] ),
    .S(_0866_),
    .Z(_0904_));
 NOR2_X1 _3187_ (.A1(_0871_),
    .A2(_0904_),
    .ZN(_0905_));
 OAI33_X1 _3188_ (.A1(_0892_),
    .A2(_0897_),
    .A3(_0900_),
    .B1(_0901_),
    .B2(_0903_),
    .B3(_0905_),
    .ZN(_0906_));
 OAI221_X1 _3189_ (.A(_0861_),
    .B1(_0890_),
    .B2(_0906_),
    .C1(_0597_),
    .C2(_0798_),
    .ZN(_0907_));
 CLKBUF_X3 _3190_ (.A(_0761_),
    .Z(_0908_));
 NAND2_X1 _3191_ (.A1(\last_valid_data[0] ),
    .A2(_0908_),
    .ZN(_0909_));
 BUF_X8 _3192_ (.A(_0607_),
    .Z(_0910_));
 CLKBUF_X3 _3193_ (.A(_0859_),
    .Z(_0911_));
 NAND2_X1 _3194_ (.A1(_0911_),
    .A2(\last_valid_data[0] ),
    .ZN(_0912_));
 OAI221_X1 _3195_ (.A(_0907_),
    .B1(_0909_),
    .B2(_0910_),
    .C1(_0912_),
    .C2(_0856_),
    .ZN(_0031_));
 BUF_X4 _3196_ (.A(_0901_),
    .Z(_0913_));
 MUX2_X1 _3197_ (.A(\mem[8][10] ),
    .B(\mem[12][10] ),
    .S(_0867_),
    .Z(_0914_));
 NOR2_X1 _3198_ (.A1(_0864_),
    .A2(_0914_),
    .ZN(_0915_));
 MUX2_X1 _3199_ (.A(\mem[9][10] ),
    .B(\mem[13][10] ),
    .S(_0873_),
    .Z(_0916_));
 NOR2_X1 _3200_ (.A1(_0872_),
    .A2(_0916_),
    .ZN(_0917_));
 BUF_X4 _3201_ (.A(_0862_),
    .Z(_0918_));
 BUF_X4 _3202_ (.A(_0918_),
    .Z(_0919_));
 BUF_X4 _3203_ (.A(_0894_),
    .Z(_0920_));
 MUX2_X1 _3204_ (.A(\mem[0][10] ),
    .B(\mem[4][10] ),
    .S(_0920_),
    .Z(_0921_));
 NOR2_X1 _3205_ (.A1(_0919_),
    .A2(_0921_),
    .ZN(_0922_));
 BUF_X4 _3206_ (.A(_0886_),
    .Z(_0923_));
 BUF_X4 _3207_ (.A(_0882_),
    .Z(_0924_));
 MUX2_X1 _3208_ (.A(\mem[1][10] ),
    .B(\mem[5][10] ),
    .S(_0924_),
    .Z(_0925_));
 NOR2_X1 _3209_ (.A1(_0923_),
    .A2(_0925_),
    .ZN(_0926_));
 OAI33_X1 _3210_ (.A1(_0913_),
    .A2(_0915_),
    .A3(_0917_),
    .B1(_0922_),
    .B2(_0926_),
    .B3(_0900_),
    .ZN(_0927_));
 BUF_X4 _3211_ (.A(_0881_),
    .Z(_0928_));
 BUF_X4 _3212_ (.A(_0918_),
    .Z(_0929_));
 MUX2_X1 _3213_ (.A(\mem[10][10] ),
    .B(\mem[14][10] ),
    .S(_0895_),
    .Z(_0930_));
 NOR2_X1 _3214_ (.A1(_0929_),
    .A2(_0930_),
    .ZN(_0931_));
 BUF_X4 _3215_ (.A(_0894_),
    .Z(_0932_));
 MUX2_X1 _3216_ (.A(\mem[11][10] ),
    .B(\mem[15][10] ),
    .S(_0932_),
    .Z(_0933_));
 NOR2_X1 _3217_ (.A1(_0893_),
    .A2(_0933_),
    .ZN(_0934_));
 CLKBUF_X3 _3218_ (.A(_0918_),
    .Z(_0935_));
 BUF_X4 _3219_ (.A(_0882_),
    .Z(_0936_));
 MUX2_X1 _3220_ (.A(\mem[2][10] ),
    .B(\mem[6][10] ),
    .S(_0936_),
    .Z(_0937_));
 NOR2_X1 _3221_ (.A1(_0935_),
    .A2(_0937_),
    .ZN(_0938_));
 MUX2_X1 _3222_ (.A(\mem[3][10] ),
    .B(\mem[7][10] ),
    .S(_0883_),
    .Z(_0939_));
 NOR2_X1 _3223_ (.A1(_0887_),
    .A2(_0939_),
    .ZN(_0940_));
 OAI33_X1 _3224_ (.A1(_0928_),
    .A2(_0931_),
    .A3(_0934_),
    .B1(_0938_),
    .B2(_0940_),
    .B3(_0880_),
    .ZN(_0941_));
 BUF_X2 _3225_ (.A(_0815_),
    .Z(_0942_));
 OAI221_X1 _3226_ (.A(_0861_),
    .B1(_0927_),
    .B2(_0941_),
    .C1(_0942_),
    .C2(_0597_),
    .ZN(_0943_));
 NAND2_X1 _3227_ (.A1(\last_valid_data[10] ),
    .A2(_0908_),
    .ZN(_0944_));
 NAND2_X1 _3228_ (.A1(_0911_),
    .A2(\last_valid_data[10] ),
    .ZN(_0945_));
 OAI221_X1 _3229_ (.A(_0943_),
    .B1(_0944_),
    .B2(_0910_),
    .C1(_0945_),
    .C2(_0856_),
    .ZN(_0032_));
 MUX2_X1 _3230_ (.A(\mem[8][11] ),
    .B(\mem[12][11] ),
    .S(_0867_),
    .Z(_0946_));
 NOR2_X1 _3231_ (.A1(_0864_),
    .A2(_0946_),
    .ZN(_0947_));
 MUX2_X1 _3232_ (.A(\mem[9][11] ),
    .B(\mem[13][11] ),
    .S(_0873_),
    .Z(_0948_));
 NOR2_X1 _3233_ (.A1(_0872_),
    .A2(_0948_),
    .ZN(_0949_));
 MUX2_X1 _3234_ (.A(\mem[0][11] ),
    .B(\mem[4][11] ),
    .S(_0920_),
    .Z(_0950_));
 NOR2_X1 _3235_ (.A1(_0919_),
    .A2(_0950_),
    .ZN(_0951_));
 MUX2_X1 _3236_ (.A(\mem[1][11] ),
    .B(\mem[5][11] ),
    .S(_0924_),
    .Z(_0952_));
 NOR2_X1 _3237_ (.A1(_0923_),
    .A2(_0952_),
    .ZN(_0953_));
 OAI33_X1 _3238_ (.A1(_0913_),
    .A2(_0947_),
    .A3(_0949_),
    .B1(_0951_),
    .B2(_0953_),
    .B3(_0900_),
    .ZN(_0954_));
 MUX2_X1 _3239_ (.A(\mem[10][11] ),
    .B(\mem[14][11] ),
    .S(_0895_),
    .Z(_0955_));
 NOR2_X1 _3240_ (.A1(_0929_),
    .A2(_0955_),
    .ZN(_0956_));
 MUX2_X1 _3241_ (.A(\mem[11][11] ),
    .B(\mem[15][11] ),
    .S(_0932_),
    .Z(_0957_));
 NOR2_X1 _3242_ (.A1(_0893_),
    .A2(_0957_),
    .ZN(_0958_));
 BUF_X4 _3243_ (.A(_0882_),
    .Z(_0959_));
 MUX2_X1 _3244_ (.A(\mem[2][11] ),
    .B(\mem[6][11] ),
    .S(_0959_),
    .Z(_0960_));
 NOR2_X1 _3245_ (.A1(_0935_),
    .A2(_0960_),
    .ZN(_0961_));
 MUX2_X1 _3246_ (.A(\mem[3][11] ),
    .B(\mem[7][11] ),
    .S(_0883_),
    .Z(_0962_));
 NOR2_X1 _3247_ (.A1(_0887_),
    .A2(_0962_),
    .ZN(_0963_));
 OAI33_X1 _3248_ (.A1(_0928_),
    .A2(_0956_),
    .A3(_0958_),
    .B1(_0961_),
    .B2(_0963_),
    .B3(_0880_),
    .ZN(_0964_));
 OAI221_X1 _3249_ (.A(_0861_),
    .B1(_0954_),
    .B2(_0964_),
    .C1(_0942_),
    .C2(_0597_),
    .ZN(_0965_));
 NAND2_X1 _3250_ (.A1(\last_valid_data[11] ),
    .A2(_0908_),
    .ZN(_0966_));
 NAND2_X1 _3251_ (.A1(_0911_),
    .A2(\last_valid_data[11] ),
    .ZN(_0967_));
 OAI221_X1 _3252_ (.A(_0965_),
    .B1(_0966_),
    .B2(_0910_),
    .C1(_0967_),
    .C2(_0856_),
    .ZN(_0033_));
 MUX2_X1 _3253_ (.A(\mem[8][12] ),
    .B(\mem[12][12] ),
    .S(_0867_),
    .Z(_0968_));
 NOR2_X1 _3254_ (.A1(_0864_),
    .A2(_0968_),
    .ZN(_0969_));
 MUX2_X1 _3255_ (.A(\mem[9][12] ),
    .B(\mem[13][12] ),
    .S(_0873_),
    .Z(_0970_));
 NOR2_X1 _3256_ (.A1(_0872_),
    .A2(_0970_),
    .ZN(_0971_));
 MUX2_X1 _3257_ (.A(\mem[0][12] ),
    .B(\mem[4][12] ),
    .S(_0920_),
    .Z(_0972_));
 NOR2_X1 _3258_ (.A1(_0919_),
    .A2(_0972_),
    .ZN(_0973_));
 MUX2_X1 _3259_ (.A(\mem[1][12] ),
    .B(\mem[5][12] ),
    .S(_0924_),
    .Z(_0974_));
 NOR2_X1 _3260_ (.A1(_0923_),
    .A2(_0974_),
    .ZN(_0975_));
 OAI33_X1 _3261_ (.A1(_0913_),
    .A2(_0969_),
    .A3(_0971_),
    .B1(_0973_),
    .B2(_0975_),
    .B3(_0900_),
    .ZN(_0976_));
 MUX2_X1 _3262_ (.A(\mem[10][12] ),
    .B(\mem[14][12] ),
    .S(_0895_),
    .Z(_0977_));
 NOR2_X1 _3263_ (.A1(_0929_),
    .A2(_0977_),
    .ZN(_0978_));
 BUF_X4 _3264_ (.A(_0894_),
    .Z(_0979_));
 MUX2_X1 _3265_ (.A(\mem[11][12] ),
    .B(\mem[15][12] ),
    .S(_0979_),
    .Z(_0980_));
 NOR2_X1 _3266_ (.A1(_0893_),
    .A2(_0980_),
    .ZN(_0981_));
 MUX2_X1 _3267_ (.A(\mem[2][12] ),
    .B(\mem[6][12] ),
    .S(_0959_),
    .Z(_0982_));
 NOR2_X1 _3268_ (.A1(_0935_),
    .A2(_0982_),
    .ZN(_0983_));
 MUX2_X1 _3269_ (.A(\mem[3][12] ),
    .B(\mem[7][12] ),
    .S(_0883_),
    .Z(_0984_));
 NOR2_X1 _3270_ (.A1(_0887_),
    .A2(_0984_),
    .ZN(_0985_));
 OAI33_X1 _3271_ (.A1(_0928_),
    .A2(_0978_),
    .A3(_0981_),
    .B1(_0983_),
    .B2(_0985_),
    .B3(_0880_),
    .ZN(_0986_));
 OAI221_X1 _3272_ (.A(_0861_),
    .B1(_0976_),
    .B2(_0986_),
    .C1(_0942_),
    .C2(_0597_),
    .ZN(_0987_));
 NAND2_X1 _3273_ (.A1(\last_valid_data[12] ),
    .A2(_0908_),
    .ZN(_0988_));
 NAND2_X1 _3274_ (.A1(_0911_),
    .A2(\last_valid_data[12] ),
    .ZN(_0989_));
 OAI221_X1 _3275_ (.A(_0987_),
    .B1(_0988_),
    .B2(_0910_),
    .C1(_0989_),
    .C2(_0856_),
    .ZN(_0034_));
 MUX2_X1 _3276_ (.A(\mem[8][13] ),
    .B(\mem[12][13] ),
    .S(_0867_),
    .Z(_0990_));
 NOR2_X1 _3277_ (.A1(_0864_),
    .A2(_0990_),
    .ZN(_0991_));
 MUX2_X1 _3278_ (.A(\mem[9][13] ),
    .B(\mem[13][13] ),
    .S(_0873_),
    .Z(_0992_));
 NOR2_X1 _3279_ (.A1(_0872_),
    .A2(_0992_),
    .ZN(_0993_));
 BUF_X4 _3280_ (.A(_0894_),
    .Z(_0994_));
 MUX2_X1 _3281_ (.A(\mem[0][13] ),
    .B(\mem[4][13] ),
    .S(_0994_),
    .Z(_0995_));
 NOR2_X1 _3282_ (.A1(_0919_),
    .A2(_0995_),
    .ZN(_0996_));
 MUX2_X1 _3283_ (.A(\mem[1][13] ),
    .B(\mem[5][13] ),
    .S(_0924_),
    .Z(_0997_));
 NOR2_X1 _3284_ (.A1(_0923_),
    .A2(_0997_),
    .ZN(_0998_));
 OAI33_X1 _3285_ (.A1(_0913_),
    .A2(_0991_),
    .A3(_0993_),
    .B1(_0996_),
    .B2(_0998_),
    .B3(_0900_),
    .ZN(_0999_));
 MUX2_X1 _3286_ (.A(\mem[10][13] ),
    .B(\mem[14][13] ),
    .S(_0895_),
    .Z(_1000_));
 NOR2_X1 _3287_ (.A1(_0929_),
    .A2(_1000_),
    .ZN(_1001_));
 MUX2_X1 _3288_ (.A(\mem[11][13] ),
    .B(\mem[15][13] ),
    .S(_0979_),
    .Z(_1002_));
 NOR2_X1 _3289_ (.A1(_0893_),
    .A2(_1002_),
    .ZN(_1003_));
 MUX2_X1 _3290_ (.A(\mem[2][13] ),
    .B(\mem[6][13] ),
    .S(_0959_),
    .Z(_1004_));
 NOR2_X1 _3291_ (.A1(_0935_),
    .A2(_1004_),
    .ZN(_1005_));
 MUX2_X1 _3292_ (.A(\mem[3][13] ),
    .B(\mem[7][13] ),
    .S(_0883_),
    .Z(_1006_));
 NOR2_X1 _3293_ (.A1(_0887_),
    .A2(_1006_),
    .ZN(_1007_));
 OAI33_X1 _3294_ (.A1(_0928_),
    .A2(_1001_),
    .A3(_1003_),
    .B1(_1005_),
    .B2(_1007_),
    .B3(_0880_),
    .ZN(_1008_));
 OAI221_X1 _3295_ (.A(_0861_),
    .B1(_0999_),
    .B2(_1008_),
    .C1(_0942_),
    .C2(_0597_),
    .ZN(_1009_));
 NAND2_X1 _3296_ (.A1(\last_valid_data[13] ),
    .A2(_0908_),
    .ZN(_1010_));
 NAND2_X1 _3297_ (.A1(_0911_),
    .A2(\last_valid_data[13] ),
    .ZN(_1011_));
 OAI221_X1 _3298_ (.A(_1009_),
    .B1(_1010_),
    .B2(_0910_),
    .C1(_1011_),
    .C2(_0856_),
    .ZN(_0035_));
 MUX2_X1 _3299_ (.A(\mem[8][14] ),
    .B(\mem[12][14] ),
    .S(_0867_),
    .Z(_1012_));
 NOR2_X1 _3300_ (.A1(_0864_),
    .A2(_1012_),
    .ZN(_1013_));
 MUX2_X1 _3301_ (.A(\mem[9][14] ),
    .B(\mem[13][14] ),
    .S(_0873_),
    .Z(_1014_));
 NOR2_X1 _3302_ (.A1(_0872_),
    .A2(_1014_),
    .ZN(_1015_));
 MUX2_X1 _3303_ (.A(\mem[0][14] ),
    .B(\mem[4][14] ),
    .S(_0994_),
    .Z(_1016_));
 NOR2_X1 _3304_ (.A1(_0919_),
    .A2(_1016_),
    .ZN(_1017_));
 MUX2_X1 _3305_ (.A(\mem[1][14] ),
    .B(\mem[5][14] ),
    .S(_0924_),
    .Z(_1018_));
 NOR2_X1 _3306_ (.A1(_0923_),
    .A2(_1018_),
    .ZN(_1019_));
 OAI33_X1 _3307_ (.A1(_0913_),
    .A2(_1013_),
    .A3(_1015_),
    .B1(_1017_),
    .B2(_1019_),
    .B3(_0900_),
    .ZN(_1020_));
 BUF_X4 _3308_ (.A(_0894_),
    .Z(_1021_));
 MUX2_X1 _3309_ (.A(\mem[10][14] ),
    .B(\mem[14][14] ),
    .S(_1021_),
    .Z(_1022_));
 NOR2_X1 _3310_ (.A1(_0929_),
    .A2(_1022_),
    .ZN(_1023_));
 MUX2_X1 _3311_ (.A(\mem[11][14] ),
    .B(\mem[15][14] ),
    .S(_0979_),
    .Z(_1024_));
 NOR2_X1 _3312_ (.A1(_0893_),
    .A2(_1024_),
    .ZN(_1025_));
 MUX2_X1 _3313_ (.A(\mem[2][14] ),
    .B(\mem[6][14] ),
    .S(_0959_),
    .Z(_1026_));
 NOR2_X1 _3314_ (.A1(_0935_),
    .A2(_1026_),
    .ZN(_1027_));
 BUF_X4 _3315_ (.A(_0886_),
    .Z(_1028_));
 MUX2_X1 _3316_ (.A(\mem[3][14] ),
    .B(\mem[7][14] ),
    .S(_0883_),
    .Z(_1029_));
 NOR2_X1 _3317_ (.A1(_1028_),
    .A2(_1029_),
    .ZN(_1030_));
 OAI33_X1 _3318_ (.A1(_0928_),
    .A2(_1023_),
    .A3(_1025_),
    .B1(_1027_),
    .B2(_1030_),
    .B3(_0880_),
    .ZN(_1031_));
 CLKBUF_X3 _3319_ (.A(_0595_),
    .Z(_1032_));
 OAI221_X1 _3320_ (.A(_0861_),
    .B1(_1020_),
    .B2(_1031_),
    .C1(_0942_),
    .C2(_1032_),
    .ZN(_1033_));
 NAND2_X1 _3321_ (.A1(\last_valid_data[14] ),
    .A2(_0908_),
    .ZN(_1034_));
 NAND2_X1 _3322_ (.A1(_0911_),
    .A2(\last_valid_data[14] ),
    .ZN(_1035_));
 OAI221_X1 _3323_ (.A(_1033_),
    .B1(_1034_),
    .B2(_0910_),
    .C1(_1035_),
    .C2(_0856_),
    .ZN(_0036_));
 MUX2_X1 _3324_ (.A(\mem[8][15] ),
    .B(\mem[12][15] ),
    .S(_0867_),
    .Z(_1036_));
 NOR2_X1 _3325_ (.A1(_0864_),
    .A2(_1036_),
    .ZN(_1037_));
 MUX2_X1 _3326_ (.A(\mem[9][15] ),
    .B(\mem[13][15] ),
    .S(_0873_),
    .Z(_1038_));
 NOR2_X1 _3327_ (.A1(_0872_),
    .A2(_1038_),
    .ZN(_1039_));
 MUX2_X1 _3328_ (.A(\mem[0][15] ),
    .B(\mem[4][15] ),
    .S(_0994_),
    .Z(_1040_));
 NOR2_X1 _3329_ (.A1(_0919_),
    .A2(_1040_),
    .ZN(_1041_));
 MUX2_X1 _3330_ (.A(\mem[1][15] ),
    .B(\mem[5][15] ),
    .S(_0924_),
    .Z(_1042_));
 NOR2_X1 _3331_ (.A1(_0923_),
    .A2(_1042_),
    .ZN(_1043_));
 OAI33_X1 _3332_ (.A1(_0913_),
    .A2(_1037_),
    .A3(_1039_),
    .B1(_1041_),
    .B2(_1043_),
    .B3(_0900_),
    .ZN(_1044_));
 MUX2_X1 _3333_ (.A(\mem[10][15] ),
    .B(\mem[14][15] ),
    .S(_1021_),
    .Z(_1045_));
 NOR2_X1 _3334_ (.A1(_0929_),
    .A2(_1045_),
    .ZN(_1046_));
 MUX2_X1 _3335_ (.A(\mem[11][15] ),
    .B(\mem[15][15] ),
    .S(_0979_),
    .Z(_1047_));
 NOR2_X1 _3336_ (.A1(_0893_),
    .A2(_1047_),
    .ZN(_1048_));
 BUF_X4 _3337_ (.A(_0918_),
    .Z(_1049_));
 MUX2_X1 _3338_ (.A(\mem[2][15] ),
    .B(\mem[6][15] ),
    .S(_0959_),
    .Z(_1050_));
 NOR2_X1 _3339_ (.A1(_1049_),
    .A2(_1050_),
    .ZN(_1051_));
 MUX2_X1 _3340_ (.A(\mem[3][15] ),
    .B(\mem[7][15] ),
    .S(_0883_),
    .Z(_1052_));
 NOR2_X1 _3341_ (.A1(_1028_),
    .A2(_1052_),
    .ZN(_1053_));
 OAI33_X1 _3342_ (.A1(_0928_),
    .A2(_1046_),
    .A3(_1048_),
    .B1(_1051_),
    .B2(_1053_),
    .B3(_0880_),
    .ZN(_1054_));
 OAI221_X1 _3343_ (.A(_0861_),
    .B1(_1044_),
    .B2(_1054_),
    .C1(_0942_),
    .C2(_1032_),
    .ZN(_1055_));
 NAND2_X1 _3344_ (.A1(\last_valid_data[15] ),
    .A2(_0908_),
    .ZN(_1056_));
 NAND2_X1 _3345_ (.A1(_0911_),
    .A2(\last_valid_data[15] ),
    .ZN(_1057_));
 OAI221_X1 _3346_ (.A(_1055_),
    .B1(_1056_),
    .B2(_0910_),
    .C1(_1057_),
    .C2(_0856_),
    .ZN(_0037_));
 MUX2_X1 _3347_ (.A(\mem[8][16] ),
    .B(\mem[12][16] ),
    .S(_0867_),
    .Z(_1058_));
 NOR2_X1 _3348_ (.A1(_0864_),
    .A2(_1058_),
    .ZN(_1059_));
 BUF_X4 _3349_ (.A(_0894_),
    .Z(_1060_));
 MUX2_X1 _3350_ (.A(\mem[9][16] ),
    .B(\mem[13][16] ),
    .S(_1060_),
    .Z(_1061_));
 NOR2_X1 _3351_ (.A1(_0872_),
    .A2(_1061_),
    .ZN(_1062_));
 BUF_X4 _3352_ (.A(_0918_),
    .Z(_1063_));
 MUX2_X1 _3353_ (.A(\mem[0][16] ),
    .B(\mem[4][16] ),
    .S(_0994_),
    .Z(_1064_));
 NOR2_X1 _3354_ (.A1(_1063_),
    .A2(_1064_),
    .ZN(_1065_));
 BUF_X4 _3355_ (.A(_0886_),
    .Z(_1066_));
 MUX2_X1 _3356_ (.A(\mem[1][16] ),
    .B(\mem[5][16] ),
    .S(_0924_),
    .Z(_1067_));
 NOR2_X1 _3357_ (.A1(_1066_),
    .A2(_1067_),
    .ZN(_1068_));
 OAI33_X1 _3358_ (.A1(_0913_),
    .A2(_1059_),
    .A3(_1062_),
    .B1(_1065_),
    .B2(_1068_),
    .B3(_0900_),
    .ZN(_1069_));
 MUX2_X1 _3359_ (.A(\mem[10][16] ),
    .B(\mem[14][16] ),
    .S(_1021_),
    .Z(_1070_));
 NOR2_X1 _3360_ (.A1(_0929_),
    .A2(_1070_),
    .ZN(_1071_));
 MUX2_X1 _3361_ (.A(\mem[11][16] ),
    .B(\mem[15][16] ),
    .S(_0979_),
    .Z(_1072_));
 NOR2_X1 _3362_ (.A1(_0893_),
    .A2(_1072_),
    .ZN(_1073_));
 MUX2_X1 _3363_ (.A(\mem[2][16] ),
    .B(\mem[6][16] ),
    .S(_0959_),
    .Z(_1074_));
 NOR2_X1 _3364_ (.A1(_1049_),
    .A2(_1074_),
    .ZN(_1075_));
 BUF_X4 _3365_ (.A(_0882_),
    .Z(_1076_));
 MUX2_X1 _3366_ (.A(\mem[3][16] ),
    .B(\mem[7][16] ),
    .S(_1076_),
    .Z(_1077_));
 NOR2_X1 _3367_ (.A1(_1028_),
    .A2(_1077_),
    .ZN(_1078_));
 OAI33_X1 _3368_ (.A1(_0928_),
    .A2(_1071_),
    .A3(_1073_),
    .B1(_1075_),
    .B2(_1078_),
    .B3(_0880_),
    .ZN(_1079_));
 OAI221_X1 _3369_ (.A(_0861_),
    .B1(_1069_),
    .B2(_1079_),
    .C1(_0942_),
    .C2(_1032_),
    .ZN(_1080_));
 NAND2_X1 _3370_ (.A1(\last_valid_data[16] ),
    .A2(_0908_),
    .ZN(_1081_));
 BUF_X8 _3371_ (.A(net68),
    .Z(_1082_));
 NAND2_X1 _3372_ (.A1(_0911_),
    .A2(\last_valid_data[16] ),
    .ZN(_1083_));
 OAI221_X1 _3373_ (.A(_1080_),
    .B1(_1081_),
    .B2(_1082_),
    .C1(_1083_),
    .C2(_0856_),
    .ZN(_0038_));
 MUX2_X1 _3374_ (.A(\mem[8][17] ),
    .B(\mem[12][17] ),
    .S(_0867_),
    .Z(_1084_));
 NOR2_X1 _3375_ (.A1(_0864_),
    .A2(_1084_),
    .ZN(_1085_));
 MUX2_X1 _3376_ (.A(\mem[9][17] ),
    .B(\mem[13][17] ),
    .S(_1060_),
    .Z(_1086_));
 NOR2_X1 _3377_ (.A1(_0872_),
    .A2(_1086_),
    .ZN(_1087_));
 MUX2_X1 _3378_ (.A(\mem[0][17] ),
    .B(\mem[4][17] ),
    .S(_0994_),
    .Z(_1088_));
 NOR2_X1 _3379_ (.A1(_1063_),
    .A2(_1088_),
    .ZN(_1089_));
 MUX2_X1 _3380_ (.A(\mem[1][17] ),
    .B(\mem[5][17] ),
    .S(_0924_),
    .Z(_1090_));
 NOR2_X1 _3381_ (.A1(_1066_),
    .A2(_1090_),
    .ZN(_1091_));
 OAI33_X1 _3382_ (.A1(_0913_),
    .A2(_1085_),
    .A3(_1087_),
    .B1(_1089_),
    .B2(_1091_),
    .B3(_0900_),
    .ZN(_1092_));
 BUF_X4 _3383_ (.A(_0918_),
    .Z(_1093_));
 MUX2_X1 _3384_ (.A(\mem[10][17] ),
    .B(\mem[14][17] ),
    .S(_1021_),
    .Z(_1094_));
 NOR2_X1 _3385_ (.A1(_1093_),
    .A2(_1094_),
    .ZN(_1095_));
 BUF_X4 _3386_ (.A(_0886_),
    .Z(_1096_));
 MUX2_X1 _3387_ (.A(\mem[11][17] ),
    .B(\mem[15][17] ),
    .S(_0979_),
    .Z(_1097_));
 NOR2_X1 _3388_ (.A1(_1096_),
    .A2(_1097_),
    .ZN(_1098_));
 MUX2_X1 _3389_ (.A(\mem[2][17] ),
    .B(\mem[6][17] ),
    .S(_0959_),
    .Z(_1099_));
 NOR2_X1 _3390_ (.A1(_1049_),
    .A2(_1099_),
    .ZN(_1100_));
 MUX2_X1 _3391_ (.A(\mem[3][17] ),
    .B(\mem[7][17] ),
    .S(_1076_),
    .Z(_1101_));
 NOR2_X1 _3392_ (.A1(_1028_),
    .A2(_1101_),
    .ZN(_1102_));
 OAI33_X1 _3393_ (.A1(_0928_),
    .A2(_1095_),
    .A3(_1098_),
    .B1(_1100_),
    .B2(_1102_),
    .B3(_0880_),
    .ZN(_1103_));
 OAI221_X1 _3394_ (.A(_0861_),
    .B1(_1092_),
    .B2(_1103_),
    .C1(_0942_),
    .C2(_1032_),
    .ZN(_1104_));
 NAND2_X1 _3395_ (.A1(\last_valid_data[17] ),
    .A2(_0908_),
    .ZN(_1105_));
 NAND2_X1 _3396_ (.A1(_0911_),
    .A2(\last_valid_data[17] ),
    .ZN(_1106_));
 CLKBUF_X3 _3397_ (.A(_0763_),
    .Z(_1107_));
 OAI221_X1 _3398_ (.A(_1104_),
    .B1(_1105_),
    .B2(_1082_),
    .C1(_1106_),
    .C2(_1107_),
    .ZN(_0039_));
 BUF_X4 _3399_ (.A(_0863_),
    .Z(_1108_));
 BUF_X4 _3400_ (.A(_0866_),
    .Z(_1109_));
 MUX2_X1 _3401_ (.A(\mem[8][18] ),
    .B(\mem[12][18] ),
    .S(_1109_),
    .Z(_1110_));
 NOR2_X1 _3402_ (.A1(_1108_),
    .A2(_1110_),
    .ZN(_1111_));
 MUX2_X1 _3403_ (.A(\mem[9][18] ),
    .B(\mem[13][18] ),
    .S(_1060_),
    .Z(_1112_));
 NOR2_X1 _3404_ (.A1(_0872_),
    .A2(_1112_),
    .ZN(_1113_));
 MUX2_X1 _3405_ (.A(\mem[0][18] ),
    .B(\mem[4][18] ),
    .S(_0994_),
    .Z(_1114_));
 NOR2_X1 _3406_ (.A1(_1063_),
    .A2(_1114_),
    .ZN(_1115_));
 MUX2_X1 _3407_ (.A(\mem[1][18] ),
    .B(\mem[5][18] ),
    .S(_0924_),
    .Z(_1116_));
 NOR2_X1 _3408_ (.A1(_1066_),
    .A2(_1116_),
    .ZN(_1117_));
 OAI33_X1 _3409_ (.A1(_0913_),
    .A2(_1111_),
    .A3(_1113_),
    .B1(_1115_),
    .B2(_1117_),
    .B3(_0900_),
    .ZN(_1118_));
 MUX2_X1 _3410_ (.A(\mem[10][18] ),
    .B(\mem[14][18] ),
    .S(_1021_),
    .Z(_1119_));
 NOR2_X1 _3411_ (.A1(_1093_),
    .A2(_1119_),
    .ZN(_1120_));
 MUX2_X1 _3412_ (.A(\mem[11][18] ),
    .B(\mem[15][18] ),
    .S(_0979_),
    .Z(_1121_));
 NOR2_X1 _3413_ (.A1(_1096_),
    .A2(_1121_),
    .ZN(_1122_));
 MUX2_X1 _3414_ (.A(\mem[2][18] ),
    .B(\mem[6][18] ),
    .S(_0959_),
    .Z(_1123_));
 NOR2_X1 _3415_ (.A1(_1049_),
    .A2(_1123_),
    .ZN(_1124_));
 MUX2_X1 _3416_ (.A(\mem[3][18] ),
    .B(\mem[7][18] ),
    .S(_1076_),
    .Z(_1125_));
 NOR2_X1 _3417_ (.A1(_1028_),
    .A2(_1125_),
    .ZN(_1126_));
 OAI33_X1 _3418_ (.A1(_0928_),
    .A2(_1120_),
    .A3(_1122_),
    .B1(_1124_),
    .B2(_1126_),
    .B3(_0880_),
    .ZN(_1127_));
 CLKBUF_X3 _3419_ (.A(_0815_),
    .Z(_1128_));
 OAI221_X1 _3420_ (.A(_0861_),
    .B1(_1118_),
    .B2(_1127_),
    .C1(_1128_),
    .C2(_1032_),
    .ZN(_1129_));
 NAND2_X1 _3421_ (.A1(\last_valid_data[18] ),
    .A2(_0908_),
    .ZN(_1130_));
 NAND2_X1 _3422_ (.A1(_0911_),
    .A2(\last_valid_data[18] ),
    .ZN(_1131_));
 OAI221_X1 _3423_ (.A(_1129_),
    .B1(_1130_),
    .B2(_1082_),
    .C1(_1131_),
    .C2(_1107_),
    .ZN(_0040_));
 CLKBUF_X3 _3424_ (.A(_0860_),
    .Z(_1132_));
 MUX2_X1 _3425_ (.A(\mem[8][19] ),
    .B(\mem[12][19] ),
    .S(_1109_),
    .Z(_1133_));
 NOR2_X1 _3426_ (.A1(_1108_),
    .A2(_1133_),
    .ZN(_1134_));
 BUF_X4 _3427_ (.A(_0871_),
    .Z(_1135_));
 MUX2_X1 _3428_ (.A(\mem[9][19] ),
    .B(\mem[13][19] ),
    .S(_1060_),
    .Z(_1136_));
 NOR2_X1 _3429_ (.A1(_1135_),
    .A2(_1136_),
    .ZN(_1137_));
 MUX2_X1 _3430_ (.A(\mem[0][19] ),
    .B(\mem[4][19] ),
    .S(_0994_),
    .Z(_1138_));
 NOR2_X1 _3431_ (.A1(_1063_),
    .A2(_1138_),
    .ZN(_1139_));
 MUX2_X1 _3432_ (.A(\mem[1][19] ),
    .B(\mem[5][19] ),
    .S(_0924_),
    .Z(_1140_));
 NOR2_X1 _3433_ (.A1(_1066_),
    .A2(_1140_),
    .ZN(_1141_));
 BUF_X4 _3434_ (.A(_0899_),
    .Z(_1142_));
 OAI33_X1 _3435_ (.A1(_0913_),
    .A2(_1134_),
    .A3(_1137_),
    .B1(_1139_),
    .B2(_1141_),
    .B3(_1142_),
    .ZN(_1143_));
 MUX2_X1 _3436_ (.A(\mem[10][19] ),
    .B(\mem[14][19] ),
    .S(_1021_),
    .Z(_1144_));
 NOR2_X1 _3437_ (.A1(_1093_),
    .A2(_1144_),
    .ZN(_1145_));
 MUX2_X1 _3438_ (.A(\mem[11][19] ),
    .B(\mem[15][19] ),
    .S(_0979_),
    .Z(_1146_));
 NOR2_X1 _3439_ (.A1(_1096_),
    .A2(_1146_),
    .ZN(_1147_));
 MUX2_X1 _3440_ (.A(\mem[2][19] ),
    .B(\mem[6][19] ),
    .S(_0959_),
    .Z(_1148_));
 NOR2_X1 _3441_ (.A1(_1049_),
    .A2(_1148_),
    .ZN(_1149_));
 MUX2_X1 _3442_ (.A(\mem[3][19] ),
    .B(\mem[7][19] ),
    .S(_1076_),
    .Z(_1150_));
 NOR2_X1 _3443_ (.A1(_1028_),
    .A2(_1150_),
    .ZN(_1151_));
 CLKBUF_X3 _3444_ (.A(_0879_),
    .Z(_1152_));
 OAI33_X1 _3445_ (.A1(_0928_),
    .A2(_1145_),
    .A3(_1147_),
    .B1(_1149_),
    .B2(_1151_),
    .B3(_1152_),
    .ZN(_1153_));
 OAI221_X1 _3446_ (.A(_1132_),
    .B1(_1143_),
    .B2(_1153_),
    .C1(_1128_),
    .C2(_1032_),
    .ZN(_1154_));
 CLKBUF_X3 _3447_ (.A(_0761_),
    .Z(_1155_));
 NAND2_X1 _3448_ (.A1(\last_valid_data[19] ),
    .A2(_1155_),
    .ZN(_1156_));
 CLKBUF_X3 _3449_ (.A(_0859_),
    .Z(_1157_));
 NAND2_X1 _3450_ (.A1(_1157_),
    .A2(\last_valid_data[19] ),
    .ZN(_1158_));
 OAI221_X1 _3451_ (.A(_1154_),
    .B1(_1156_),
    .B2(_1082_),
    .C1(_1158_),
    .C2(_1107_),
    .ZN(_0041_));
 BUF_X4 _3452_ (.A(_0901_),
    .Z(_1159_));
 MUX2_X1 _3453_ (.A(\mem[8][1] ),
    .B(\mem[12][1] ),
    .S(_1109_),
    .Z(_1160_));
 NOR2_X1 _3454_ (.A1(_1108_),
    .A2(_1160_),
    .ZN(_1161_));
 MUX2_X1 _3455_ (.A(\mem[9][1] ),
    .B(\mem[13][1] ),
    .S(_1060_),
    .Z(_1162_));
 NOR2_X1 _3456_ (.A1(_1135_),
    .A2(_1162_),
    .ZN(_1163_));
 MUX2_X1 _3457_ (.A(\mem[0][1] ),
    .B(\mem[4][1] ),
    .S(_0994_),
    .Z(_1164_));
 NOR2_X1 _3458_ (.A1(_1063_),
    .A2(_1164_),
    .ZN(_1165_));
 BUF_X4 _3459_ (.A(_0882_),
    .Z(_1166_));
 MUX2_X1 _3460_ (.A(\mem[1][1] ),
    .B(\mem[5][1] ),
    .S(_1166_),
    .Z(_1167_));
 NOR2_X1 _3461_ (.A1(_1066_),
    .A2(_1167_),
    .ZN(_1168_));
 OAI33_X1 _3462_ (.A1(_1159_),
    .A2(_1161_),
    .A3(_1163_),
    .B1(_1165_),
    .B2(_1168_),
    .B3(_1142_),
    .ZN(_1169_));
 BUF_X4 _3463_ (.A(_0881_),
    .Z(_1170_));
 MUX2_X1 _3464_ (.A(\mem[10][1] ),
    .B(\mem[14][1] ),
    .S(_1021_),
    .Z(_1171_));
 NOR2_X1 _3465_ (.A1(_1093_),
    .A2(_1171_),
    .ZN(_1172_));
 MUX2_X1 _3466_ (.A(\mem[11][1] ),
    .B(\mem[15][1] ),
    .S(_0979_),
    .Z(_1173_));
 NOR2_X1 _3467_ (.A1(_1096_),
    .A2(_1173_),
    .ZN(_1174_));
 MUX2_X1 _3468_ (.A(\mem[2][1] ),
    .B(\mem[6][1] ),
    .S(_0959_),
    .Z(_1175_));
 NOR2_X1 _3469_ (.A1(_1049_),
    .A2(_1175_),
    .ZN(_1176_));
 MUX2_X1 _3470_ (.A(\mem[3][1] ),
    .B(\mem[7][1] ),
    .S(_1076_),
    .Z(_1177_));
 NOR2_X1 _3471_ (.A1(_1028_),
    .A2(_1177_),
    .ZN(_1178_));
 OAI33_X1 _3472_ (.A1(_1170_),
    .A2(_1172_),
    .A3(_1174_),
    .B1(_1176_),
    .B2(_1178_),
    .B3(_1152_),
    .ZN(_1179_));
 OAI221_X1 _3473_ (.A(_1132_),
    .B1(_1169_),
    .B2(_1179_),
    .C1(_1128_),
    .C2(_1032_),
    .ZN(_1180_));
 NAND2_X1 _3474_ (.A1(\last_valid_data[1] ),
    .A2(_1155_),
    .ZN(_1181_));
 NAND2_X1 _3475_ (.A1(_1157_),
    .A2(\last_valid_data[1] ),
    .ZN(_1182_));
 OAI221_X1 _3476_ (.A(_1180_),
    .B1(_1181_),
    .B2(_1082_),
    .C1(_1182_),
    .C2(_1107_),
    .ZN(_0042_));
 MUX2_X1 _3477_ (.A(\mem[8][20] ),
    .B(\mem[12][20] ),
    .S(_1109_),
    .Z(_1183_));
 NOR2_X1 _3478_ (.A1(_1108_),
    .A2(_1183_),
    .ZN(_1184_));
 MUX2_X1 _3479_ (.A(\mem[9][20] ),
    .B(\mem[13][20] ),
    .S(_1060_),
    .Z(_1185_));
 NOR2_X1 _3480_ (.A1(_1135_),
    .A2(_1185_),
    .ZN(_1186_));
 MUX2_X1 _3481_ (.A(\mem[0][20] ),
    .B(\mem[4][20] ),
    .S(_0994_),
    .Z(_1187_));
 NOR2_X1 _3482_ (.A1(_1063_),
    .A2(_1187_),
    .ZN(_1188_));
 MUX2_X1 _3483_ (.A(\mem[1][20] ),
    .B(\mem[5][20] ),
    .S(_1166_),
    .Z(_1189_));
 NOR2_X1 _3484_ (.A1(_1066_),
    .A2(_1189_),
    .ZN(_1190_));
 OAI33_X1 _3485_ (.A1(_1159_),
    .A2(_1184_),
    .A3(_1186_),
    .B1(_1188_),
    .B2(_1190_),
    .B3(_1142_),
    .ZN(_1191_));
 MUX2_X1 _3486_ (.A(\mem[10][20] ),
    .B(\mem[14][20] ),
    .S(_1021_),
    .Z(_1192_));
 NOR2_X1 _3487_ (.A1(_1093_),
    .A2(_1192_),
    .ZN(_1193_));
 MUX2_X1 _3488_ (.A(\mem[11][20] ),
    .B(\mem[15][20] ),
    .S(_0979_),
    .Z(_1194_));
 NOR2_X1 _3489_ (.A1(_1096_),
    .A2(_1194_),
    .ZN(_1195_));
 BUF_X4 _3490_ (.A(_0882_),
    .Z(_1196_));
 MUX2_X1 _3491_ (.A(\mem[2][20] ),
    .B(\mem[6][20] ),
    .S(_1196_),
    .Z(_1197_));
 NOR2_X1 _3492_ (.A1(_1049_),
    .A2(_1197_),
    .ZN(_1198_));
 MUX2_X1 _3493_ (.A(\mem[3][20] ),
    .B(\mem[7][20] ),
    .S(_1076_),
    .Z(_1199_));
 NOR2_X1 _3494_ (.A1(_1028_),
    .A2(_1199_),
    .ZN(_1200_));
 OAI33_X1 _3495_ (.A1(_1170_),
    .A2(_1193_),
    .A3(_1195_),
    .B1(_1198_),
    .B2(_1200_),
    .B3(_1152_),
    .ZN(_1201_));
 OAI221_X1 _3496_ (.A(_1132_),
    .B1(_1191_),
    .B2(_1201_),
    .C1(_1128_),
    .C2(_1032_),
    .ZN(_1202_));
 NAND2_X1 _3497_ (.A1(\last_valid_data[20] ),
    .A2(_1155_),
    .ZN(_1203_));
 NAND2_X1 _3498_ (.A1(_1157_),
    .A2(\last_valid_data[20] ),
    .ZN(_1204_));
 OAI221_X1 _3499_ (.A(_1202_),
    .B1(_1203_),
    .B2(_1082_),
    .C1(_1204_),
    .C2(_1107_),
    .ZN(_0043_));
 MUX2_X1 _3500_ (.A(\mem[8][21] ),
    .B(\mem[12][21] ),
    .S(_1109_),
    .Z(_1205_));
 NOR2_X1 _3501_ (.A1(_1108_),
    .A2(_1205_),
    .ZN(_1206_));
 MUX2_X1 _3502_ (.A(\mem[9][21] ),
    .B(\mem[13][21] ),
    .S(_1060_),
    .Z(_1207_));
 NOR2_X1 _3503_ (.A1(_1135_),
    .A2(_1207_),
    .ZN(_1208_));
 MUX2_X1 _3504_ (.A(\mem[0][21] ),
    .B(\mem[4][21] ),
    .S(_0994_),
    .Z(_1209_));
 NOR2_X1 _3505_ (.A1(_1063_),
    .A2(_1209_),
    .ZN(_1210_));
 MUX2_X1 _3506_ (.A(\mem[1][21] ),
    .B(\mem[5][21] ),
    .S(_1166_),
    .Z(_1211_));
 NOR2_X1 _3507_ (.A1(_1066_),
    .A2(_1211_),
    .ZN(_1212_));
 OAI33_X1 _3508_ (.A1(_1159_),
    .A2(_1206_),
    .A3(_1208_),
    .B1(_1210_),
    .B2(_1212_),
    .B3(_1142_),
    .ZN(_1213_));
 MUX2_X1 _3509_ (.A(\mem[10][21] ),
    .B(\mem[14][21] ),
    .S(_1021_),
    .Z(_1214_));
 NOR2_X1 _3510_ (.A1(_1093_),
    .A2(_1214_),
    .ZN(_1215_));
 BUF_X4 _3511_ (.A(_0882_),
    .Z(_1216_));
 MUX2_X1 _3512_ (.A(\mem[11][21] ),
    .B(\mem[15][21] ),
    .S(_1216_),
    .Z(_1217_));
 NOR2_X1 _3513_ (.A1(_1096_),
    .A2(_1217_),
    .ZN(_1218_));
 MUX2_X1 _3514_ (.A(\mem[2][21] ),
    .B(\mem[6][21] ),
    .S(_1196_),
    .Z(_1219_));
 NOR2_X1 _3515_ (.A1(_1049_),
    .A2(_1219_),
    .ZN(_1220_));
 MUX2_X1 _3516_ (.A(\mem[3][21] ),
    .B(\mem[7][21] ),
    .S(_1076_),
    .Z(_1221_));
 NOR2_X1 _3517_ (.A1(_1028_),
    .A2(_1221_),
    .ZN(_1222_));
 OAI33_X1 _3518_ (.A1(_1170_),
    .A2(_1215_),
    .A3(_1218_),
    .B1(_1220_),
    .B2(_1222_),
    .B3(_1152_),
    .ZN(_1223_));
 OAI221_X1 _3519_ (.A(_1132_),
    .B1(_1213_),
    .B2(_1223_),
    .C1(_1128_),
    .C2(_1032_),
    .ZN(_1224_));
 NAND2_X1 _3520_ (.A1(\last_valid_data[21] ),
    .A2(_1155_),
    .ZN(_1225_));
 NAND2_X1 _3521_ (.A1(_1157_),
    .A2(\last_valid_data[21] ),
    .ZN(_1226_));
 OAI221_X1 _3522_ (.A(_1224_),
    .B1(_1225_),
    .B2(_1082_),
    .C1(_1226_),
    .C2(_1107_),
    .ZN(_0044_));
 MUX2_X1 _3523_ (.A(\mem[8][22] ),
    .B(\mem[12][22] ),
    .S(_1109_),
    .Z(_1227_));
 NOR2_X1 _3524_ (.A1(_1108_),
    .A2(_1227_),
    .ZN(_1228_));
 MUX2_X1 _3525_ (.A(\mem[9][22] ),
    .B(\mem[13][22] ),
    .S(_1060_),
    .Z(_1229_));
 NOR2_X1 _3526_ (.A1(_1135_),
    .A2(_1229_),
    .ZN(_1230_));
 BUF_X4 _3527_ (.A(_0894_),
    .Z(_1231_));
 MUX2_X1 _3528_ (.A(\mem[0][22] ),
    .B(\mem[4][22] ),
    .S(_1231_),
    .Z(_1232_));
 NOR2_X1 _3529_ (.A1(_1063_),
    .A2(_1232_),
    .ZN(_1233_));
 MUX2_X1 _3530_ (.A(\mem[1][22] ),
    .B(\mem[5][22] ),
    .S(_1166_),
    .Z(_1234_));
 NOR2_X1 _3531_ (.A1(_1066_),
    .A2(_1234_),
    .ZN(_1235_));
 OAI33_X1 _3532_ (.A1(_1159_),
    .A2(_1228_),
    .A3(_1230_),
    .B1(_1233_),
    .B2(_1235_),
    .B3(_1142_),
    .ZN(_1236_));
 MUX2_X1 _3533_ (.A(\mem[10][22] ),
    .B(\mem[14][22] ),
    .S(_1021_),
    .Z(_1237_));
 NOR2_X1 _3534_ (.A1(_1093_),
    .A2(_1237_),
    .ZN(_1238_));
 MUX2_X1 _3535_ (.A(\mem[11][22] ),
    .B(\mem[15][22] ),
    .S(_1216_),
    .Z(_1239_));
 NOR2_X1 _3536_ (.A1(_1096_),
    .A2(_1239_),
    .ZN(_1240_));
 MUX2_X1 _3537_ (.A(\mem[2][22] ),
    .B(\mem[6][22] ),
    .S(_1196_),
    .Z(_1241_));
 NOR2_X1 _3538_ (.A1(_1049_),
    .A2(_1241_),
    .ZN(_1242_));
 MUX2_X1 _3539_ (.A(\mem[3][22] ),
    .B(\mem[7][22] ),
    .S(_1076_),
    .Z(_1243_));
 NOR2_X1 _3540_ (.A1(_1028_),
    .A2(_1243_),
    .ZN(_1244_));
 OAI33_X1 _3541_ (.A1(_1170_),
    .A2(_1238_),
    .A3(_1240_),
    .B1(_1242_),
    .B2(_1244_),
    .B3(_1152_),
    .ZN(_1245_));
 OAI221_X1 _3542_ (.A(_1132_),
    .B1(_1236_),
    .B2(_1245_),
    .C1(_1128_),
    .C2(_1032_),
    .ZN(_1246_));
 NAND2_X1 _3543_ (.A1(\last_valid_data[22] ),
    .A2(_1155_),
    .ZN(_1247_));
 NAND2_X1 _3544_ (.A1(_1157_),
    .A2(\last_valid_data[22] ),
    .ZN(_1248_));
 OAI221_X1 _3545_ (.A(_1246_),
    .B1(_1247_),
    .B2(_1082_),
    .C1(_1248_),
    .C2(_1107_),
    .ZN(_0045_));
 MUX2_X1 _3546_ (.A(\mem[8][23] ),
    .B(\mem[12][23] ),
    .S(_1109_),
    .Z(_1249_));
 NOR2_X1 _3547_ (.A1(_1108_),
    .A2(_1249_),
    .ZN(_1250_));
 MUX2_X1 _3548_ (.A(\mem[9][23] ),
    .B(\mem[13][23] ),
    .S(_1060_),
    .Z(_1251_));
 NOR2_X1 _3549_ (.A1(_1135_),
    .A2(_1251_),
    .ZN(_1252_));
 MUX2_X1 _3550_ (.A(\mem[0][23] ),
    .B(\mem[4][23] ),
    .S(_1231_),
    .Z(_1253_));
 NOR2_X1 _3551_ (.A1(_1063_),
    .A2(_1253_),
    .ZN(_1254_));
 MUX2_X1 _3552_ (.A(\mem[1][23] ),
    .B(\mem[5][23] ),
    .S(_1166_),
    .Z(_1255_));
 NOR2_X1 _3553_ (.A1(_1066_),
    .A2(_1255_),
    .ZN(_1256_));
 OAI33_X1 _3554_ (.A1(_1159_),
    .A2(_1250_),
    .A3(_1252_),
    .B1(_1254_),
    .B2(_1256_),
    .B3(_1142_),
    .ZN(_1257_));
 BUF_X4 _3555_ (.A(_0894_),
    .Z(_1258_));
 MUX2_X1 _3556_ (.A(\mem[10][23] ),
    .B(\mem[14][23] ),
    .S(_1258_),
    .Z(_1259_));
 NOR2_X1 _3557_ (.A1(_1093_),
    .A2(_1259_),
    .ZN(_1260_));
 MUX2_X1 _3558_ (.A(\mem[11][23] ),
    .B(\mem[15][23] ),
    .S(_1216_),
    .Z(_1261_));
 NOR2_X1 _3559_ (.A1(_1096_),
    .A2(_1261_),
    .ZN(_1262_));
 MUX2_X1 _3560_ (.A(\mem[2][23] ),
    .B(\mem[6][23] ),
    .S(_1196_),
    .Z(_1263_));
 NOR2_X1 _3561_ (.A1(_1049_),
    .A2(_1263_),
    .ZN(_1264_));
 CLKBUF_X3 _3562_ (.A(_0886_),
    .Z(_1265_));
 MUX2_X1 _3563_ (.A(\mem[3][23] ),
    .B(\mem[7][23] ),
    .S(_1076_),
    .Z(_1266_));
 NOR2_X1 _3564_ (.A1(_1265_),
    .A2(_1266_),
    .ZN(_1267_));
 OAI33_X1 _3565_ (.A1(_1170_),
    .A2(_1260_),
    .A3(_1262_),
    .B1(_1264_),
    .B2(_1267_),
    .B3(_1152_),
    .ZN(_1268_));
 CLKBUF_X3 _3566_ (.A(_0595_),
    .Z(_1269_));
 OAI221_X1 _3567_ (.A(_1132_),
    .B1(_1257_),
    .B2(_1268_),
    .C1(_1128_),
    .C2(_1269_),
    .ZN(_1270_));
 NAND2_X1 _3568_ (.A1(\last_valid_data[23] ),
    .A2(_1155_),
    .ZN(_1271_));
 NAND2_X1 _3569_ (.A1(_1157_),
    .A2(\last_valid_data[23] ),
    .ZN(_1272_));
 OAI221_X1 _3570_ (.A(_1270_),
    .B1(_1271_),
    .B2(_1082_),
    .C1(_1272_),
    .C2(_1107_),
    .ZN(_0046_));
 MUX2_X1 _3571_ (.A(\mem[8][24] ),
    .B(\mem[12][24] ),
    .S(_1109_),
    .Z(_1273_));
 NOR2_X1 _3572_ (.A1(_1108_),
    .A2(_1273_),
    .ZN(_1274_));
 MUX2_X1 _3573_ (.A(\mem[9][24] ),
    .B(\mem[13][24] ),
    .S(_1060_),
    .Z(_1275_));
 NOR2_X1 _3574_ (.A1(_1135_),
    .A2(_1275_),
    .ZN(_1276_));
 MUX2_X1 _3575_ (.A(\mem[0][24] ),
    .B(\mem[4][24] ),
    .S(_1231_),
    .Z(_1277_));
 NOR2_X1 _3576_ (.A1(_1063_),
    .A2(_1277_),
    .ZN(_1278_));
 MUX2_X1 _3577_ (.A(\mem[1][24] ),
    .B(\mem[5][24] ),
    .S(_1166_),
    .Z(_1279_));
 NOR2_X1 _3578_ (.A1(_1066_),
    .A2(_1279_),
    .ZN(_1280_));
 OAI33_X1 _3579_ (.A1(_1159_),
    .A2(_1274_),
    .A3(_1276_),
    .B1(_1278_),
    .B2(_1280_),
    .B3(_1142_),
    .ZN(_1281_));
 MUX2_X1 _3580_ (.A(\mem[10][24] ),
    .B(\mem[14][24] ),
    .S(_1258_),
    .Z(_1282_));
 NOR2_X1 _3581_ (.A1(_1093_),
    .A2(_1282_),
    .ZN(_1283_));
 MUX2_X1 _3582_ (.A(\mem[11][24] ),
    .B(\mem[15][24] ),
    .S(_1216_),
    .Z(_1284_));
 NOR2_X1 _3583_ (.A1(_1096_),
    .A2(_1284_),
    .ZN(_1285_));
 CLKBUF_X3 _3584_ (.A(_0918_),
    .Z(_1286_));
 MUX2_X1 _3585_ (.A(\mem[2][24] ),
    .B(\mem[6][24] ),
    .S(_1196_),
    .Z(_1287_));
 NOR2_X1 _3586_ (.A1(_1286_),
    .A2(_1287_),
    .ZN(_1288_));
 MUX2_X1 _3587_ (.A(\mem[3][24] ),
    .B(\mem[7][24] ),
    .S(_1076_),
    .Z(_1289_));
 NOR2_X1 _3588_ (.A1(_1265_),
    .A2(_1289_),
    .ZN(_1290_));
 OAI33_X1 _3589_ (.A1(_1170_),
    .A2(_1283_),
    .A3(_1285_),
    .B1(_1288_),
    .B2(_1290_),
    .B3(_1152_),
    .ZN(_1291_));
 OAI221_X1 _3590_ (.A(_1132_),
    .B1(_1281_),
    .B2(_1291_),
    .C1(_1128_),
    .C2(_1269_),
    .ZN(_1292_));
 NAND2_X1 _3591_ (.A1(\last_valid_data[24] ),
    .A2(_1155_),
    .ZN(_1293_));
 NAND2_X1 _3592_ (.A1(_1157_),
    .A2(\last_valid_data[24] ),
    .ZN(_1294_));
 OAI221_X1 _3593_ (.A(_1292_),
    .B1(_1293_),
    .B2(_1082_),
    .C1(_1294_),
    .C2(_1107_),
    .ZN(_0047_));
 MUX2_X1 _3594_ (.A(\mem[8][25] ),
    .B(\mem[12][25] ),
    .S(_1109_),
    .Z(_1295_));
 NOR2_X1 _3595_ (.A1(_1108_),
    .A2(_1295_),
    .ZN(_1296_));
 BUF_X4 _3596_ (.A(_0894_),
    .Z(_1297_));
 MUX2_X1 _3597_ (.A(\mem[9][25] ),
    .B(\mem[13][25] ),
    .S(_1297_),
    .Z(_1298_));
 NOR2_X1 _3598_ (.A1(_1135_),
    .A2(_1298_),
    .ZN(_1299_));
 BUF_X4 _3599_ (.A(_0918_),
    .Z(_1300_));
 MUX2_X1 _3600_ (.A(\mem[0][25] ),
    .B(\mem[4][25] ),
    .S(_1231_),
    .Z(_1301_));
 NOR2_X1 _3601_ (.A1(_1300_),
    .A2(_1301_),
    .ZN(_1302_));
 BUF_X4 _3602_ (.A(_0886_),
    .Z(_1303_));
 MUX2_X1 _3603_ (.A(\mem[1][25] ),
    .B(\mem[5][25] ),
    .S(_1166_),
    .Z(_1304_));
 NOR2_X1 _3604_ (.A1(_1303_),
    .A2(_1304_),
    .ZN(_1305_));
 OAI33_X1 _3605_ (.A1(_1159_),
    .A2(_1296_),
    .A3(_1299_),
    .B1(_1302_),
    .B2(_1305_),
    .B3(_1142_),
    .ZN(_1306_));
 MUX2_X1 _3606_ (.A(\mem[10][25] ),
    .B(\mem[14][25] ),
    .S(_1258_),
    .Z(_1307_));
 NOR2_X1 _3607_ (.A1(_1093_),
    .A2(_1307_),
    .ZN(_1308_));
 MUX2_X1 _3608_ (.A(\mem[11][25] ),
    .B(\mem[15][25] ),
    .S(_1216_),
    .Z(_1309_));
 NOR2_X1 _3609_ (.A1(_1096_),
    .A2(_1309_),
    .ZN(_1310_));
 MUX2_X1 _3610_ (.A(\mem[2][25] ),
    .B(\mem[6][25] ),
    .S(_1196_),
    .Z(_1311_));
 NOR2_X1 _3611_ (.A1(_1286_),
    .A2(_1311_),
    .ZN(_1312_));
 BUF_X4 _3612_ (.A(_0865_),
    .Z(_1313_));
 MUX2_X1 _3613_ (.A(\mem[3][25] ),
    .B(\mem[7][25] ),
    .S(_1313_),
    .Z(_1314_));
 NOR2_X1 _3614_ (.A1(_1265_),
    .A2(_1314_),
    .ZN(_1315_));
 OAI33_X1 _3615_ (.A1(_1170_),
    .A2(_1308_),
    .A3(_1310_),
    .B1(_1312_),
    .B2(_1315_),
    .B3(_1152_),
    .ZN(_1316_));
 OAI221_X1 _3616_ (.A(_1132_),
    .B1(_1306_),
    .B2(_1316_),
    .C1(_1128_),
    .C2(_1269_),
    .ZN(_1317_));
 NAND2_X1 _3617_ (.A1(\last_valid_data[25] ),
    .A2(_1155_),
    .ZN(_1318_));
 CLKBUF_X3 _3618_ (.A(_0606_),
    .Z(_1319_));
 NAND2_X1 _3619_ (.A1(_1157_),
    .A2(\last_valid_data[25] ),
    .ZN(_1320_));
 OAI221_X1 _3620_ (.A(_1317_),
    .B1(_1318_),
    .B2(_1319_),
    .C1(_1320_),
    .C2(_1107_),
    .ZN(_0048_));
 MUX2_X1 _3621_ (.A(\mem[8][26] ),
    .B(\mem[12][26] ),
    .S(_1109_),
    .Z(_1321_));
 NOR2_X1 _3622_ (.A1(_1108_),
    .A2(_1321_),
    .ZN(_1322_));
 MUX2_X1 _3623_ (.A(\mem[9][26] ),
    .B(\mem[13][26] ),
    .S(_1297_),
    .Z(_1323_));
 NOR2_X1 _3624_ (.A1(_1135_),
    .A2(_1323_),
    .ZN(_1324_));
 MUX2_X1 _3625_ (.A(\mem[0][26] ),
    .B(\mem[4][26] ),
    .S(_1231_),
    .Z(_1325_));
 NOR2_X1 _3626_ (.A1(_1300_),
    .A2(_1325_),
    .ZN(_1326_));
 MUX2_X1 _3627_ (.A(\mem[1][26] ),
    .B(\mem[5][26] ),
    .S(_1166_),
    .Z(_1327_));
 NOR2_X1 _3628_ (.A1(_1303_),
    .A2(_1327_),
    .ZN(_1328_));
 OAI33_X1 _3629_ (.A1(_1159_),
    .A2(_1322_),
    .A3(_1324_),
    .B1(_1326_),
    .B2(_1328_),
    .B3(_1142_),
    .ZN(_1329_));
 CLKBUF_X3 _3630_ (.A(_0918_),
    .Z(_1330_));
 MUX2_X1 _3631_ (.A(\mem[10][26] ),
    .B(\mem[14][26] ),
    .S(_1258_),
    .Z(_1331_));
 NOR2_X1 _3632_ (.A1(_1330_),
    .A2(_1331_),
    .ZN(_1332_));
 CLKBUF_X3 _3633_ (.A(_0886_),
    .Z(_1333_));
 MUX2_X1 _3634_ (.A(\mem[11][26] ),
    .B(\mem[15][26] ),
    .S(_1216_),
    .Z(_1334_));
 NOR2_X1 _3635_ (.A1(_1333_),
    .A2(_1334_),
    .ZN(_1335_));
 MUX2_X1 _3636_ (.A(\mem[2][26] ),
    .B(\mem[6][26] ),
    .S(_1196_),
    .Z(_1336_));
 NOR2_X1 _3637_ (.A1(_1286_),
    .A2(_1336_),
    .ZN(_1337_));
 MUX2_X1 _3638_ (.A(\mem[3][26] ),
    .B(\mem[7][26] ),
    .S(_1313_),
    .Z(_1338_));
 NOR2_X1 _3639_ (.A1(_1265_),
    .A2(_1338_),
    .ZN(_1339_));
 OAI33_X1 _3640_ (.A1(_1170_),
    .A2(_1332_),
    .A3(_1335_),
    .B1(_1337_),
    .B2(_1339_),
    .B3(_1152_),
    .ZN(_1340_));
 OAI221_X1 _3641_ (.A(_1132_),
    .B1(_1329_),
    .B2(_1340_),
    .C1(_1128_),
    .C2(_1269_),
    .ZN(_1341_));
 NAND2_X1 _3642_ (.A1(\last_valid_data[26] ),
    .A2(_1155_),
    .ZN(_1342_));
 NAND2_X1 _3643_ (.A1(_1157_),
    .A2(\last_valid_data[26] ),
    .ZN(_1343_));
 CLKBUF_X3 _3644_ (.A(_0763_),
    .Z(_1344_));
 OAI221_X1 _3645_ (.A(_1341_),
    .B1(_1342_),
    .B2(_1319_),
    .C1(_1343_),
    .C2(_1344_),
    .ZN(_0049_));
 BUF_X4 _3646_ (.A(_0918_),
    .Z(_1345_));
 BUF_X4 _3647_ (.A(_0866_),
    .Z(_1346_));
 MUX2_X1 _3648_ (.A(\mem[8][27] ),
    .B(\mem[12][27] ),
    .S(_1346_),
    .Z(_1347_));
 NOR2_X1 _3649_ (.A1(_1345_),
    .A2(_1347_),
    .ZN(_1348_));
 MUX2_X1 _3650_ (.A(\mem[9][27] ),
    .B(\mem[13][27] ),
    .S(_1297_),
    .Z(_1349_));
 NOR2_X1 _3651_ (.A1(_1135_),
    .A2(_1349_),
    .ZN(_1350_));
 MUX2_X1 _3652_ (.A(\mem[0][27] ),
    .B(\mem[4][27] ),
    .S(_1231_),
    .Z(_1351_));
 NOR2_X1 _3653_ (.A1(_1300_),
    .A2(_1351_),
    .ZN(_1352_));
 MUX2_X1 _3654_ (.A(\mem[1][27] ),
    .B(\mem[5][27] ),
    .S(_1166_),
    .Z(_1353_));
 NOR2_X1 _3655_ (.A1(_1303_),
    .A2(_1353_),
    .ZN(_1354_));
 OAI33_X1 _3656_ (.A1(_1159_),
    .A2(_1348_),
    .A3(_1350_),
    .B1(_1352_),
    .B2(_1354_),
    .B3(_1142_),
    .ZN(_1355_));
 MUX2_X1 _3657_ (.A(\mem[10][27] ),
    .B(\mem[14][27] ),
    .S(_1258_),
    .Z(_1356_));
 NOR2_X1 _3658_ (.A1(_1330_),
    .A2(_1356_),
    .ZN(_1357_));
 MUX2_X1 _3659_ (.A(\mem[11][27] ),
    .B(\mem[15][27] ),
    .S(_1216_),
    .Z(_1358_));
 NOR2_X1 _3660_ (.A1(_1333_),
    .A2(_1358_),
    .ZN(_1359_));
 MUX2_X1 _3661_ (.A(\mem[2][27] ),
    .B(\mem[6][27] ),
    .S(_1196_),
    .Z(_1360_));
 NOR2_X1 _3662_ (.A1(_1286_),
    .A2(_1360_),
    .ZN(_1361_));
 MUX2_X1 _3663_ (.A(\mem[3][27] ),
    .B(\mem[7][27] ),
    .S(_1313_),
    .Z(_1362_));
 NOR2_X1 _3664_ (.A1(_1265_),
    .A2(_1362_),
    .ZN(_1363_));
 OAI33_X1 _3665_ (.A1(_1170_),
    .A2(_1357_),
    .A3(_1359_),
    .B1(_1361_),
    .B2(_1363_),
    .B3(_1152_),
    .ZN(_1364_));
 CLKBUF_X3 _3666_ (.A(_0815_),
    .Z(_1365_));
 OAI221_X1 _3667_ (.A(_1132_),
    .B1(_1355_),
    .B2(_1364_),
    .C1(_1365_),
    .C2(_1269_),
    .ZN(_1366_));
 NAND2_X1 _3668_ (.A1(\last_valid_data[27] ),
    .A2(_1155_),
    .ZN(_1367_));
 NAND2_X1 _3669_ (.A1(_1157_),
    .A2(\last_valid_data[27] ),
    .ZN(_1368_));
 OAI221_X1 _3670_ (.A(_1366_),
    .B1(_1367_),
    .B2(_1319_),
    .C1(_1368_),
    .C2(_1344_),
    .ZN(_0050_));
 CLKBUF_X3 _3671_ (.A(_0860_),
    .Z(_1369_));
 MUX2_X1 _3672_ (.A(\mem[8][28] ),
    .B(\mem[12][28] ),
    .S(_1346_),
    .Z(_1370_));
 NOR2_X1 _3673_ (.A1(_1345_),
    .A2(_1370_),
    .ZN(_1371_));
 CLKBUF_X3 _3674_ (.A(_0886_),
    .Z(_1372_));
 MUX2_X1 _3675_ (.A(\mem[9][28] ),
    .B(\mem[13][28] ),
    .S(_1297_),
    .Z(_1373_));
 NOR2_X1 _3676_ (.A1(_1372_),
    .A2(_1373_),
    .ZN(_1374_));
 MUX2_X1 _3677_ (.A(\mem[0][28] ),
    .B(\mem[4][28] ),
    .S(_1231_),
    .Z(_1375_));
 NOR2_X1 _3678_ (.A1(_1300_),
    .A2(_1375_),
    .ZN(_1376_));
 MUX2_X1 _3679_ (.A(\mem[1][28] ),
    .B(\mem[5][28] ),
    .S(_1166_),
    .Z(_1377_));
 NOR2_X1 _3680_ (.A1(_1303_),
    .A2(_1377_),
    .ZN(_1378_));
 CLKBUF_X3 _3681_ (.A(_0899_),
    .Z(_1379_));
 OAI33_X1 _3682_ (.A1(_1159_),
    .A2(_1371_),
    .A3(_1374_),
    .B1(_1376_),
    .B2(_1378_),
    .B3(_1379_),
    .ZN(_1380_));
 MUX2_X1 _3683_ (.A(\mem[10][28] ),
    .B(\mem[14][28] ),
    .S(_1258_),
    .Z(_1381_));
 NOR2_X1 _3684_ (.A1(_1330_),
    .A2(_1381_),
    .ZN(_1382_));
 MUX2_X1 _3685_ (.A(\mem[11][28] ),
    .B(\mem[15][28] ),
    .S(_1216_),
    .Z(_1383_));
 NOR2_X1 _3686_ (.A1(_1333_),
    .A2(_1383_),
    .ZN(_1384_));
 MUX2_X1 _3687_ (.A(\mem[2][28] ),
    .B(\mem[6][28] ),
    .S(_1196_),
    .Z(_1385_));
 NOR2_X1 _3688_ (.A1(_1286_),
    .A2(_1385_),
    .ZN(_1386_));
 MUX2_X1 _3689_ (.A(\mem[3][28] ),
    .B(\mem[7][28] ),
    .S(_1313_),
    .Z(_1387_));
 NOR2_X1 _3690_ (.A1(_1265_),
    .A2(_1387_),
    .ZN(_1388_));
 CLKBUF_X3 _3691_ (.A(_0879_),
    .Z(_1389_));
 OAI33_X1 _3692_ (.A1(_1170_),
    .A2(_1382_),
    .A3(_1384_),
    .B1(_1386_),
    .B2(_1388_),
    .B3(_1389_),
    .ZN(_1390_));
 OAI221_X1 _3693_ (.A(_1369_),
    .B1(_1380_),
    .B2(_1390_),
    .C1(_1365_),
    .C2(_1269_),
    .ZN(_1391_));
 CLKBUF_X3 _3694_ (.A(_0761_),
    .Z(_1392_));
 NAND2_X1 _3695_ (.A1(\last_valid_data[28] ),
    .A2(_1392_),
    .ZN(_1393_));
 CLKBUF_X3 _3696_ (.A(_0859_),
    .Z(_1394_));
 NAND2_X1 _3697_ (.A1(_1394_),
    .A2(\last_valid_data[28] ),
    .ZN(_1395_));
 OAI221_X1 _3698_ (.A(_1391_),
    .B1(_1393_),
    .B2(_1319_),
    .C1(_1395_),
    .C2(_1344_),
    .ZN(_0051_));
 CLKBUF_X3 _3699_ (.A(_0901_),
    .Z(_1396_));
 MUX2_X1 _3700_ (.A(\mem[8][29] ),
    .B(\mem[12][29] ),
    .S(_1346_),
    .Z(_1397_));
 NOR2_X1 _3701_ (.A1(_1345_),
    .A2(_1397_),
    .ZN(_1398_));
 MUX2_X1 _3702_ (.A(\mem[9][29] ),
    .B(\mem[13][29] ),
    .S(_1297_),
    .Z(_1399_));
 NOR2_X1 _3703_ (.A1(_1372_),
    .A2(_1399_),
    .ZN(_1400_));
 MUX2_X1 _3704_ (.A(\mem[0][29] ),
    .B(\mem[4][29] ),
    .S(_1231_),
    .Z(_1401_));
 NOR2_X1 _3705_ (.A1(_1300_),
    .A2(_1401_),
    .ZN(_1402_));
 CLKBUF_X3 _3706_ (.A(_0882_),
    .Z(_1403_));
 MUX2_X1 _3707_ (.A(\mem[1][29] ),
    .B(\mem[5][29] ),
    .S(_1403_),
    .Z(_1404_));
 NOR2_X1 _3708_ (.A1(_1303_),
    .A2(_1404_),
    .ZN(_1405_));
 OAI33_X1 _3709_ (.A1(_1396_),
    .A2(_1398_),
    .A3(_1400_),
    .B1(_1402_),
    .B2(_1405_),
    .B3(_1379_),
    .ZN(_1406_));
 CLKBUF_X3 _3710_ (.A(_0881_),
    .Z(_1407_));
 MUX2_X1 _3711_ (.A(\mem[10][29] ),
    .B(\mem[14][29] ),
    .S(_1258_),
    .Z(_1408_));
 NOR2_X1 _3712_ (.A1(_1330_),
    .A2(_1408_),
    .ZN(_1409_));
 MUX2_X1 _3713_ (.A(\mem[11][29] ),
    .B(\mem[15][29] ),
    .S(_1216_),
    .Z(_1410_));
 NOR2_X1 _3714_ (.A1(_1333_),
    .A2(_1410_),
    .ZN(_1411_));
 MUX2_X1 _3715_ (.A(\mem[2][29] ),
    .B(\mem[6][29] ),
    .S(_1196_),
    .Z(_1412_));
 NOR2_X1 _3716_ (.A1(_1286_),
    .A2(_1412_),
    .ZN(_1413_));
 MUX2_X1 _3717_ (.A(\mem[3][29] ),
    .B(\mem[7][29] ),
    .S(_1313_),
    .Z(_1414_));
 NOR2_X1 _3718_ (.A1(_1265_),
    .A2(_1414_),
    .ZN(_1415_));
 OAI33_X1 _3719_ (.A1(_1407_),
    .A2(_1409_),
    .A3(_1411_),
    .B1(_1413_),
    .B2(_1415_),
    .B3(_1389_),
    .ZN(_1416_));
 OAI221_X1 _3720_ (.A(_1369_),
    .B1(_1406_),
    .B2(_1416_),
    .C1(_1365_),
    .C2(_1269_),
    .ZN(_1417_));
 NAND2_X1 _3721_ (.A1(\last_valid_data[29] ),
    .A2(_1392_),
    .ZN(_1418_));
 NAND2_X1 _3722_ (.A1(_1394_),
    .A2(\last_valid_data[29] ),
    .ZN(_1419_));
 OAI221_X1 _3723_ (.A(_1417_),
    .B1(_1418_),
    .B2(_1319_),
    .C1(_1419_),
    .C2(_1344_),
    .ZN(_0052_));
 MUX2_X1 _3724_ (.A(\mem[8][2] ),
    .B(\mem[12][2] ),
    .S(_1346_),
    .Z(_1420_));
 NOR2_X1 _3725_ (.A1(_1345_),
    .A2(_1420_),
    .ZN(_1421_));
 MUX2_X1 _3726_ (.A(\mem[9][2] ),
    .B(\mem[13][2] ),
    .S(_1297_),
    .Z(_1422_));
 NOR2_X1 _3727_ (.A1(_1372_),
    .A2(_1422_),
    .ZN(_1423_));
 MUX2_X1 _3728_ (.A(\mem[0][2] ),
    .B(\mem[4][2] ),
    .S(_1231_),
    .Z(_1424_));
 NOR2_X1 _3729_ (.A1(_1300_),
    .A2(_1424_),
    .ZN(_1425_));
 MUX2_X1 _3730_ (.A(\mem[1][2] ),
    .B(\mem[5][2] ),
    .S(_1403_),
    .Z(_1426_));
 NOR2_X1 _3731_ (.A1(_1303_),
    .A2(_1426_),
    .ZN(_1427_));
 OAI33_X1 _3732_ (.A1(_1396_),
    .A2(_1421_),
    .A3(_1423_),
    .B1(_1425_),
    .B2(_1427_),
    .B3(_1379_),
    .ZN(_1428_));
 MUX2_X1 _3733_ (.A(\mem[10][2] ),
    .B(\mem[14][2] ),
    .S(_1258_),
    .Z(_1429_));
 NOR2_X1 _3734_ (.A1(_1330_),
    .A2(_1429_),
    .ZN(_1430_));
 MUX2_X1 _3735_ (.A(\mem[11][2] ),
    .B(\mem[15][2] ),
    .S(_1216_),
    .Z(_1431_));
 NOR2_X1 _3736_ (.A1(_1333_),
    .A2(_1431_),
    .ZN(_1432_));
 BUF_X4 _3737_ (.A(_0882_),
    .Z(_1433_));
 MUX2_X1 _3738_ (.A(\mem[2][2] ),
    .B(\mem[6][2] ),
    .S(_1433_),
    .Z(_1434_));
 NOR2_X1 _3739_ (.A1(_1286_),
    .A2(_1434_),
    .ZN(_1435_));
 MUX2_X1 _3740_ (.A(\mem[3][2] ),
    .B(\mem[7][2] ),
    .S(_1313_),
    .Z(_1436_));
 NOR2_X1 _3741_ (.A1(_1265_),
    .A2(_1436_),
    .ZN(_1437_));
 OAI33_X1 _3742_ (.A1(_1407_),
    .A2(_1430_),
    .A3(_1432_),
    .B1(_1435_),
    .B2(_1437_),
    .B3(_1389_),
    .ZN(_1438_));
 OAI221_X1 _3743_ (.A(_1369_),
    .B1(_1428_),
    .B2(_1438_),
    .C1(_1365_),
    .C2(_1269_),
    .ZN(_1439_));
 NAND2_X1 _3744_ (.A1(\last_valid_data[2] ),
    .A2(_1392_),
    .ZN(_1440_));
 NAND2_X1 _3745_ (.A1(_1394_),
    .A2(\last_valid_data[2] ),
    .ZN(_1441_));
 OAI221_X1 _3746_ (.A(_1439_),
    .B1(_1440_),
    .B2(_1319_),
    .C1(_1441_),
    .C2(_1344_),
    .ZN(_0053_));
 MUX2_X1 _3747_ (.A(\mem[8][30] ),
    .B(\mem[12][30] ),
    .S(_1346_),
    .Z(_1442_));
 NOR2_X1 _3748_ (.A1(_1345_),
    .A2(_1442_),
    .ZN(_1443_));
 MUX2_X1 _3749_ (.A(\mem[9][30] ),
    .B(\mem[13][30] ),
    .S(_1297_),
    .Z(_1444_));
 NOR2_X1 _3750_ (.A1(_1372_),
    .A2(_1444_),
    .ZN(_1445_));
 MUX2_X1 _3751_ (.A(\mem[0][30] ),
    .B(\mem[4][30] ),
    .S(_1231_),
    .Z(_1446_));
 NOR2_X1 _3752_ (.A1(_1300_),
    .A2(_1446_),
    .ZN(_1447_));
 MUX2_X1 _3753_ (.A(\mem[1][30] ),
    .B(\mem[5][30] ),
    .S(_1403_),
    .Z(_1448_));
 NOR2_X1 _3754_ (.A1(_1303_),
    .A2(_1448_),
    .ZN(_1449_));
 OAI33_X1 _3755_ (.A1(_1396_),
    .A2(_1443_),
    .A3(_1445_),
    .B1(_1447_),
    .B2(_1449_),
    .B3(_1379_),
    .ZN(_1450_));
 MUX2_X1 _3756_ (.A(\mem[10][30] ),
    .B(\mem[14][30] ),
    .S(_1258_),
    .Z(_1451_));
 NOR2_X1 _3757_ (.A1(_1330_),
    .A2(_1451_),
    .ZN(_1452_));
 MUX2_X1 _3758_ (.A(\mem[11][30] ),
    .B(\mem[15][30] ),
    .S(_0936_),
    .Z(_1453_));
 NOR2_X1 _3759_ (.A1(_1333_),
    .A2(_1453_),
    .ZN(_1454_));
 MUX2_X1 _3760_ (.A(\mem[2][30] ),
    .B(\mem[6][30] ),
    .S(_1433_),
    .Z(_1455_));
 NOR2_X1 _3761_ (.A1(_1286_),
    .A2(_1455_),
    .ZN(_1456_));
 MUX2_X1 _3762_ (.A(\mem[3][30] ),
    .B(\mem[7][30] ),
    .S(_1313_),
    .Z(_1457_));
 NOR2_X1 _3763_ (.A1(_1265_),
    .A2(_1457_),
    .ZN(_1458_));
 OAI33_X1 _3764_ (.A1(_1407_),
    .A2(_1452_),
    .A3(_1454_),
    .B1(_1456_),
    .B2(_1458_),
    .B3(_1389_),
    .ZN(_1459_));
 OAI221_X1 _3765_ (.A(_1369_),
    .B1(_1450_),
    .B2(_1459_),
    .C1(_1365_),
    .C2(_1269_),
    .ZN(_1460_));
 NAND2_X1 _3766_ (.A1(\last_valid_data[30] ),
    .A2(_1392_),
    .ZN(_1461_));
 NAND2_X1 _3767_ (.A1(_1394_),
    .A2(\last_valid_data[30] ),
    .ZN(_1462_));
 OAI221_X1 _3768_ (.A(_1460_),
    .B1(_1461_),
    .B2(_1319_),
    .C1(_1462_),
    .C2(_1344_),
    .ZN(_0054_));
 MUX2_X1 _3769_ (.A(\mem[8][31] ),
    .B(\mem[12][31] ),
    .S(_1346_),
    .Z(_1463_));
 NOR2_X1 _3770_ (.A1(_1345_),
    .A2(_1463_),
    .ZN(_1464_));
 MUX2_X1 _3771_ (.A(\mem[9][31] ),
    .B(\mem[13][31] ),
    .S(_1297_),
    .Z(_1465_));
 NOR2_X1 _3772_ (.A1(_1372_),
    .A2(_1465_),
    .ZN(_1466_));
 MUX2_X1 _3773_ (.A(\mem[0][31] ),
    .B(\mem[4][31] ),
    .S(_0932_),
    .Z(_1467_));
 NOR2_X1 _3774_ (.A1(_1300_),
    .A2(_1467_),
    .ZN(_1468_));
 MUX2_X1 _3775_ (.A(\mem[1][31] ),
    .B(\mem[5][31] ),
    .S(_1403_),
    .Z(_1469_));
 NOR2_X1 _3776_ (.A1(_1303_),
    .A2(_1469_),
    .ZN(_1470_));
 OAI33_X1 _3777_ (.A1(_1396_),
    .A2(_1464_),
    .A3(_1466_),
    .B1(_1468_),
    .B2(_1470_),
    .B3(_1379_),
    .ZN(_1471_));
 MUX2_X1 _3778_ (.A(\mem[10][31] ),
    .B(\mem[14][31] ),
    .S(_1258_),
    .Z(_1472_));
 NOR2_X1 _3779_ (.A1(_1330_),
    .A2(_1472_),
    .ZN(_1473_));
 MUX2_X1 _3780_ (.A(\mem[11][31] ),
    .B(\mem[15][31] ),
    .S(_0936_),
    .Z(_1474_));
 NOR2_X1 _3781_ (.A1(_1333_),
    .A2(_1474_),
    .ZN(_1475_));
 MUX2_X1 _3782_ (.A(\mem[2][31] ),
    .B(\mem[6][31] ),
    .S(_1433_),
    .Z(_1476_));
 NOR2_X1 _3783_ (.A1(_1286_),
    .A2(_1476_),
    .ZN(_1477_));
 MUX2_X1 _3784_ (.A(\mem[3][31] ),
    .B(\mem[7][31] ),
    .S(_1313_),
    .Z(_1478_));
 NOR2_X1 _3785_ (.A1(_1265_),
    .A2(_1478_),
    .ZN(_1479_));
 OAI33_X1 _3786_ (.A1(_1407_),
    .A2(_1473_),
    .A3(_1475_),
    .B1(_1477_),
    .B2(_1479_),
    .B3(_1389_),
    .ZN(_1480_));
 OAI221_X1 _3787_ (.A(_1369_),
    .B1(_1471_),
    .B2(_1480_),
    .C1(_1365_),
    .C2(_1269_),
    .ZN(_1481_));
 NAND2_X1 _3788_ (.A1(\last_valid_data[31] ),
    .A2(_1392_),
    .ZN(_1482_));
 NAND2_X1 _3789_ (.A1(_1394_),
    .A2(\last_valid_data[31] ),
    .ZN(_1483_));
 OAI221_X1 _3790_ (.A(_1481_),
    .B1(_1482_),
    .B2(_1319_),
    .C1(_1483_),
    .C2(_1344_),
    .ZN(_0055_));
 MUX2_X1 _3791_ (.A(\mem[8][3] ),
    .B(\mem[12][3] ),
    .S(_1346_),
    .Z(_1484_));
 NOR2_X1 _3792_ (.A1(_1345_),
    .A2(_1484_),
    .ZN(_1485_));
 MUX2_X1 _3793_ (.A(\mem[9][3] ),
    .B(\mem[13][3] ),
    .S(_1297_),
    .Z(_1486_));
 NOR2_X1 _3794_ (.A1(_1372_),
    .A2(_1486_),
    .ZN(_1487_));
 MUX2_X1 _3795_ (.A(\mem[0][3] ),
    .B(\mem[4][3] ),
    .S(_0932_),
    .Z(_1488_));
 NOR2_X1 _3796_ (.A1(_1300_),
    .A2(_1488_),
    .ZN(_1489_));
 MUX2_X1 _3797_ (.A(\mem[1][3] ),
    .B(\mem[5][3] ),
    .S(_1403_),
    .Z(_1490_));
 NOR2_X1 _3798_ (.A1(_1303_),
    .A2(_1490_),
    .ZN(_1491_));
 OAI33_X1 _3799_ (.A1(_1396_),
    .A2(_1485_),
    .A3(_1487_),
    .B1(_1489_),
    .B2(_1491_),
    .B3(_1379_),
    .ZN(_1492_));
 MUX2_X1 _3800_ (.A(\mem[10][3] ),
    .B(\mem[14][3] ),
    .S(_0920_),
    .Z(_1493_));
 NOR2_X1 _3801_ (.A1(_1330_),
    .A2(_1493_),
    .ZN(_1494_));
 MUX2_X1 _3802_ (.A(\mem[11][3] ),
    .B(\mem[15][3] ),
    .S(_0936_),
    .Z(_1495_));
 NOR2_X1 _3803_ (.A1(_1333_),
    .A2(_1495_),
    .ZN(_1496_));
 MUX2_X1 _3804_ (.A(\mem[2][3] ),
    .B(\mem[6][3] ),
    .S(_1433_),
    .Z(_1497_));
 NOR2_X1 _3805_ (.A1(_1286_),
    .A2(_1497_),
    .ZN(_1498_));
 MUX2_X1 _3806_ (.A(\mem[3][3] ),
    .B(\mem[7][3] ),
    .S(_1313_),
    .Z(_1499_));
 NOR2_X1 _3807_ (.A1(_0871_),
    .A2(_1499_),
    .ZN(_1500_));
 OAI33_X1 _3808_ (.A1(_1407_),
    .A2(_1494_),
    .A3(_1496_),
    .B1(_1498_),
    .B2(_1500_),
    .B3(_1389_),
    .ZN(_1501_));
 OAI221_X1 _3809_ (.A(_1369_),
    .B1(_1492_),
    .B2(_1501_),
    .C1(_1365_),
    .C2(_0596_),
    .ZN(_1502_));
 NAND2_X1 _3810_ (.A1(\last_valid_data[3] ),
    .A2(_1392_),
    .ZN(_1503_));
 NAND2_X1 _3811_ (.A1(_1394_),
    .A2(\last_valid_data[3] ),
    .ZN(_1504_));
 OAI221_X1 _3812_ (.A(_1502_),
    .B1(_1503_),
    .B2(_1319_),
    .C1(_1504_),
    .C2(_1344_),
    .ZN(_0056_));
 MUX2_X1 _3813_ (.A(\mem[8][4] ),
    .B(\mem[12][4] ),
    .S(_1346_),
    .Z(_1505_));
 NOR2_X1 _3814_ (.A1(_1345_),
    .A2(_1505_),
    .ZN(_1506_));
 MUX2_X1 _3815_ (.A(\mem[9][4] ),
    .B(\mem[13][4] ),
    .S(_1297_),
    .Z(_1507_));
 NOR2_X1 _3816_ (.A1(_1372_),
    .A2(_1507_),
    .ZN(_1508_));
 MUX2_X1 _3817_ (.A(\mem[0][4] ),
    .B(\mem[4][4] ),
    .S(_0932_),
    .Z(_1509_));
 NOR2_X1 _3818_ (.A1(_1300_),
    .A2(_1509_),
    .ZN(_1510_));
 MUX2_X1 _3819_ (.A(\mem[1][4] ),
    .B(\mem[5][4] ),
    .S(_1403_),
    .Z(_1511_));
 NOR2_X1 _3820_ (.A1(_1303_),
    .A2(_1511_),
    .ZN(_1512_));
 OAI33_X1 _3821_ (.A1(_1396_),
    .A2(_1506_),
    .A3(_1508_),
    .B1(_1510_),
    .B2(_1512_),
    .B3(_1379_),
    .ZN(_1513_));
 MUX2_X1 _3822_ (.A(\mem[10][4] ),
    .B(\mem[14][4] ),
    .S(_0920_),
    .Z(_1514_));
 NOR2_X1 _3823_ (.A1(_1330_),
    .A2(_1514_),
    .ZN(_1515_));
 MUX2_X1 _3824_ (.A(\mem[11][4] ),
    .B(\mem[15][4] ),
    .S(_0936_),
    .Z(_1516_));
 NOR2_X1 _3825_ (.A1(_1333_),
    .A2(_1516_),
    .ZN(_1517_));
 MUX2_X1 _3826_ (.A(\mem[2][4] ),
    .B(\mem[6][4] ),
    .S(_1433_),
    .Z(_1518_));
 NOR2_X1 _3827_ (.A1(_0863_),
    .A2(_1518_),
    .ZN(_1519_));
 MUX2_X1 _3828_ (.A(\mem[3][4] ),
    .B(\mem[7][4] ),
    .S(_1313_),
    .Z(_1520_));
 NOR2_X1 _3829_ (.A1(_0871_),
    .A2(_1520_),
    .ZN(_1521_));
 OAI33_X1 _3830_ (.A1(_1407_),
    .A2(_1515_),
    .A3(_1517_),
    .B1(_1519_),
    .B2(_1521_),
    .B3(_1389_),
    .ZN(_1522_));
 OAI221_X1 _3831_ (.A(_1369_),
    .B1(_1513_),
    .B2(_1522_),
    .C1(_1365_),
    .C2(_0596_),
    .ZN(_1523_));
 NAND2_X1 _3832_ (.A1(\last_valid_data[4] ),
    .A2(_1392_),
    .ZN(_1524_));
 NAND2_X1 _3833_ (.A1(_1394_),
    .A2(\last_valid_data[4] ),
    .ZN(_1525_));
 OAI221_X1 _3834_ (.A(_1523_),
    .B1(_1524_),
    .B2(_1319_),
    .C1(_1525_),
    .C2(_1344_),
    .ZN(_0057_));
 MUX2_X1 _3835_ (.A(\mem[8][5] ),
    .B(\mem[12][5] ),
    .S(_1346_),
    .Z(_1526_));
 NOR2_X1 _3836_ (.A1(_1345_),
    .A2(_1526_),
    .ZN(_1527_));
 MUX2_X1 _3837_ (.A(\mem[9][5] ),
    .B(\mem[13][5] ),
    .S(_0895_),
    .Z(_1528_));
 NOR2_X1 _3838_ (.A1(_1372_),
    .A2(_1528_),
    .ZN(_1529_));
 MUX2_X1 _3839_ (.A(\mem[0][5] ),
    .B(\mem[4][5] ),
    .S(_0932_),
    .Z(_1530_));
 NOR2_X1 _3840_ (.A1(_0935_),
    .A2(_1530_),
    .ZN(_1531_));
 MUX2_X1 _3841_ (.A(\mem[1][5] ),
    .B(\mem[5][5] ),
    .S(_1403_),
    .Z(_1532_));
 NOR2_X1 _3842_ (.A1(_0887_),
    .A2(_1532_),
    .ZN(_1533_));
 OAI33_X1 _3843_ (.A1(_1396_),
    .A2(_1527_),
    .A3(_1529_),
    .B1(_1531_),
    .B2(_1533_),
    .B3(_1379_),
    .ZN(_1534_));
 MUX2_X1 _3844_ (.A(\mem[10][5] ),
    .B(\mem[14][5] ),
    .S(_0920_),
    .Z(_1535_));
 NOR2_X1 _3845_ (.A1(_1330_),
    .A2(_1535_),
    .ZN(_1536_));
 MUX2_X1 _3846_ (.A(\mem[11][5] ),
    .B(\mem[15][5] ),
    .S(_0936_),
    .Z(_1537_));
 NOR2_X1 _3847_ (.A1(_1333_),
    .A2(_1537_),
    .ZN(_1538_));
 MUX2_X1 _3848_ (.A(\mem[2][5] ),
    .B(\mem[6][5] ),
    .S(_1433_),
    .Z(_1539_));
 NOR2_X1 _3849_ (.A1(_0863_),
    .A2(_1539_),
    .ZN(_1540_));
 MUX2_X1 _3850_ (.A(\mem[3][5] ),
    .B(\mem[7][5] ),
    .S(_0866_),
    .Z(_1541_));
 NOR2_X1 _3851_ (.A1(_0871_),
    .A2(_1541_),
    .ZN(_1542_));
 OAI33_X1 _3852_ (.A1(_1407_),
    .A2(_1536_),
    .A3(_1538_),
    .B1(_1540_),
    .B2(_1542_),
    .B3(_1389_),
    .ZN(_1543_));
 OAI221_X1 _3853_ (.A(_1369_),
    .B1(_1534_),
    .B2(_1543_),
    .C1(_1365_),
    .C2(_0596_),
    .ZN(_1544_));
 NAND2_X1 _3854_ (.A1(\last_valid_data[5] ),
    .A2(_1392_),
    .ZN(_1545_));
 NAND2_X1 _3855_ (.A1(_1394_),
    .A2(\last_valid_data[5] ),
    .ZN(_1546_));
 OAI221_X1 _3856_ (.A(_1544_),
    .B1(_1545_),
    .B2(net68),
    .C1(_1546_),
    .C2(_1344_),
    .ZN(_0058_));
 MUX2_X1 _3857_ (.A(\mem[8][6] ),
    .B(\mem[12][6] ),
    .S(_1346_),
    .Z(_1547_));
 NOR2_X1 _3858_ (.A1(_1345_),
    .A2(_1547_),
    .ZN(_1548_));
 MUX2_X1 _3859_ (.A(\mem[9][6] ),
    .B(\mem[13][6] ),
    .S(_0895_),
    .Z(_1549_));
 NOR2_X1 _3860_ (.A1(_1372_),
    .A2(_1549_),
    .ZN(_1550_));
 MUX2_X1 _3861_ (.A(\mem[0][6] ),
    .B(\mem[4][6] ),
    .S(_0932_),
    .Z(_1551_));
 NOR2_X1 _3862_ (.A1(_0935_),
    .A2(_1551_),
    .ZN(_1552_));
 MUX2_X1 _3863_ (.A(\mem[1][6] ),
    .B(\mem[5][6] ),
    .S(_1403_),
    .Z(_1553_));
 NOR2_X1 _3864_ (.A1(_0887_),
    .A2(_1553_),
    .ZN(_1554_));
 OAI33_X1 _3865_ (.A1(_1396_),
    .A2(_1548_),
    .A3(_1550_),
    .B1(_1552_),
    .B2(_1554_),
    .B3(_1379_),
    .ZN(_1555_));
 MUX2_X1 _3866_ (.A(\mem[10][6] ),
    .B(\mem[14][6] ),
    .S(_0920_),
    .Z(_1556_));
 NOR2_X1 _3867_ (.A1(_0919_),
    .A2(_1556_),
    .ZN(_1557_));
 MUX2_X1 _3868_ (.A(\mem[11][6] ),
    .B(\mem[15][6] ),
    .S(_0936_),
    .Z(_1558_));
 NOR2_X1 _3869_ (.A1(_0923_),
    .A2(_1558_),
    .ZN(_1559_));
 MUX2_X1 _3870_ (.A(\mem[2][6] ),
    .B(\mem[6][6] ),
    .S(_1433_),
    .Z(_1560_));
 NOR2_X1 _3871_ (.A1(_0863_),
    .A2(_1560_),
    .ZN(_1561_));
 MUX2_X1 _3872_ (.A(\mem[3][6] ),
    .B(\mem[7][6] ),
    .S(_0866_),
    .Z(_1562_));
 NOR2_X1 _3873_ (.A1(_0871_),
    .A2(_1562_),
    .ZN(_1563_));
 OAI33_X1 _3874_ (.A1(_1407_),
    .A2(_1557_),
    .A3(_1559_),
    .B1(_1561_),
    .B2(_1563_),
    .B3(_1389_),
    .ZN(_1564_));
 OAI221_X1 _3875_ (.A(_1369_),
    .B1(_1555_),
    .B2(_1564_),
    .C1(_1365_),
    .C2(_0596_),
    .ZN(_1565_));
 NAND2_X1 _3876_ (.A1(\last_valid_data[6] ),
    .A2(_1392_),
    .ZN(_1566_));
 NAND2_X1 _3877_ (.A1(_1394_),
    .A2(\last_valid_data[6] ),
    .ZN(_1567_));
 OAI221_X1 _3878_ (.A(_1565_),
    .B1(_1566_),
    .B2(net68),
    .C1(_1567_),
    .C2(_0772_),
    .ZN(_0059_));
 MUX2_X1 _3879_ (.A(\mem[8][7] ),
    .B(\mem[12][7] ),
    .S(_0873_),
    .Z(_1568_));
 NOR2_X1 _3880_ (.A1(_0929_),
    .A2(_1568_),
    .ZN(_1569_));
 MUX2_X1 _3881_ (.A(\mem[9][7] ),
    .B(\mem[13][7] ),
    .S(_0895_),
    .Z(_1570_));
 NOR2_X1 _3882_ (.A1(_1372_),
    .A2(_1570_),
    .ZN(_1571_));
 MUX2_X1 _3883_ (.A(\mem[0][7] ),
    .B(\mem[4][7] ),
    .S(_0932_),
    .Z(_1572_));
 NOR2_X1 _3884_ (.A1(_0935_),
    .A2(_1572_),
    .ZN(_1573_));
 MUX2_X1 _3885_ (.A(\mem[1][7] ),
    .B(\mem[5][7] ),
    .S(_1403_),
    .Z(_1574_));
 NOR2_X1 _3886_ (.A1(_0887_),
    .A2(_1574_),
    .ZN(_1575_));
 OAI33_X1 _3887_ (.A1(_1396_),
    .A2(_1569_),
    .A3(_1571_),
    .B1(_1573_),
    .B2(_1575_),
    .B3(_1379_),
    .ZN(_1576_));
 MUX2_X1 _3888_ (.A(\mem[10][7] ),
    .B(\mem[14][7] ),
    .S(_0920_),
    .Z(_1577_));
 NOR2_X1 _3889_ (.A1(_0919_),
    .A2(_1577_),
    .ZN(_1578_));
 MUX2_X1 _3890_ (.A(\mem[11][7] ),
    .B(\mem[15][7] ),
    .S(_0936_),
    .Z(_1579_));
 NOR2_X1 _3891_ (.A1(_0923_),
    .A2(_1579_),
    .ZN(_1580_));
 MUX2_X1 _3892_ (.A(\mem[2][7] ),
    .B(\mem[6][7] ),
    .S(_1433_),
    .Z(_1581_));
 NOR2_X1 _3893_ (.A1(_0863_),
    .A2(_1581_),
    .ZN(_1582_));
 MUX2_X1 _3894_ (.A(\mem[3][7] ),
    .B(\mem[7][7] ),
    .S(_0866_),
    .Z(_1583_));
 NOR2_X1 _3895_ (.A1(_0871_),
    .A2(_1583_),
    .ZN(_1584_));
 OAI33_X1 _3896_ (.A1(_1407_),
    .A2(_1578_),
    .A3(_1580_),
    .B1(_1582_),
    .B2(_1584_),
    .B3(_1389_),
    .ZN(_1585_));
 OAI221_X1 _3897_ (.A(_1369_),
    .B1(_1576_),
    .B2(_1585_),
    .C1(_0798_),
    .C2(_0596_),
    .ZN(_1586_));
 NAND2_X1 _3898_ (.A1(\last_valid_data[7] ),
    .A2(_1392_),
    .ZN(_1587_));
 NAND2_X1 _3899_ (.A1(_1394_),
    .A2(\last_valid_data[7] ),
    .ZN(_1588_));
 OAI221_X1 _3900_ (.A(_1586_),
    .B1(_1587_),
    .B2(net68),
    .C1(_1588_),
    .C2(_0772_),
    .ZN(_0060_));
 MUX2_X1 _3901_ (.A(\mem[8][8] ),
    .B(\mem[12][8] ),
    .S(_0873_),
    .Z(_1589_));
 NOR2_X1 _3902_ (.A1(_0929_),
    .A2(_1589_),
    .ZN(_1590_));
 MUX2_X1 _3903_ (.A(\mem[9][8] ),
    .B(\mem[13][8] ),
    .S(_0895_),
    .Z(_1591_));
 NOR2_X1 _3904_ (.A1(_0893_),
    .A2(_1591_),
    .ZN(_1592_));
 MUX2_X1 _3905_ (.A(\mem[0][8] ),
    .B(\mem[4][8] ),
    .S(_0932_),
    .Z(_1593_));
 NOR2_X1 _3906_ (.A1(_0935_),
    .A2(_1593_),
    .ZN(_1594_));
 MUX2_X1 _3907_ (.A(\mem[1][8] ),
    .B(\mem[5][8] ),
    .S(_1403_),
    .Z(_1595_));
 NOR2_X1 _3908_ (.A1(_0887_),
    .A2(_1595_),
    .ZN(_1596_));
 OAI33_X1 _3909_ (.A1(_1396_),
    .A2(_1590_),
    .A3(_1592_),
    .B1(_1594_),
    .B2(_1596_),
    .B3(_0899_),
    .ZN(_1597_));
 MUX2_X1 _3910_ (.A(\mem[10][8] ),
    .B(\mem[14][8] ),
    .S(_0920_),
    .Z(_1598_));
 NOR2_X1 _3911_ (.A1(_0919_),
    .A2(_1598_),
    .ZN(_1599_));
 MUX2_X1 _3912_ (.A(\mem[11][8] ),
    .B(\mem[15][8] ),
    .S(_0936_),
    .Z(_1600_));
 NOR2_X1 _3913_ (.A1(_0923_),
    .A2(_1600_),
    .ZN(_1601_));
 MUX2_X1 _3914_ (.A(\mem[2][8] ),
    .B(\mem[6][8] ),
    .S(_1433_),
    .Z(_1602_));
 NOR2_X1 _3915_ (.A1(_0863_),
    .A2(_1602_),
    .ZN(_1603_));
 MUX2_X1 _3916_ (.A(\mem[3][8] ),
    .B(\mem[7][8] ),
    .S(_0866_),
    .Z(_1604_));
 NOR2_X1 _3917_ (.A1(_0871_),
    .A2(_1604_),
    .ZN(_1605_));
 OAI33_X1 _3918_ (.A1(_1407_),
    .A2(_1599_),
    .A3(_1601_),
    .B1(_1603_),
    .B2(_1605_),
    .B3(_0879_),
    .ZN(_1606_));
 OAI221_X1 _3919_ (.A(_0860_),
    .B1(_1597_),
    .B2(_1606_),
    .C1(_0798_),
    .C2(_0596_),
    .ZN(_1607_));
 NAND2_X1 _3920_ (.A1(\last_valid_data[8] ),
    .A2(_0769_),
    .ZN(_1608_));
 NAND2_X1 _3921_ (.A1(_0859_),
    .A2(\last_valid_data[8] ),
    .ZN(_1609_));
 OAI221_X1 _3922_ (.A(_1607_),
    .B1(_1608_),
    .B2(net68),
    .C1(_1609_),
    .C2(_0772_),
    .ZN(_0061_));
 MUX2_X1 _3923_ (.A(\mem[8][9] ),
    .B(\mem[12][9] ),
    .S(_0873_),
    .Z(_1610_));
 NOR2_X1 _3924_ (.A1(_0929_),
    .A2(_1610_),
    .ZN(_1611_));
 MUX2_X1 _3925_ (.A(\mem[9][9] ),
    .B(\mem[13][9] ),
    .S(_0895_),
    .Z(_1612_));
 NOR2_X1 _3926_ (.A1(_0893_),
    .A2(_1612_),
    .ZN(_1613_));
 MUX2_X1 _3927_ (.A(\mem[0][9] ),
    .B(\mem[4][9] ),
    .S(_0932_),
    .Z(_1614_));
 NOR2_X1 _3928_ (.A1(_0935_),
    .A2(_1614_),
    .ZN(_1615_));
 MUX2_X1 _3929_ (.A(\mem[1][9] ),
    .B(\mem[5][9] ),
    .S(_0883_),
    .Z(_1616_));
 NOR2_X1 _3930_ (.A1(_0887_),
    .A2(_1616_),
    .ZN(_1617_));
 OAI33_X1 _3931_ (.A1(_0901_),
    .A2(_1611_),
    .A3(_1613_),
    .B1(_1615_),
    .B2(_1617_),
    .B3(_0899_),
    .ZN(_1618_));
 MUX2_X1 _3932_ (.A(\mem[10][9] ),
    .B(\mem[14][9] ),
    .S(_0920_),
    .Z(_1619_));
 NOR2_X1 _3933_ (.A1(_0919_),
    .A2(_1619_),
    .ZN(_1620_));
 MUX2_X1 _3934_ (.A(\mem[11][9] ),
    .B(\mem[15][9] ),
    .S(_0936_),
    .Z(_1621_));
 NOR2_X1 _3935_ (.A1(_0923_),
    .A2(_1621_),
    .ZN(_1622_));
 MUX2_X1 _3936_ (.A(\mem[2][9] ),
    .B(\mem[6][9] ),
    .S(_1433_),
    .Z(_1623_));
 NOR2_X1 _3937_ (.A1(_0863_),
    .A2(_1623_),
    .ZN(_1624_));
 MUX2_X1 _3938_ (.A(\mem[3][9] ),
    .B(\mem[7][9] ),
    .S(_0866_),
    .Z(_1625_));
 NOR2_X1 _3939_ (.A1(_0871_),
    .A2(_1625_),
    .ZN(_1626_));
 OAI33_X1 _3940_ (.A1(_0881_),
    .A2(_1620_),
    .A3(_1622_),
    .B1(_1624_),
    .B2(_1626_),
    .B3(_0879_),
    .ZN(_1627_));
 OAI221_X1 _3941_ (.A(_0860_),
    .B1(_1618_),
    .B2(_1627_),
    .C1(_0798_),
    .C2(_0596_),
    .ZN(_1628_));
 NAND2_X1 _3942_ (.A1(\last_valid_data[9] ),
    .A2(_0769_),
    .ZN(_1629_));
 NAND2_X1 _3943_ (.A1(_0859_),
    .A2(\last_valid_data[9] ),
    .ZN(_1630_));
 OAI221_X1 _3944_ (.A(_1628_),
    .B1(_1629_),
    .B2(net68),
    .C1(_1630_),
    .C2(_0772_),
    .ZN(_0062_));
 BUF_X2 _3945_ (.A(last_valid_data_available),
    .Z(_1631_));
 CLKBUF_X3 _3946_ (.A(_1631_),
    .Z(_1632_));
 INV_X1 _3947_ (.A(_1632_),
    .ZN(_1633_));
 AOI21_X1 _3948_ (.A(_0856_),
    .B1(_0766_),
    .B2(_1633_),
    .ZN(_0063_));
 AND2_X1 _3949_ (.A1(_0006_),
    .A2(_0828_),
    .ZN(_1634_));
 MUX2_X1 _3950_ (.A(_1634_),
    .B(_0765_),
    .S(_0766_),
    .Z(_0576_));
 AND2_X1 _3951_ (.A1(\rd_ptr[4] ),
    .A2(_0828_),
    .ZN(_1635_));
 NOR2_X1 _3952_ (.A1(\rd_ptr[4] ),
    .A2(_0830_),
    .ZN(_1636_));
 NAND4_X1 _3953_ (.A1(_0608_),
    .A2(_2310_),
    .A3(\rd_ptr[2] ),
    .A4(\rd_ptr[3] ),
    .ZN(_1637_));
 AOI21_X1 _3954_ (.A(_1637_),
    .B1(_0602_),
    .B2(_0593_),
    .ZN(_1638_));
 MUX2_X1 _3955_ (.A(_1635_),
    .B(_1636_),
    .S(_1638_),
    .Z(_0577_));
 AND2_X1 _3956_ (.A1(\wr_ptr[0] ),
    .A2(_0828_),
    .ZN(_1639_));
 AND2_X1 _3957_ (.A1(_0004_),
    .A2(_0769_),
    .ZN(_1640_));
 AOI21_X1 _3958_ (.A(_0614_),
    .B1(_0595_),
    .B2(_0601_),
    .ZN(_1641_));
 MUX2_X1 _3959_ (.A(_1639_),
    .B(_1640_),
    .S(_1641_),
    .Z(_0578_));
 AND2_X1 _3960_ (.A1(\wr_ptr[1] ),
    .A2(_0828_),
    .ZN(_1642_));
 AND2_X1 _3961_ (.A1(_0005_),
    .A2(_0767_),
    .ZN(_1643_));
 MUX2_X1 _3962_ (.A(_1642_),
    .B(_1643_),
    .S(_1641_),
    .Z(_0579_));
 NOR2_X1 _3963_ (.A1(_0686_),
    .A2(_0763_),
    .ZN(_1644_));
 NOR2_X1 _3964_ (.A1(_0616_),
    .A2(_0830_),
    .ZN(_1645_));
 NAND2_X1 _3965_ (.A1(_0613_),
    .A2(_0693_),
    .ZN(_1646_));
 AOI21_X1 _3966_ (.A(_1646_),
    .B1(_0602_),
    .B2(_0797_),
    .ZN(_1647_));
 MUX2_X1 _3967_ (.A(_1644_),
    .B(_1645_),
    .S(_1647_),
    .Z(_0580_));
 AND2_X1 _3968_ (.A1(_0615_),
    .A2(_0828_),
    .ZN(_1648_));
 NOR2_X1 _3969_ (.A1(_0615_),
    .A2(_0830_),
    .ZN(_1649_));
 NAND4_X1 _3970_ (.A1(_0613_),
    .A2(_0616_),
    .A3(\wr_ptr[1] ),
    .A4(\wr_ptr[0] ),
    .ZN(_1650_));
 AOI21_X1 _3971_ (.A(_1650_),
    .B1(_0602_),
    .B2(_0595_),
    .ZN(_1651_));
 MUX2_X1 _3972_ (.A(_1648_),
    .B(_1649_),
    .S(_1651_),
    .Z(_0581_));
 AND2_X1 _3973_ (.A1(\wr_ptr[4] ),
    .A2(_0761_),
    .ZN(_1652_));
 NOR2_X1 _3974_ (.A1(\wr_ptr[4] ),
    .A2(_0830_),
    .ZN(_1653_));
 AOI21_X1 _3975_ (.A(_0713_),
    .B1(_0602_),
    .B2(_0595_),
    .ZN(_1654_));
 MUX2_X1 _3976_ (.A(_1652_),
    .B(_1653_),
    .S(_1654_),
    .Z(_0582_));
 XOR2_X1 _3977_ (.A(_2321_),
    .B(_0598_),
    .Z(_1655_));
 NOR4_X1 _3978_ (.A1(net6),
    .A2(net7),
    .A3(_0597_),
    .A4(_1655_),
    .ZN(net2));
 NAND2_X1 _3979_ (.A1(_0598_),
    .A2(net6),
    .ZN(_1656_));
 OAI21_X1 _3980_ (.A(_0593_),
    .B1(_1656_),
    .B2(_0587_),
    .ZN(net3));
 NOR2_X1 _3981_ (.A1(_0614_),
    .A2(net63),
    .ZN(net28));
 BUF_X4 _3982_ (.A(_0798_),
    .Z(_1657_));
 OAI22_X1 _3983_ (.A1(net8),
    .A2(_1657_),
    .B1(_0906_),
    .B2(_0890_),
    .ZN(_1658_));
 NAND2_X1 _3984_ (.A1(_1632_),
    .A2(\last_valid_data[0] ),
    .ZN(_1659_));
 OAI21_X1 _3985_ (.A(_1658_),
    .B1(_1659_),
    .B2(net61),
    .ZN(net29));
 OAI22_X1 _3986_ (.A1(net8),
    .A2(_1657_),
    .B1(_0927_),
    .B2(_0941_),
    .ZN(_1660_));
 NAND2_X1 _3987_ (.A1(_1632_),
    .A2(\last_valid_data[10] ),
    .ZN(_1661_));
 OAI21_X1 _3988_ (.A(_1660_),
    .B1(_1661_),
    .B2(net61),
    .ZN(net30));
 OAI22_X1 _3989_ (.A1(net8),
    .A2(_1657_),
    .B1(_0954_),
    .B2(_0964_),
    .ZN(_1662_));
 NAND2_X1 _3990_ (.A1(_1632_),
    .A2(\last_valid_data[11] ),
    .ZN(_1663_));
 OAI21_X1 _3991_ (.A(_1662_),
    .B1(_1663_),
    .B2(net61),
    .ZN(net31));
 OAI22_X1 _3992_ (.A1(net8),
    .A2(_1657_),
    .B1(_0976_),
    .B2(_0986_),
    .ZN(_1664_));
 NAND2_X1 _3993_ (.A1(_1632_),
    .A2(\last_valid_data[12] ),
    .ZN(_1665_));
 OAI21_X1 _3994_ (.A(_1664_),
    .B1(_1665_),
    .B2(net61),
    .ZN(net32));
 OAI22_X1 _3995_ (.A1(net8),
    .A2(_1657_),
    .B1(_0999_),
    .B2(_1008_),
    .ZN(_1666_));
 NAND2_X1 _3996_ (.A1(_1632_),
    .A2(\last_valid_data[13] ),
    .ZN(_1667_));
 OAI21_X1 _3997_ (.A(_1666_),
    .B1(_1667_),
    .B2(net61),
    .ZN(net33));
 OAI22_X1 _3998_ (.A1(net8),
    .A2(_1657_),
    .B1(_1020_),
    .B2(_1031_),
    .ZN(_1668_));
 NAND2_X1 _3999_ (.A1(_1632_),
    .A2(\last_valid_data[14] ),
    .ZN(_1669_));
 OAI21_X1 _4000_ (.A(_1668_),
    .B1(_1669_),
    .B2(net61),
    .ZN(net34));
 OAI22_X1 _4001_ (.A1(net8),
    .A2(_1657_),
    .B1(_1044_),
    .B2(_1054_),
    .ZN(_1670_));
 NAND2_X1 _4002_ (.A1(_1632_),
    .A2(\last_valid_data[15] ),
    .ZN(_1671_));
 OAI21_X1 _4003_ (.A(_1670_),
    .B1(_1671_),
    .B2(net61),
    .ZN(net35));
 OAI22_X1 _4004_ (.A1(net8),
    .A2(_1657_),
    .B1(_1069_),
    .B2(_1079_),
    .ZN(_1672_));
 NAND2_X1 _4005_ (.A1(_1632_),
    .A2(\last_valid_data[16] ),
    .ZN(_1673_));
 OAI21_X1 _4006_ (.A(_1672_),
    .B1(_1673_),
    .B2(net61),
    .ZN(net36));
 OAI22_X1 _4007_ (.A1(net8),
    .A2(_1657_),
    .B1(_1092_),
    .B2(_1103_),
    .ZN(_1674_));
 NAND2_X1 _4008_ (.A1(_1632_),
    .A2(\last_valid_data[17] ),
    .ZN(_1675_));
 OAI21_X1 _4009_ (.A(_1674_),
    .B1(_1675_),
    .B2(net61),
    .ZN(net37));
 CLKBUF_X3 _4010_ (.A(_0596_),
    .Z(_1676_));
 OAI22_X1 _4011_ (.A1(_1676_),
    .A2(_1657_),
    .B1(_1118_),
    .B2(_1127_),
    .ZN(_1677_));
 CLKBUF_X3 _4012_ (.A(_1631_),
    .Z(_1678_));
 NAND2_X1 _4013_ (.A1(_1678_),
    .A2(\last_valid_data[18] ),
    .ZN(_1679_));
 BUF_X32 _4014_ (.A(_0607_),
    .Z(_1680_));
 OAI21_X2 _4015_ (.A(_1677_),
    .B1(_1679_),
    .B2(_1680_),
    .ZN(net38));
 BUF_X8 _4016_ (.A(_0798_),
    .Z(_1681_));
 OAI22_X2 _4017_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1143_),
    .B2(_1153_),
    .ZN(_1682_));
 NAND2_X1 _4018_ (.A1(_1678_),
    .A2(\last_valid_data[19] ),
    .ZN(_1683_));
 OAI21_X2 _4019_ (.A(_1682_),
    .B1(_1683_),
    .B2(_1680_),
    .ZN(net39));
 OAI22_X2 _4020_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1169_),
    .B2(_1179_),
    .ZN(_1684_));
 NAND2_X1 _4021_ (.A1(_1678_),
    .A2(\last_valid_data[1] ),
    .ZN(_1685_));
 OAI21_X2 _4022_ (.A(_1684_),
    .B1(_1685_),
    .B2(net67),
    .ZN(net40));
 OAI22_X2 _4023_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1191_),
    .B2(_1201_),
    .ZN(_1686_));
 NAND2_X1 _4024_ (.A1(_1678_),
    .A2(\last_valid_data[20] ),
    .ZN(_1687_));
 OAI21_X2 _4025_ (.A(_1686_),
    .B1(_1687_),
    .B2(net67),
    .ZN(net41));
 OAI22_X2 _4026_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1213_),
    .B2(_1223_),
    .ZN(_1688_));
 NAND2_X1 _4027_ (.A1(_1678_),
    .A2(\last_valid_data[21] ),
    .ZN(_1689_));
 OAI21_X2 _4028_ (.A(_1688_),
    .B1(_1689_),
    .B2(net67),
    .ZN(net42));
 OAI22_X2 _4029_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1236_),
    .B2(_1245_),
    .ZN(_1690_));
 NAND2_X1 _4030_ (.A1(_1678_),
    .A2(\last_valid_data[22] ),
    .ZN(_1691_));
 OAI21_X2 _4031_ (.A(_1690_),
    .B1(_1691_),
    .B2(net67),
    .ZN(net43));
 OAI22_X2 _4032_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1257_),
    .B2(_1268_),
    .ZN(_1692_));
 NAND2_X1 _4033_ (.A1(_1678_),
    .A2(\last_valid_data[23] ),
    .ZN(_1693_));
 OAI21_X2 _4034_ (.A(_1692_),
    .B1(_1693_),
    .B2(_1680_),
    .ZN(net44));
 OAI22_X2 _4035_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1281_),
    .B2(_1291_),
    .ZN(_1694_));
 NAND2_X1 _4036_ (.A1(_1678_),
    .A2(\last_valid_data[24] ),
    .ZN(_1695_));
 OAI21_X2 _4037_ (.A(_1694_),
    .B1(_1695_),
    .B2(net67),
    .ZN(net45));
 OAI22_X2 _4038_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1306_),
    .B2(_1316_),
    .ZN(_1696_));
 NAND2_X1 _4039_ (.A1(_1678_),
    .A2(\last_valid_data[25] ),
    .ZN(_1697_));
 OAI21_X2 _4040_ (.A(_1696_),
    .B1(_1697_),
    .B2(_1680_),
    .ZN(net46));
 OAI22_X2 _4041_ (.A1(_1676_),
    .A2(_1681_),
    .B1(_1329_),
    .B2(_1340_),
    .ZN(_1698_));
 NAND2_X1 _4042_ (.A1(_1678_),
    .A2(\last_valid_data[26] ),
    .ZN(_1699_));
 OAI21_X2 _4043_ (.A(_1698_),
    .B1(_1699_),
    .B2(_1680_),
    .ZN(net47));
 CLKBUF_X3 _4044_ (.A(_0596_),
    .Z(_1700_));
 OAI22_X2 _4045_ (.A1(_1700_),
    .A2(_1681_),
    .B1(_1355_),
    .B2(_1364_),
    .ZN(_1701_));
 CLKBUF_X3 _4046_ (.A(_1631_),
    .Z(_1702_));
 NAND2_X1 _4047_ (.A1(_1702_),
    .A2(\last_valid_data[27] ),
    .ZN(_1703_));
 BUF_X32 _4048_ (.A(_0607_),
    .Z(_1704_));
 OAI21_X4 _4049_ (.A(_1701_),
    .B1(_1703_),
    .B2(net66),
    .ZN(net48));
 BUF_X8 _4050_ (.A(_0798_),
    .Z(_1705_));
 OAI22_X2 _4051_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1380_),
    .B2(_1390_),
    .ZN(_1706_));
 NAND2_X1 _4052_ (.A1(_1702_),
    .A2(\last_valid_data[28] ),
    .ZN(_1707_));
 OAI21_X2 _4053_ (.A(_1706_),
    .B1(_1707_),
    .B2(net66),
    .ZN(net49));
 OAI22_X2 _4054_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1406_),
    .B2(_1416_),
    .ZN(_1708_));
 NAND2_X1 _4055_ (.A1(_1702_),
    .A2(\last_valid_data[29] ),
    .ZN(_1709_));
 OAI21_X4 _4056_ (.A(_1708_),
    .B1(_1709_),
    .B2(_1704_),
    .ZN(net50));
 OAI22_X2 _4057_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1428_),
    .B2(_1438_),
    .ZN(_1710_));
 NAND2_X1 _4058_ (.A1(_1702_),
    .A2(\last_valid_data[2] ),
    .ZN(_1711_));
 OAI21_X4 _4059_ (.A(_1710_),
    .B1(_1711_),
    .B2(_1704_),
    .ZN(net51));
 OAI22_X2 _4060_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1450_),
    .B2(_1459_),
    .ZN(_1712_));
 NAND2_X1 _4061_ (.A1(_1702_),
    .A2(\last_valid_data[30] ),
    .ZN(_1713_));
 OAI21_X4 _4062_ (.A(_1712_),
    .B1(_1713_),
    .B2(_1704_),
    .ZN(net52));
 OAI22_X2 _4063_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1471_),
    .B2(_1480_),
    .ZN(_1714_));
 NAND2_X1 _4064_ (.A1(_1702_),
    .A2(\last_valid_data[31] ),
    .ZN(_1715_));
 OAI21_X4 _4065_ (.A(_1714_),
    .B1(_1715_),
    .B2(_1704_),
    .ZN(net53));
 OAI22_X2 _4066_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1492_),
    .B2(_1501_),
    .ZN(_1716_));
 NAND2_X1 _4067_ (.A1(_1702_),
    .A2(\last_valid_data[3] ),
    .ZN(_1717_));
 OAI21_X4 _4068_ (.A(_1716_),
    .B1(_1717_),
    .B2(_1704_),
    .ZN(net54));
 OAI22_X4 _4069_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1513_),
    .B2(_1522_),
    .ZN(_1718_));
 NAND2_X1 _4070_ (.A1(_1702_),
    .A2(\last_valid_data[4] ),
    .ZN(_1719_));
 OAI21_X4 _4071_ (.A(_1718_),
    .B1(_1719_),
    .B2(net66),
    .ZN(net55));
 OAI22_X4 _4072_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1534_),
    .B2(_1543_),
    .ZN(_1720_));
 NAND2_X1 _4073_ (.A1(_1702_),
    .A2(\last_valid_data[5] ),
    .ZN(_1721_));
 OAI21_X4 _4074_ (.A(_1720_),
    .B1(net66),
    .B2(_1721_),
    .ZN(net56));
 OAI22_X4 _4075_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1555_),
    .B2(_1564_),
    .ZN(_1722_));
 NAND2_X1 _4076_ (.A1(_1702_),
    .A2(\last_valid_data[6] ),
    .ZN(_1723_));
 OAI21_X4 _4077_ (.A(_1722_),
    .B1(net66),
    .B2(_1723_),
    .ZN(net57));
 OAI22_X2 _4078_ (.A1(_0597_),
    .A2(_1705_),
    .B1(_1576_),
    .B2(_1585_),
    .ZN(_1724_));
 NAND2_X1 _4079_ (.A1(_1631_),
    .A2(\last_valid_data[7] ),
    .ZN(_1725_));
 OAI21_X1 _4080_ (.A(_1724_),
    .B1(_1725_),
    .B2(_0910_),
    .ZN(net58));
 OAI22_X1 _4081_ (.A1(_0597_),
    .A2(_0942_),
    .B1(_1597_),
    .B2(_1606_),
    .ZN(_1726_));
 NAND2_X1 _4082_ (.A1(_1631_),
    .A2(\last_valid_data[8] ),
    .ZN(_1727_));
 OAI21_X1 _4083_ (.A(_1726_),
    .B1(_1727_),
    .B2(_0910_),
    .ZN(net59));
 OAI22_X1 _4084_ (.A1(_0597_),
    .A2(_0942_),
    .B1(_1618_),
    .B2(_1627_),
    .ZN(_1728_));
 NAND2_X1 _4085_ (.A1(_1631_),
    .A2(\last_valid_data[9] ),
    .ZN(_1729_));
 OAI21_X1 _4086_ (.A(_1728_),
    .B1(_1729_),
    .B2(_0910_),
    .ZN(net60));
 FA_X1 _4087_ (.A(_2299_),
    .B(\wr_ptr[1] ),
    .CI(_2300_),
    .CO(_2301_),
    .S(net5));
 HA_X1 _4088_ (.A(_2302_),
    .B(\wr_ptr[3] ),
    .CO(_2303_),
    .S(_2304_));
 HA_X1 _4089_ (.A(_2299_),
    .B(\wr_ptr[1] ),
    .CO(_2305_),
    .S(_2306_));
 HA_X1 _4090_ (.A(_2307_),
    .B(\wr_ptr[2] ),
    .CO(_2308_),
    .S(_2309_));
 HA_X1 _4091_ (.A(net65),
    .B(\rd_ptr[1] ),
    .CO(_2310_),
    .S(_0007_));
 HA_X1 _4092_ (.A(net10),
    .B(net17),
    .CO(_2311_),
    .S(_0009_));
 HA_X1 _4093_ (.A(_0004_),
    .B(_2312_),
    .CO(_2313_),
    .S(_0005_));
 HA_X1 _4094_ (.A(_0004_),
    .B(\wr_ptr[1] ),
    .CO(_2314_),
    .S(_2315_));
 HA_X1 _4095_ (.A(\wr_ptr[0] ),
    .B(_2312_),
    .CO(_2316_),
    .S(_2317_));
 HA_X1 _4096_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_2318_),
    .S(_2319_));
 HA_X1 _4097_ (.A(\rd_ptr[0] ),
    .B(_0004_),
    .CO(_2320_),
    .S(_2321_));
 DFF_X1 _4098_ (.D(_0010_),
    .CK(clknet_leaf_36_clk),
    .Q(_0000_),
    .QN(_2298_));
 DFF_X1 _4099_ (.D(_0011_),
    .CK(clknet_leaf_36_clk),
    .Q(_0001_),
    .QN(_2297_));
 DFF_X1 _4100_ (.D(_0012_),
    .CK(clknet_leaf_35_clk),
    .Q(_0002_),
    .QN(_2296_));
 DFF_X1 _4101_ (.D(_0013_),
    .CK(clknet_leaf_36_clk),
    .Q(_0003_),
    .QN(_2295_));
 DFF_X2 \error_count[0]$_SDFFE_PN0P_  (.D(_0014_),
    .CK(clknet_leaf_39_clk),
    .Q(net10),
    .QN(_0008_));
 DFF_X1 \error_count[10]$_SDFFE_PN0P_  (.D(_0015_),
    .CK(clknet_leaf_37_clk),
    .Q(net11),
    .QN(_2294_));
 DFF_X1 \error_count[11]$_SDFFE_PN0P_  (.D(_0016_),
    .CK(clknet_leaf_37_clk),
    .Q(net12),
    .QN(_2293_));
 DFF_X1 \error_count[12]$_SDFFE_PN0P_  (.D(_0017_),
    .CK(clknet_leaf_37_clk),
    .Q(net13),
    .QN(_2292_));
 DFF_X1 \error_count[13]$_SDFFE_PN0P_  (.D(_0018_),
    .CK(clknet_leaf_37_clk),
    .Q(net14),
    .QN(_2291_));
 DFF_X1 \error_count[14]$_SDFFE_PN0P_  (.D(_0019_),
    .CK(clknet_leaf_37_clk),
    .Q(net15),
    .QN(_2290_));
 DFF_X1 \error_count[15]$_SDFFE_PN0P_  (.D(_0020_),
    .CK(clknet_leaf_37_clk),
    .Q(net16),
    .QN(_2289_));
 DFF_X2 \error_count[1]$_SDFFE_PN0P_  (.D(_0021_),
    .CK(clknet_leaf_38_clk),
    .Q(net17),
    .QN(_2288_));
 DFF_X1 \error_count[2]$_SDFFE_PN0P_  (.D(_0022_),
    .CK(clknet_leaf_39_clk),
    .Q(net18),
    .QN(_2287_));
 DFF_X1 \error_count[3]$_SDFFE_PN0P_  (.D(_0023_),
    .CK(clknet_leaf_38_clk),
    .Q(net19),
    .QN(_2286_));
 DFF_X1 \error_count[4]$_SDFFE_PN0P_  (.D(_0024_),
    .CK(clknet_leaf_38_clk),
    .Q(net20),
    .QN(_2285_));
 DFF_X1 \error_count[5]$_SDFFE_PN0P_  (.D(_0025_),
    .CK(clknet_leaf_37_clk),
    .Q(net21),
    .QN(_2284_));
 DFF_X1 \error_count[6]$_SDFFE_PN0P_  (.D(_0026_),
    .CK(clknet_leaf_38_clk),
    .Q(net22),
    .QN(_2283_));
 DFF_X2 \error_count[7]$_SDFFE_PN0P_  (.D(_0027_),
    .CK(clknet_leaf_38_clk),
    .Q(net23),
    .QN(_2282_));
 DFF_X1 \error_count[8]$_SDFFE_PN0P_  (.D(_0028_),
    .CK(clknet_leaf_38_clk),
    .Q(net24),
    .QN(_2281_));
 DFF_X1 \error_count[9]$_SDFFE_PN0P_  (.D(_0029_),
    .CK(clknet_leaf_39_clk),
    .Q(net25),
    .QN(_2280_));
 DFF_X1 \error_detected$_SDFF_PN0_  (.D(_0030_),
    .CK(clknet_leaf_38_clk),
    .Q(net26),
    .QN(_2279_));
 DFF_X1 \last_valid_data[0]$_SDFFE_PN0P_  (.D(_0031_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[0] ),
    .QN(_2278_));
 DFF_X1 \last_valid_data[10]$_SDFFE_PN0P_  (.D(_0032_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[10] ),
    .QN(_2277_));
 DFF_X1 \last_valid_data[11]$_SDFFE_PN0P_  (.D(_0033_),
    .CK(clknet_leaf_42_clk),
    .Q(\last_valid_data[11] ),
    .QN(_2276_));
 DFF_X1 \last_valid_data[12]$_SDFFE_PN0P_  (.D(_0034_),
    .CK(clknet_leaf_42_clk),
    .Q(\last_valid_data[12] ),
    .QN(_2275_));
 DFF_X1 \last_valid_data[13]$_SDFFE_PN0P_  (.D(_0035_),
    .CK(clknet_leaf_52_clk),
    .Q(\last_valid_data[13] ),
    .QN(_2274_));
 DFF_X1 \last_valid_data[14]$_SDFFE_PN0P_  (.D(_0036_),
    .CK(clknet_leaf_42_clk),
    .Q(\last_valid_data[14] ),
    .QN(_2273_));
 DFF_X1 \last_valid_data[15]$_SDFFE_PN0P_  (.D(_0037_),
    .CK(clknet_leaf_42_clk),
    .Q(\last_valid_data[15] ),
    .QN(_2272_));
 DFF_X1 \last_valid_data[16]$_SDFFE_PN0P_  (.D(_0038_),
    .CK(clknet_leaf_41_clk),
    .Q(\last_valid_data[16] ),
    .QN(_2271_));
 DFF_X1 \last_valid_data[17]$_SDFFE_PN0P_  (.D(_0039_),
    .CK(clknet_leaf_41_clk),
    .Q(\last_valid_data[17] ),
    .QN(_2270_));
 DFF_X1 \last_valid_data[18]$_SDFFE_PN0P_  (.D(_0040_),
    .CK(clknet_leaf_44_clk),
    .Q(\last_valid_data[18] ),
    .QN(_2269_));
 DFF_X1 \last_valid_data[19]$_SDFFE_PN0P_  (.D(_0041_),
    .CK(clknet_leaf_30_clk),
    .Q(\last_valid_data[19] ),
    .QN(_2268_));
 DFF_X1 \last_valid_data[1]$_SDFFE_PN0P_  (.D(_0042_),
    .CK(clknet_leaf_33_clk),
    .Q(\last_valid_data[1] ),
    .QN(_2267_));
 DFF_X1 \last_valid_data[20]$_SDFFE_PN0P_  (.D(_0043_),
    .CK(clknet_leaf_33_clk),
    .Q(\last_valid_data[20] ),
    .QN(_2266_));
 DFF_X1 \last_valid_data[21]$_SDFFE_PN0P_  (.D(_0044_),
    .CK(clknet_leaf_26_clk),
    .Q(\last_valid_data[21] ),
    .QN(_2265_));
 DFF_X1 \last_valid_data[22]$_SDFFE_PN0P_  (.D(_0045_),
    .CK(clknet_leaf_26_clk),
    .Q(\last_valid_data[22] ),
    .QN(_2264_));
 DFF_X1 \last_valid_data[23]$_SDFFE_PN0P_  (.D(_0046_),
    .CK(clknet_leaf_27_clk),
    .Q(\last_valid_data[23] ),
    .QN(_2263_));
 DFF_X1 \last_valid_data[24]$_SDFFE_PN0P_  (.D(_0047_),
    .CK(clknet_leaf_27_clk),
    .Q(\last_valid_data[24] ),
    .QN(_2262_));
 DFF_X1 \last_valid_data[25]$_SDFFE_PN0P_  (.D(_0048_),
    .CK(clknet_leaf_27_clk),
    .Q(\last_valid_data[25] ),
    .QN(_2261_));
 DFF_X1 \last_valid_data[26]$_SDFFE_PN0P_  (.D(_0049_),
    .CK(clknet_leaf_10_clk),
    .Q(\last_valid_data[26] ),
    .QN(_2260_));
 DFF_X1 \last_valid_data[27]$_SDFFE_PN0P_  (.D(_0050_),
    .CK(clknet_leaf_10_clk),
    .Q(\last_valid_data[27] ),
    .QN(_2259_));
 DFF_X1 \last_valid_data[28]$_SDFFE_PN0P_  (.D(_0051_),
    .CK(clknet_leaf_6_clk),
    .Q(\last_valid_data[28] ),
    .QN(_2258_));
 DFF_X1 \last_valid_data[29]$_SDFFE_PN0P_  (.D(_0052_),
    .CK(clknet_leaf_6_clk),
    .Q(\last_valid_data[29] ),
    .QN(_2257_));
 DFF_X1 \last_valid_data[2]$_SDFFE_PN0P_  (.D(_0053_),
    .CK(clknet_leaf_12_clk),
    .Q(\last_valid_data[2] ),
    .QN(_2256_));
 DFF_X1 \last_valid_data[30]$_SDFFE_PN0P_  (.D(_0054_),
    .CK(clknet_leaf_12_clk),
    .Q(\last_valid_data[30] ),
    .QN(_2255_));
 DFF_X1 \last_valid_data[31]$_SDFFE_PN0P_  (.D(_0055_),
    .CK(clknet_leaf_13_clk),
    .Q(\last_valid_data[31] ),
    .QN(_2254_));
 DFF_X1 \last_valid_data[3]$_SDFFE_PN0P_  (.D(_0056_),
    .CK(clknet_leaf_10_clk),
    .Q(\last_valid_data[3] ),
    .QN(_2253_));
 DFF_X1 \last_valid_data[4]$_SDFFE_PN0P_  (.D(_0057_),
    .CK(clknet_leaf_10_clk),
    .Q(\last_valid_data[4] ),
    .QN(_2252_));
 DFF_X1 \last_valid_data[5]$_SDFFE_PN0P_  (.D(_0058_),
    .CK(clknet_leaf_9_clk),
    .Q(\last_valid_data[5] ),
    .QN(_2251_));
 DFF_X1 \last_valid_data[6]$_SDFFE_PN0P_  (.D(_0059_),
    .CK(clknet_leaf_9_clk),
    .Q(\last_valid_data[6] ),
    .QN(_2250_));
 DFF_X1 \last_valid_data[7]$_SDFFE_PN0P_  (.D(_0060_),
    .CK(clknet_leaf_46_clk),
    .Q(\last_valid_data[7] ),
    .QN(_2249_));
 DFF_X1 \last_valid_data[8]$_SDFFE_PN0P_  (.D(_0061_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[8] ),
    .QN(_2248_));
 DFF_X1 \last_valid_data[9]$_SDFFE_PN0P_  (.D(_0062_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[9] ),
    .QN(_2247_));
 DFF_X1 \last_valid_data_available$_SDFFE_PN0P_  (.D(_0063_),
    .CK(clknet_leaf_39_clk),
    .Q(last_valid_data_available),
    .QN(_2246_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[0][0] ),
    .QN(_2245_));
 DFF_X1 \mem[0][10]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[0][10] ),
    .QN(_2244_));
 DFF_X1 \mem[0][11]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[0][11] ),
    .QN(_2243_));
 DFF_X1 \mem[0][12]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[0][12] ),
    .QN(_2242_));
 DFF_X1 \mem[0][13]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[0][13] ),
    .QN(_2241_));
 DFF_X1 \mem[0][14]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[0][14] ),
    .QN(_2240_));
 DFF_X1 \mem[0][15]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[0][15] ),
    .QN(_2239_));
 DFF_X1 \mem[0][16]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_leaf_41_clk),
    .Q(\mem[0][16] ),
    .QN(_2238_));
 DFF_X1 \mem[0][17]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[0][17] ),
    .QN(_2237_));
 DFF_X1 \mem[0][18]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[0][18] ),
    .QN(_2236_));
 DFF_X1 \mem[0][19]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[0][19] ),
    .QN(_2235_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[0][1] ),
    .QN(_2234_));
 DFF_X1 \mem[0][20]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[0][20] ),
    .QN(_2233_));
 DFF_X1 \mem[0][21]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[0][21] ),
    .QN(_2232_));
 DFF_X1 \mem[0][22]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[0][22] ),
    .QN(_2231_));
 DFF_X1 \mem[0][23]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[0][23] ),
    .QN(_2230_));
 DFF_X1 \mem[0][24]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[0][24] ),
    .QN(_2229_));
 DFF_X1 \mem[0][25]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[0][25] ),
    .QN(_2228_));
 DFF_X1 \mem[0][26]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[0][26] ),
    .QN(_2227_));
 DFF_X1 \mem[0][27]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[0][27] ),
    .QN(_2226_));
 DFF_X1 \mem[0][28]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[0][28] ),
    .QN(_2225_));
 DFF_X1 \mem[0][29]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[0][29] ),
    .QN(_2224_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[0][2] ),
    .QN(_2223_));
 DFF_X1 \mem[0][30]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[0][30] ),
    .QN(_2222_));
 DFF_X1 \mem[0][31]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[0][31] ),
    .QN(_2221_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[0][3] ),
    .QN(_2220_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[0][4] ),
    .QN(_2219_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[0][5] ),
    .QN(_2218_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[0][6] ),
    .QN(_2217_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[0][7] ),
    .QN(_2216_));
 DFF_X1 \mem[0][8]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[0][8] ),
    .QN(_2215_));
 DFF_X1 \mem[0][9]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[0][9] ),
    .QN(_2214_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[10][0] ),
    .QN(_2213_));
 DFF_X1 \mem[10][10]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[10][10] ),
    .QN(_2212_));
 DFF_X1 \mem[10][11]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[10][11] ),
    .QN(_2211_));
 DFF_X1 \mem[10][12]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[10][12] ),
    .QN(_2210_));
 DFF_X1 \mem[10][13]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[10][13] ),
    .QN(_2209_));
 DFF_X1 \mem[10][14]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[10][14] ),
    .QN(_2208_));
 DFF_X1 \mem[10][15]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[10][15] ),
    .QN(_2207_));
 DFF_X1 \mem[10][16]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[10][16] ),
    .QN(_2206_));
 DFF_X1 \mem[10][17]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[10][17] ),
    .QN(_2205_));
 DFF_X1 \mem[10][18]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[10][18] ),
    .QN(_2204_));
 DFF_X1 \mem[10][19]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[10][19] ),
    .QN(_2203_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[10][1] ),
    .QN(_2202_));
 DFF_X1 \mem[10][20]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[10][20] ),
    .QN(_2201_));
 DFF_X1 \mem[10][21]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[10][21] ),
    .QN(_2200_));
 DFF_X1 \mem[10][22]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[10][22] ),
    .QN(_2199_));
 DFF_X1 \mem[10][23]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[10][23] ),
    .QN(_2198_));
 DFF_X1 \mem[10][24]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[10][24] ),
    .QN(_2197_));
 DFF_X1 \mem[10][25]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[10][25] ),
    .QN(_2196_));
 DFF_X1 \mem[10][26]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[10][26] ),
    .QN(_2195_));
 DFF_X1 \mem[10][27]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[10][27] ),
    .QN(_2194_));
 DFF_X1 \mem[10][28]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[10][28] ),
    .QN(_2193_));
 DFF_X1 \mem[10][29]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[10][29] ),
    .QN(_2192_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[10][2] ),
    .QN(_2191_));
 DFF_X1 \mem[10][30]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[10][30] ),
    .QN(_2190_));
 DFF_X1 \mem[10][31]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[10][31] ),
    .QN(_2189_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[10][3] ),
    .QN(_2188_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[10][4] ),
    .QN(_2187_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[10][5] ),
    .QN(_2186_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[10][6] ),
    .QN(_2185_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[10][7] ),
    .QN(_2184_));
 DFF_X1 \mem[10][8]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[10][8] ),
    .QN(_2183_));
 DFF_X1 \mem[10][9]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[10][9] ),
    .QN(_2182_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[11][0] ),
    .QN(_2181_));
 DFF_X1 \mem[11][10]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[11][10] ),
    .QN(_2180_));
 DFF_X1 \mem[11][11]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[11][11] ),
    .QN(_2179_));
 DFF_X1 \mem[11][12]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[11][12] ),
    .QN(_2178_));
 DFF_X1 \mem[11][13]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[11][13] ),
    .QN(_2177_));
 DFF_X1 \mem[11][14]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[11][14] ),
    .QN(_2176_));
 DFF_X1 \mem[11][15]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[11][15] ),
    .QN(_2175_));
 DFF_X1 \mem[11][16]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[11][16] ),
    .QN(_2174_));
 DFF_X1 \mem[11][17]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[11][17] ),
    .QN(_2173_));
 DFF_X1 \mem[11][18]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[11][18] ),
    .QN(_2172_));
 DFF_X1 \mem[11][19]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[11][19] ),
    .QN(_2171_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[11][1] ),
    .QN(_2170_));
 DFF_X1 \mem[11][20]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[11][20] ),
    .QN(_2169_));
 DFF_X1 \mem[11][21]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[11][21] ),
    .QN(_2168_));
 DFF_X1 \mem[11][22]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[11][22] ),
    .QN(_2167_));
 DFF_X1 \mem[11][23]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[11][23] ),
    .QN(_2166_));
 DFF_X1 \mem[11][24]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[11][24] ),
    .QN(_2165_));
 DFF_X1 \mem[11][25]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[11][25] ),
    .QN(_2164_));
 DFF_X1 \mem[11][26]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[11][26] ),
    .QN(_2163_));
 DFF_X1 \mem[11][27]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[11][27] ),
    .QN(_2162_));
 DFF_X1 \mem[11][28]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[11][28] ),
    .QN(_2161_));
 DFF_X1 \mem[11][29]$_DFFE_PP_  (.D(_0149_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[11][29] ),
    .QN(_2160_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0150_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[11][2] ),
    .QN(_2159_));
 DFF_X1 \mem[11][30]$_DFFE_PP_  (.D(_0151_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[11][30] ),
    .QN(_2158_));
 DFF_X1 \mem[11][31]$_DFFE_PP_  (.D(_0152_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[11][31] ),
    .QN(_2157_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0153_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[11][3] ),
    .QN(_2156_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0154_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[11][4] ),
    .QN(_2155_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0155_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[11][5] ),
    .QN(_2154_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0156_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[11][6] ),
    .QN(_2153_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0157_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[11][7] ),
    .QN(_2152_));
 DFF_X1 \mem[11][8]$_DFFE_PP_  (.D(_0158_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[11][8] ),
    .QN(_2151_));
 DFF_X1 \mem[11][9]$_DFFE_PP_  (.D(_0159_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[11][9] ),
    .QN(_2150_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0160_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[12][0] ),
    .QN(_2149_));
 DFF_X1 \mem[12][10]$_DFFE_PP_  (.D(_0161_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[12][10] ),
    .QN(_2148_));
 DFF_X1 \mem[12][11]$_DFFE_PP_  (.D(_0162_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[12][11] ),
    .QN(_2147_));
 DFF_X1 \mem[12][12]$_DFFE_PP_  (.D(_0163_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[12][12] ),
    .QN(_2146_));
 DFF_X1 \mem[12][13]$_DFFE_PP_  (.D(_0164_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[12][13] ),
    .QN(_2145_));
 DFF_X1 \mem[12][14]$_DFFE_PP_  (.D(_0165_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[12][14] ),
    .QN(_2144_));
 DFF_X1 \mem[12][15]$_DFFE_PP_  (.D(_0166_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[12][15] ),
    .QN(_2143_));
 DFF_X1 \mem[12][16]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[12][16] ),
    .QN(_2142_));
 DFF_X1 \mem[12][17]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[12][17] ),
    .QN(_2141_));
 DFF_X1 \mem[12][18]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[12][18] ),
    .QN(_2140_));
 DFF_X1 \mem[12][19]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[12][19] ),
    .QN(_2139_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[12][1] ),
    .QN(_2138_));
 DFF_X1 \mem[12][20]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[12][20] ),
    .QN(_2137_));
 DFF_X1 \mem[12][21]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[12][21] ),
    .QN(_2136_));
 DFF_X1 \mem[12][22]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[12][22] ),
    .QN(_2135_));
 DFF_X1 \mem[12][23]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[12][23] ),
    .QN(_2134_));
 DFF_X1 \mem[12][24]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[12][24] ),
    .QN(_2133_));
 DFF_X1 \mem[12][25]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[12][25] ),
    .QN(_2132_));
 DFF_X1 \mem[12][26]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[12][26] ),
    .QN(_2131_));
 DFF_X1 \mem[12][27]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[12][27] ),
    .QN(_2130_));
 DFF_X1 \mem[12][28]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[12][28] ),
    .QN(_2129_));
 DFF_X1 \mem[12][29]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[12][29] ),
    .QN(_2128_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[12][2] ),
    .QN(_2127_));
 DFF_X1 \mem[12][30]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[12][30] ),
    .QN(_2126_));
 DFF_X1 \mem[12][31]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[12][31] ),
    .QN(_2125_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[12][3] ),
    .QN(_2124_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[12][4] ),
    .QN(_2123_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[12][5] ),
    .QN(_2122_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[12][6] ),
    .QN(_2121_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[12][7] ),
    .QN(_2120_));
 DFF_X1 \mem[12][8]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[12][8] ),
    .QN(_2119_));
 DFF_X1 \mem[12][9]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[12][9] ),
    .QN(_2118_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0192_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[13][0] ),
    .QN(_2117_));
 DFF_X1 \mem[13][10]$_DFFE_PP_  (.D(_0193_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[13][10] ),
    .QN(_2116_));
 DFF_X1 \mem[13][11]$_DFFE_PP_  (.D(_0194_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[13][11] ),
    .QN(_2115_));
 DFF_X1 \mem[13][12]$_DFFE_PP_  (.D(_0195_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[13][12] ),
    .QN(_2114_));
 DFF_X1 \mem[13][13]$_DFFE_PP_  (.D(_0196_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[13][13] ),
    .QN(_2113_));
 DFF_X1 \mem[13][14]$_DFFE_PP_  (.D(_0197_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[13][14] ),
    .QN(_2112_));
 DFF_X1 \mem[13][15]$_DFFE_PP_  (.D(_0198_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[13][15] ),
    .QN(_2111_));
 DFF_X1 \mem[13][16]$_DFFE_PP_  (.D(_0199_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[13][16] ),
    .QN(_2110_));
 DFF_X1 \mem[13][17]$_DFFE_PP_  (.D(_0200_),
    .CK(clknet_leaf_43_clk),
    .Q(\mem[13][17] ),
    .QN(_2109_));
 DFF_X1 \mem[13][18]$_DFFE_PP_  (.D(_0201_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[13][18] ),
    .QN(_2108_));
 DFF_X1 \mem[13][19]$_DFFE_PP_  (.D(_0202_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[13][19] ),
    .QN(_2107_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0203_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[13][1] ),
    .QN(_2106_));
 DFF_X1 \mem[13][20]$_DFFE_PP_  (.D(_0204_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[13][20] ),
    .QN(_2105_));
 DFF_X1 \mem[13][21]$_DFFE_PP_  (.D(_0205_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[13][21] ),
    .QN(_2104_));
 DFF_X1 \mem[13][22]$_DFFE_PP_  (.D(_0206_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[13][22] ),
    .QN(_2103_));
 DFF_X1 \mem[13][23]$_DFFE_PP_  (.D(_0207_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[13][23] ),
    .QN(_2102_));
 DFF_X1 \mem[13][24]$_DFFE_PP_  (.D(_0208_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[13][24] ),
    .QN(_2101_));
 DFF_X1 \mem[13][25]$_DFFE_PP_  (.D(_0209_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[13][25] ),
    .QN(_2100_));
 DFF_X1 \mem[13][26]$_DFFE_PP_  (.D(_0210_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[13][26] ),
    .QN(_2099_));
 DFF_X1 \mem[13][27]$_DFFE_PP_  (.D(_0211_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[13][27] ),
    .QN(_2098_));
 DFF_X1 \mem[13][28]$_DFFE_PP_  (.D(_0212_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[13][28] ),
    .QN(_2097_));
 DFF_X1 \mem[13][29]$_DFFE_PP_  (.D(_0213_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[13][29] ),
    .QN(_2096_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0214_),
    .CK(clknet_leaf_79_clk),
    .Q(\mem[13][2] ),
    .QN(_2095_));
 DFF_X1 \mem[13][30]$_DFFE_PP_  (.D(_0215_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[13][30] ),
    .QN(_2094_));
 DFF_X1 \mem[13][31]$_DFFE_PP_  (.D(_0216_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[13][31] ),
    .QN(_2093_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0217_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[13][3] ),
    .QN(_2092_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0218_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[13][4] ),
    .QN(_2091_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0219_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[13][5] ),
    .QN(_2090_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0220_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[13][6] ),
    .QN(_2089_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0221_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[13][7] ),
    .QN(_2088_));
 DFF_X1 \mem[13][8]$_DFFE_PP_  (.D(_0222_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[13][8] ),
    .QN(_2087_));
 DFF_X1 \mem[13][9]$_DFFE_PP_  (.D(_0223_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[13][9] ),
    .QN(_2086_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0224_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[14][0] ),
    .QN(_2085_));
 DFF_X1 \mem[14][10]$_DFFE_PP_  (.D(_0225_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[14][10] ),
    .QN(_2084_));
 DFF_X1 \mem[14][11]$_DFFE_PP_  (.D(_0226_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[14][11] ),
    .QN(_2083_));
 DFF_X1 \mem[14][12]$_DFFE_PP_  (.D(_0227_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[14][12] ),
    .QN(_2082_));
 DFF_X1 \mem[14][13]$_DFFE_PP_  (.D(_0228_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[14][13] ),
    .QN(_2081_));
 DFF_X1 \mem[14][14]$_DFFE_PP_  (.D(_0229_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[14][14] ),
    .QN(_2080_));
 DFF_X1 \mem[14][15]$_DFFE_PP_  (.D(_0230_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[14][15] ),
    .QN(_2079_));
 DFF_X1 \mem[14][16]$_DFFE_PP_  (.D(_0231_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[14][16] ),
    .QN(_2078_));
 DFF_X1 \mem[14][17]$_DFFE_PP_  (.D(_0232_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[14][17] ),
    .QN(_2077_));
 DFF_X1 \mem[14][18]$_DFFE_PP_  (.D(_0233_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[14][18] ),
    .QN(_2076_));
 DFF_X1 \mem[14][19]$_DFFE_PP_  (.D(_0234_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[14][19] ),
    .QN(_2075_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0235_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[14][1] ),
    .QN(_2074_));
 DFF_X1 \mem[14][20]$_DFFE_PP_  (.D(_0236_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[14][20] ),
    .QN(_2073_));
 DFF_X1 \mem[14][21]$_DFFE_PP_  (.D(_0237_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[14][21] ),
    .QN(_2072_));
 DFF_X1 \mem[14][22]$_DFFE_PP_  (.D(_0238_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[14][22] ),
    .QN(_2071_));
 DFF_X1 \mem[14][23]$_DFFE_PP_  (.D(_0239_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[14][23] ),
    .QN(_2070_));
 DFF_X1 \mem[14][24]$_DFFE_PP_  (.D(_0240_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[14][24] ),
    .QN(_2069_));
 DFF_X1 \mem[14][25]$_DFFE_PP_  (.D(_0241_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[14][25] ),
    .QN(_2068_));
 DFF_X1 \mem[14][26]$_DFFE_PP_  (.D(_0242_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[14][26] ),
    .QN(_2067_));
 DFF_X1 \mem[14][27]$_DFFE_PP_  (.D(_0243_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[14][27] ),
    .QN(_2066_));
 DFF_X1 \mem[14][28]$_DFFE_PP_  (.D(_0244_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[14][28] ),
    .QN(_2065_));
 DFF_X1 \mem[14][29]$_DFFE_PP_  (.D(_0245_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[14][29] ),
    .QN(_2064_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0246_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[14][2] ),
    .QN(_2063_));
 DFF_X1 \mem[14][30]$_DFFE_PP_  (.D(_0247_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[14][30] ),
    .QN(_2062_));
 DFF_X1 \mem[14][31]$_DFFE_PP_  (.D(_0248_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[14][31] ),
    .QN(_2061_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0249_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[14][3] ),
    .QN(_2060_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0250_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[14][4] ),
    .QN(_2059_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0251_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[14][5] ),
    .QN(_2058_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0252_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[14][6] ),
    .QN(_2057_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0253_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[14][7] ),
    .QN(_2056_));
 DFF_X1 \mem[14][8]$_DFFE_PP_  (.D(_0254_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[14][8] ),
    .QN(_2055_));
 DFF_X1 \mem[14][9]$_DFFE_PP_  (.D(_0255_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[14][9] ),
    .QN(_2054_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0256_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[15][0] ),
    .QN(_2053_));
 DFF_X1 \mem[15][10]$_DFFE_PP_  (.D(_0257_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[15][10] ),
    .QN(_2052_));
 DFF_X1 \mem[15][11]$_DFFE_PP_  (.D(_0258_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[15][11] ),
    .QN(_2051_));
 DFF_X1 \mem[15][12]$_DFFE_PP_  (.D(_0259_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[15][12] ),
    .QN(_2050_));
 DFF_X1 \mem[15][13]$_DFFE_PP_  (.D(_0260_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[15][13] ),
    .QN(_2049_));
 DFF_X1 \mem[15][14]$_DFFE_PP_  (.D(_0261_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[15][14] ),
    .QN(_2048_));
 DFF_X1 \mem[15][15]$_DFFE_PP_  (.D(_0262_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[15][15] ),
    .QN(_2047_));
 DFF_X1 \mem[15][16]$_DFFE_PP_  (.D(_0263_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[15][16] ),
    .QN(_2046_));
 DFF_X1 \mem[15][17]$_DFFE_PP_  (.D(_0264_),
    .CK(clknet_leaf_41_clk),
    .Q(\mem[15][17] ),
    .QN(_2045_));
 DFF_X1 \mem[15][18]$_DFFE_PP_  (.D(_0265_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[15][18] ),
    .QN(_2044_));
 DFF_X1 \mem[15][19]$_DFFE_PP_  (.D(_0266_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[15][19] ),
    .QN(_2043_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0267_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[15][1] ),
    .QN(_2042_));
 DFF_X1 \mem[15][20]$_DFFE_PP_  (.D(_0268_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[15][20] ),
    .QN(_2041_));
 DFF_X1 \mem[15][21]$_DFFE_PP_  (.D(_0269_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[15][21] ),
    .QN(_2040_));
 DFF_X1 \mem[15][22]$_DFFE_PP_  (.D(_0270_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[15][22] ),
    .QN(_2039_));
 DFF_X1 \mem[15][23]$_DFFE_PP_  (.D(_0271_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[15][23] ),
    .QN(_2038_));
 DFF_X1 \mem[15][24]$_DFFE_PP_  (.D(_0272_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[15][24] ),
    .QN(_2037_));
 DFF_X1 \mem[15][25]$_DFFE_PP_  (.D(_0273_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[15][25] ),
    .QN(_2036_));
 DFF_X1 \mem[15][26]$_DFFE_PP_  (.D(_0274_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[15][26] ),
    .QN(_2035_));
 DFF_X1 \mem[15][27]$_DFFE_PP_  (.D(_0275_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[15][27] ),
    .QN(_2034_));
 DFF_X1 \mem[15][28]$_DFFE_PP_  (.D(_0276_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[15][28] ),
    .QN(_2033_));
 DFF_X1 \mem[15][29]$_DFFE_PP_  (.D(_0277_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[15][29] ),
    .QN(_2032_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0278_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[15][2] ),
    .QN(_2031_));
 DFF_X1 \mem[15][30]$_DFFE_PP_  (.D(_0279_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[15][30] ),
    .QN(_2030_));
 DFF_X1 \mem[15][31]$_DFFE_PP_  (.D(_0280_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[15][31] ),
    .QN(_2029_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0281_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[15][3] ),
    .QN(_2028_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0282_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[15][4] ),
    .QN(_2027_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0283_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[15][5] ),
    .QN(_2026_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0284_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[15][6] ),
    .QN(_2025_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0285_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[15][7] ),
    .QN(_2024_));
 DFF_X1 \mem[15][8]$_DFFE_PP_  (.D(_0286_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[15][8] ),
    .QN(_2023_));
 DFF_X1 \mem[15][9]$_DFFE_PP_  (.D(_0287_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[15][9] ),
    .QN(_2022_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0288_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[1][0] ),
    .QN(_2021_));
 DFF_X1 \mem[1][10]$_DFFE_PP_  (.D(_0289_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[1][10] ),
    .QN(_2020_));
 DFF_X1 \mem[1][11]$_DFFE_PP_  (.D(_0290_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[1][11] ),
    .QN(_2019_));
 DFF_X1 \mem[1][12]$_DFFE_PP_  (.D(_0291_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[1][12] ),
    .QN(_2018_));
 DFF_X1 \mem[1][13]$_DFFE_PP_  (.D(_0292_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[1][13] ),
    .QN(_2017_));
 DFF_X1 \mem[1][14]$_DFFE_PP_  (.D(_0293_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[1][14] ),
    .QN(_2016_));
 DFF_X1 \mem[1][15]$_DFFE_PP_  (.D(_0294_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[1][15] ),
    .QN(_2015_));
 DFF_X1 \mem[1][16]$_DFFE_PP_  (.D(_0295_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[1][16] ),
    .QN(_2014_));
 DFF_X1 \mem[1][17]$_DFFE_PP_  (.D(_0296_),
    .CK(clknet_leaf_41_clk),
    .Q(\mem[1][17] ),
    .QN(_2013_));
 DFF_X1 \mem[1][18]$_DFFE_PP_  (.D(_0297_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[1][18] ),
    .QN(_2012_));
 DFF_X1 \mem[1][19]$_DFFE_PP_  (.D(_0298_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[1][19] ),
    .QN(_2011_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0299_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[1][1] ),
    .QN(_2010_));
 DFF_X1 \mem[1][20]$_DFFE_PP_  (.D(_0300_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[1][20] ),
    .QN(_2009_));
 DFF_X1 \mem[1][21]$_DFFE_PP_  (.D(_0301_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[1][21] ),
    .QN(_2008_));
 DFF_X1 \mem[1][22]$_DFFE_PP_  (.D(_0302_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[1][22] ),
    .QN(_2007_));
 DFF_X1 \mem[1][23]$_DFFE_PP_  (.D(_0303_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[1][23] ),
    .QN(_2006_));
 DFF_X1 \mem[1][24]$_DFFE_PP_  (.D(_0304_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[1][24] ),
    .QN(_2005_));
 DFF_X1 \mem[1][25]$_DFFE_PP_  (.D(_0305_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[1][25] ),
    .QN(_2004_));
 DFF_X1 \mem[1][26]$_DFFE_PP_  (.D(_0306_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[1][26] ),
    .QN(_2003_));
 DFF_X1 \mem[1][27]$_DFFE_PP_  (.D(_0307_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[1][27] ),
    .QN(_2002_));
 DFF_X1 \mem[1][28]$_DFFE_PP_  (.D(_0308_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[1][28] ),
    .QN(_2001_));
 DFF_X1 \mem[1][29]$_DFFE_PP_  (.D(_0309_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[1][29] ),
    .QN(_2000_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0310_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[1][2] ),
    .QN(_1999_));
 DFF_X1 \mem[1][30]$_DFFE_PP_  (.D(_0311_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[1][30] ),
    .QN(_1998_));
 DFF_X1 \mem[1][31]$_DFFE_PP_  (.D(_0312_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[1][31] ),
    .QN(_1997_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0313_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[1][3] ),
    .QN(_1996_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0314_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[1][4] ),
    .QN(_1995_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0315_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[1][5] ),
    .QN(_1994_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0316_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[1][6] ),
    .QN(_1993_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0317_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[1][7] ),
    .QN(_1992_));
 DFF_X1 \mem[1][8]$_DFFE_PP_  (.D(_0318_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[1][8] ),
    .QN(_1991_));
 DFF_X1 \mem[1][9]$_DFFE_PP_  (.D(_0319_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[1][9] ),
    .QN(_1990_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0320_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[2][0] ),
    .QN(_1989_));
 DFF_X1 \mem[2][10]$_DFFE_PP_  (.D(_0321_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[2][10] ),
    .QN(_1988_));
 DFF_X1 \mem[2][11]$_DFFE_PP_  (.D(_0322_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[2][11] ),
    .QN(_1987_));
 DFF_X1 \mem[2][12]$_DFFE_PP_  (.D(_0323_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[2][12] ),
    .QN(_1986_));
 DFF_X1 \mem[2][13]$_DFFE_PP_  (.D(_0324_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[2][13] ),
    .QN(_1985_));
 DFF_X1 \mem[2][14]$_DFFE_PP_  (.D(_0325_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[2][14] ),
    .QN(_1984_));
 DFF_X1 \mem[2][15]$_DFFE_PP_  (.D(_0326_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[2][15] ),
    .QN(_1983_));
 DFF_X1 \mem[2][16]$_DFFE_PP_  (.D(_0327_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[2][16] ),
    .QN(_1982_));
 DFF_X1 \mem[2][17]$_DFFE_PP_  (.D(_0328_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[2][17] ),
    .QN(_1981_));
 DFF_X1 \mem[2][18]$_DFFE_PP_  (.D(_0329_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[2][18] ),
    .QN(_1980_));
 DFF_X1 \mem[2][19]$_DFFE_PP_  (.D(_0330_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[2][19] ),
    .QN(_1979_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0331_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[2][1] ),
    .QN(_1978_));
 DFF_X1 \mem[2][20]$_DFFE_PP_  (.D(_0332_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[2][20] ),
    .QN(_1977_));
 DFF_X1 \mem[2][21]$_DFFE_PP_  (.D(_0333_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[2][21] ),
    .QN(_1976_));
 DFF_X1 \mem[2][22]$_DFFE_PP_  (.D(_0334_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[2][22] ),
    .QN(_1975_));
 DFF_X1 \mem[2][23]$_DFFE_PP_  (.D(_0335_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[2][23] ),
    .QN(_1974_));
 DFF_X1 \mem[2][24]$_DFFE_PP_  (.D(_0336_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[2][24] ),
    .QN(_1973_));
 DFF_X1 \mem[2][25]$_DFFE_PP_  (.D(_0337_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[2][25] ),
    .QN(_1972_));
 DFF_X1 \mem[2][26]$_DFFE_PP_  (.D(_0338_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[2][26] ),
    .QN(_1971_));
 DFF_X1 \mem[2][27]$_DFFE_PP_  (.D(_0339_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[2][27] ),
    .QN(_1970_));
 DFF_X1 \mem[2][28]$_DFFE_PP_  (.D(_0340_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[2][28] ),
    .QN(_1969_));
 DFF_X1 \mem[2][29]$_DFFE_PP_  (.D(_0341_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[2][29] ),
    .QN(_1968_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0342_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[2][2] ),
    .QN(_1967_));
 DFF_X1 \mem[2][30]$_DFFE_PP_  (.D(_0343_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[2][30] ),
    .QN(_1966_));
 DFF_X1 \mem[2][31]$_DFFE_PP_  (.D(_0344_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[2][31] ),
    .QN(_1965_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0345_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[2][3] ),
    .QN(_1964_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0346_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[2][4] ),
    .QN(_1963_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0347_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[2][5] ),
    .QN(_1962_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0348_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[2][6] ),
    .QN(_1961_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0349_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[2][7] ),
    .QN(_1960_));
 DFF_X1 \mem[2][8]$_DFFE_PP_  (.D(_0350_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[2][8] ),
    .QN(_1959_));
 DFF_X1 \mem[2][9]$_DFFE_PP_  (.D(_0351_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[2][9] ),
    .QN(_1958_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0352_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[3][0] ),
    .QN(_1957_));
 DFF_X1 \mem[3][10]$_DFFE_PP_  (.D(_0353_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[3][10] ),
    .QN(_1956_));
 DFF_X1 \mem[3][11]$_DFFE_PP_  (.D(_0354_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[3][11] ),
    .QN(_1955_));
 DFF_X1 \mem[3][12]$_DFFE_PP_  (.D(_0355_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[3][12] ),
    .QN(_1954_));
 DFF_X1 \mem[3][13]$_DFFE_PP_  (.D(_0356_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[3][13] ),
    .QN(_1953_));
 DFF_X1 \mem[3][14]$_DFFE_PP_  (.D(_0357_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[3][14] ),
    .QN(_1952_));
 DFF_X1 \mem[3][15]$_DFFE_PP_  (.D(_0358_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[3][15] ),
    .QN(_1951_));
 DFF_X1 \mem[3][16]$_DFFE_PP_  (.D(_0359_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[3][16] ),
    .QN(_1950_));
 DFF_X1 \mem[3][17]$_DFFE_PP_  (.D(_0360_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[3][17] ),
    .QN(_1949_));
 DFF_X1 \mem[3][18]$_DFFE_PP_  (.D(_0361_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[3][18] ),
    .QN(_1948_));
 DFF_X1 \mem[3][19]$_DFFE_PP_  (.D(_0362_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[3][19] ),
    .QN(_1947_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0363_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[3][1] ),
    .QN(_1946_));
 DFF_X1 \mem[3][20]$_DFFE_PP_  (.D(_0364_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[3][20] ),
    .QN(_1945_));
 DFF_X1 \mem[3][21]$_DFFE_PP_  (.D(_0365_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[3][21] ),
    .QN(_1944_));
 DFF_X1 \mem[3][22]$_DFFE_PP_  (.D(_0366_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[3][22] ),
    .QN(_1943_));
 DFF_X1 \mem[3][23]$_DFFE_PP_  (.D(_0367_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[3][23] ),
    .QN(_1942_));
 DFF_X1 \mem[3][24]$_DFFE_PP_  (.D(_0368_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[3][24] ),
    .QN(_1941_));
 DFF_X1 \mem[3][25]$_DFFE_PP_  (.D(_0369_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[3][25] ),
    .QN(_1940_));
 DFF_X1 \mem[3][26]$_DFFE_PP_  (.D(_0370_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[3][26] ),
    .QN(_1939_));
 DFF_X1 \mem[3][27]$_DFFE_PP_  (.D(_0371_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[3][27] ),
    .QN(_1938_));
 DFF_X1 \mem[3][28]$_DFFE_PP_  (.D(_0372_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[3][28] ),
    .QN(_1937_));
 DFF_X1 \mem[3][29]$_DFFE_PP_  (.D(_0373_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[3][29] ),
    .QN(_1936_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0374_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[3][2] ),
    .QN(_1935_));
 DFF_X1 \mem[3][30]$_DFFE_PP_  (.D(_0375_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[3][30] ),
    .QN(_1934_));
 DFF_X1 \mem[3][31]$_DFFE_PP_  (.D(_0376_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[3][31] ),
    .QN(_1933_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0377_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[3][3] ),
    .QN(_1932_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0378_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[3][4] ),
    .QN(_1931_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0379_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[3][5] ),
    .QN(_1930_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0380_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[3][6] ),
    .QN(_1929_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0381_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[3][7] ),
    .QN(_1928_));
 DFF_X1 \mem[3][8]$_DFFE_PP_  (.D(_0382_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[3][8] ),
    .QN(_1927_));
 DFF_X1 \mem[3][9]$_DFFE_PP_  (.D(_0383_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[3][9] ),
    .QN(_1926_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0384_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[4][0] ),
    .QN(_1925_));
 DFF_X1 \mem[4][10]$_DFFE_PP_  (.D(_0385_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[4][10] ),
    .QN(_1924_));
 DFF_X1 \mem[4][11]$_DFFE_PP_  (.D(_0386_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[4][11] ),
    .QN(_1923_));
 DFF_X1 \mem[4][12]$_DFFE_PP_  (.D(_0387_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[4][12] ),
    .QN(_1922_));
 DFF_X1 \mem[4][13]$_DFFE_PP_  (.D(_0388_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[4][13] ),
    .QN(_1921_));
 DFF_X1 \mem[4][14]$_DFFE_PP_  (.D(_0389_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[4][14] ),
    .QN(_1920_));
 DFF_X1 \mem[4][15]$_DFFE_PP_  (.D(_0390_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[4][15] ),
    .QN(_1919_));
 DFF_X1 \mem[4][16]$_DFFE_PP_  (.D(_0391_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[4][16] ),
    .QN(_1918_));
 DFF_X1 \mem[4][17]$_DFFE_PP_  (.D(_0392_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[4][17] ),
    .QN(_1917_));
 DFF_X1 \mem[4][18]$_DFFE_PP_  (.D(_0393_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[4][18] ),
    .QN(_1916_));
 DFF_X1 \mem[4][19]$_DFFE_PP_  (.D(_0394_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[4][19] ),
    .QN(_1915_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0395_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[4][1] ),
    .QN(_1914_));
 DFF_X1 \mem[4][20]$_DFFE_PP_  (.D(_0396_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[4][20] ),
    .QN(_1913_));
 DFF_X1 \mem[4][21]$_DFFE_PP_  (.D(_0397_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[4][21] ),
    .QN(_1912_));
 DFF_X1 \mem[4][22]$_DFFE_PP_  (.D(_0398_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[4][22] ),
    .QN(_1911_));
 DFF_X1 \mem[4][23]$_DFFE_PP_  (.D(_0399_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[4][23] ),
    .QN(_1910_));
 DFF_X1 \mem[4][24]$_DFFE_PP_  (.D(_0400_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[4][24] ),
    .QN(_1909_));
 DFF_X1 \mem[4][25]$_DFFE_PP_  (.D(_0401_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[4][25] ),
    .QN(_1908_));
 DFF_X1 \mem[4][26]$_DFFE_PP_  (.D(_0402_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[4][26] ),
    .QN(_1907_));
 DFF_X1 \mem[4][27]$_DFFE_PP_  (.D(_0403_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[4][27] ),
    .QN(_1906_));
 DFF_X1 \mem[4][28]$_DFFE_PP_  (.D(_0404_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[4][28] ),
    .QN(_1905_));
 DFF_X1 \mem[4][29]$_DFFE_PP_  (.D(_0405_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[4][29] ),
    .QN(_1904_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0406_),
    .CK(clknet_leaf_79_clk),
    .Q(\mem[4][2] ),
    .QN(_1903_));
 DFF_X1 \mem[4][30]$_DFFE_PP_  (.D(_0407_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[4][30] ),
    .QN(_1902_));
 DFF_X1 \mem[4][31]$_DFFE_PP_  (.D(_0408_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[4][31] ),
    .QN(_1901_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0409_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[4][3] ),
    .QN(_1900_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0410_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[4][4] ),
    .QN(_1899_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0411_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[4][5] ),
    .QN(_1898_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0412_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[4][6] ),
    .QN(_1897_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0413_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[4][7] ),
    .QN(_1896_));
 DFF_X1 \mem[4][8]$_DFFE_PP_  (.D(_0414_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[4][8] ),
    .QN(_1895_));
 DFF_X1 \mem[4][9]$_DFFE_PP_  (.D(_0415_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[4][9] ),
    .QN(_1894_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0416_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[5][0] ),
    .QN(_1893_));
 DFF_X1 \mem[5][10]$_DFFE_PP_  (.D(_0417_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[5][10] ),
    .QN(_1892_));
 DFF_X1 \mem[5][11]$_DFFE_PP_  (.D(_0418_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[5][11] ),
    .QN(_1891_));
 DFF_X1 \mem[5][12]$_DFFE_PP_  (.D(_0419_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[5][12] ),
    .QN(_1890_));
 DFF_X1 \mem[5][13]$_DFFE_PP_  (.D(_0420_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[5][13] ),
    .QN(_1889_));
 DFF_X1 \mem[5][14]$_DFFE_PP_  (.D(_0421_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[5][14] ),
    .QN(_1888_));
 DFF_X1 \mem[5][15]$_DFFE_PP_  (.D(_0422_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[5][15] ),
    .QN(_1887_));
 DFF_X1 \mem[5][16]$_DFFE_PP_  (.D(_0423_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[5][16] ),
    .QN(_1886_));
 DFF_X1 \mem[5][17]$_DFFE_PP_  (.D(_0424_),
    .CK(clknet_leaf_41_clk),
    .Q(\mem[5][17] ),
    .QN(_1885_));
 DFF_X1 \mem[5][18]$_DFFE_PP_  (.D(_0425_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[5][18] ),
    .QN(_1884_));
 DFF_X1 \mem[5][19]$_DFFE_PP_  (.D(_0426_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[5][19] ),
    .QN(_1883_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0427_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[5][1] ),
    .QN(_1882_));
 DFF_X1 \mem[5][20]$_DFFE_PP_  (.D(_0428_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[5][20] ),
    .QN(_1881_));
 DFF_X1 \mem[5][21]$_DFFE_PP_  (.D(_0429_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[5][21] ),
    .QN(_1880_));
 DFF_X1 \mem[5][22]$_DFFE_PP_  (.D(_0430_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[5][22] ),
    .QN(_1879_));
 DFF_X1 \mem[5][23]$_DFFE_PP_  (.D(_0431_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[5][23] ),
    .QN(_1878_));
 DFF_X1 \mem[5][24]$_DFFE_PP_  (.D(_0432_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[5][24] ),
    .QN(_1877_));
 DFF_X1 \mem[5][25]$_DFFE_PP_  (.D(_0433_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[5][25] ),
    .QN(_1876_));
 DFF_X1 \mem[5][26]$_DFFE_PP_  (.D(_0434_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[5][26] ),
    .QN(_1875_));
 DFF_X1 \mem[5][27]$_DFFE_PP_  (.D(_0435_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[5][27] ),
    .QN(_1874_));
 DFF_X1 \mem[5][28]$_DFFE_PP_  (.D(_0436_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[5][28] ),
    .QN(_1873_));
 DFF_X1 \mem[5][29]$_DFFE_PP_  (.D(_0437_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[5][29] ),
    .QN(_1872_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0438_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[5][2] ),
    .QN(_1871_));
 DFF_X1 \mem[5][30]$_DFFE_PP_  (.D(_0439_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[5][30] ),
    .QN(_1870_));
 DFF_X1 \mem[5][31]$_DFFE_PP_  (.D(_0440_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[5][31] ),
    .QN(_1869_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0441_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[5][3] ),
    .QN(_1868_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0442_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[5][4] ),
    .QN(_1867_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0443_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[5][5] ),
    .QN(_1866_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0444_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[5][6] ),
    .QN(_1865_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0445_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[5][7] ),
    .QN(_1864_));
 DFF_X1 \mem[5][8]$_DFFE_PP_  (.D(_0446_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[5][8] ),
    .QN(_1863_));
 DFF_X1 \mem[5][9]$_DFFE_PP_  (.D(_0447_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[5][9] ),
    .QN(_1862_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0448_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[6][0] ),
    .QN(_1861_));
 DFF_X1 \mem[6][10]$_DFFE_PP_  (.D(_0449_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[6][10] ),
    .QN(_1860_));
 DFF_X1 \mem[6][11]$_DFFE_PP_  (.D(_0450_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[6][11] ),
    .QN(_1859_));
 DFF_X1 \mem[6][12]$_DFFE_PP_  (.D(_0451_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[6][12] ),
    .QN(_1858_));
 DFF_X1 \mem[6][13]$_DFFE_PP_  (.D(_0452_),
    .CK(clknet_leaf_49_clk),
    .Q(\mem[6][13] ),
    .QN(_1857_));
 DFF_X1 \mem[6][14]$_DFFE_PP_  (.D(_0453_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[6][14] ),
    .QN(_1856_));
 DFF_X1 \mem[6][15]$_DFFE_PP_  (.D(_0454_),
    .CK(clknet_leaf_43_clk),
    .Q(\mem[6][15] ),
    .QN(_1855_));
 DFF_X1 \mem[6][16]$_DFFE_PP_  (.D(_0455_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[6][16] ),
    .QN(_1854_));
 DFF_X1 \mem[6][17]$_DFFE_PP_  (.D(_0456_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[6][17] ),
    .QN(_1853_));
 DFF_X1 \mem[6][18]$_DFFE_PP_  (.D(_0457_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[6][18] ),
    .QN(_1852_));
 DFF_X1 \mem[6][19]$_DFFE_PP_  (.D(_0458_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[6][19] ),
    .QN(_1851_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0459_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[6][1] ),
    .QN(_1850_));
 DFF_X1 \mem[6][20]$_DFFE_PP_  (.D(_0460_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[6][20] ),
    .QN(_1849_));
 DFF_X1 \mem[6][21]$_DFFE_PP_  (.D(_0461_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[6][21] ),
    .QN(_1848_));
 DFF_X1 \mem[6][22]$_DFFE_PP_  (.D(_0462_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[6][22] ),
    .QN(_1847_));
 DFF_X1 \mem[6][23]$_DFFE_PP_  (.D(_0463_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[6][23] ),
    .QN(_1846_));
 DFF_X1 \mem[6][24]$_DFFE_PP_  (.D(_0464_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[6][24] ),
    .QN(_1845_));
 DFF_X1 \mem[6][25]$_DFFE_PP_  (.D(_0465_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[6][25] ),
    .QN(_1844_));
 DFF_X1 \mem[6][26]$_DFFE_PP_  (.D(_0466_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[6][26] ),
    .QN(_1843_));
 DFF_X1 \mem[6][27]$_DFFE_PP_  (.D(_0467_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[6][27] ),
    .QN(_1842_));
 DFF_X1 \mem[6][28]$_DFFE_PP_  (.D(_0468_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[6][28] ),
    .QN(_1841_));
 DFF_X1 \mem[6][29]$_DFFE_PP_  (.D(_0469_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[6][29] ),
    .QN(_1840_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0470_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[6][2] ),
    .QN(_1839_));
 DFF_X1 \mem[6][30]$_DFFE_PP_  (.D(_0471_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[6][30] ),
    .QN(_1838_));
 DFF_X1 \mem[6][31]$_DFFE_PP_  (.D(_0472_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[6][31] ),
    .QN(_1837_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0473_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[6][3] ),
    .QN(_1836_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0474_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[6][4] ),
    .QN(_1835_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0475_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[6][5] ),
    .QN(_1834_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0476_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[6][6] ),
    .QN(_1833_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0477_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[6][7] ),
    .QN(_1832_));
 DFF_X1 \mem[6][8]$_DFFE_PP_  (.D(_0478_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[6][8] ),
    .QN(_1831_));
 DFF_X1 \mem[6][9]$_DFFE_PP_  (.D(_0479_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[6][9] ),
    .QN(_1830_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0480_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[7][0] ),
    .QN(_1829_));
 DFF_X1 \mem[7][10]$_DFFE_PP_  (.D(_0481_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[7][10] ),
    .QN(_1828_));
 DFF_X1 \mem[7][11]$_DFFE_PP_  (.D(_0482_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[7][11] ),
    .QN(_1827_));
 DFF_X1 \mem[7][12]$_DFFE_PP_  (.D(_0483_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[7][12] ),
    .QN(_1826_));
 DFF_X1 \mem[7][13]$_DFFE_PP_  (.D(_0484_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[7][13] ),
    .QN(_1825_));
 DFF_X1 \mem[7][14]$_DFFE_PP_  (.D(_0485_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[7][14] ),
    .QN(_1824_));
 DFF_X1 \mem[7][15]$_DFFE_PP_  (.D(_0486_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[7][15] ),
    .QN(_1823_));
 DFF_X1 \mem[7][16]$_DFFE_PP_  (.D(_0487_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[7][16] ),
    .QN(_1822_));
 DFF_X1 \mem[7][17]$_DFFE_PP_  (.D(_0488_),
    .CK(clknet_leaf_40_clk),
    .Q(\mem[7][17] ),
    .QN(_1821_));
 DFF_X1 \mem[7][18]$_DFFE_PP_  (.D(_0489_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[7][18] ),
    .QN(_1820_));
 DFF_X1 \mem[7][19]$_DFFE_PP_  (.D(_0490_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[7][19] ),
    .QN(_1819_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0491_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[7][1] ),
    .QN(_1818_));
 DFF_X1 \mem[7][20]$_DFFE_PP_  (.D(_0492_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[7][20] ),
    .QN(_1817_));
 DFF_X1 \mem[7][21]$_DFFE_PP_  (.D(_0493_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[7][21] ),
    .QN(_1816_));
 DFF_X1 \mem[7][22]$_DFFE_PP_  (.D(_0494_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[7][22] ),
    .QN(_1815_));
 DFF_X1 \mem[7][23]$_DFFE_PP_  (.D(_0495_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[7][23] ),
    .QN(_1814_));
 DFF_X1 \mem[7][24]$_DFFE_PP_  (.D(_0496_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[7][24] ),
    .QN(_1813_));
 DFF_X1 \mem[7][25]$_DFFE_PP_  (.D(_0497_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[7][25] ),
    .QN(_1812_));
 DFF_X1 \mem[7][26]$_DFFE_PP_  (.D(_0498_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[7][26] ),
    .QN(_1811_));
 DFF_X1 \mem[7][27]$_DFFE_PP_  (.D(_0499_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[7][27] ),
    .QN(_1810_));
 DFF_X1 \mem[7][28]$_DFFE_PP_  (.D(_0500_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[7][28] ),
    .QN(_1809_));
 DFF_X1 \mem[7][29]$_DFFE_PP_  (.D(_0501_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[7][29] ),
    .QN(_1808_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0502_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[7][2] ),
    .QN(_1807_));
 DFF_X1 \mem[7][30]$_DFFE_PP_  (.D(_0503_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[7][30] ),
    .QN(_1806_));
 DFF_X1 \mem[7][31]$_DFFE_PP_  (.D(_0504_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[7][31] ),
    .QN(_1805_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0505_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[7][3] ),
    .QN(_1804_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0506_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[7][4] ),
    .QN(_1803_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0507_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[7][5] ),
    .QN(_1802_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0508_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[7][6] ),
    .QN(_1801_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0509_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[7][7] ),
    .QN(_1800_));
 DFF_X1 \mem[7][8]$_DFFE_PP_  (.D(_0510_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[7][8] ),
    .QN(_1799_));
 DFF_X1 \mem[7][9]$_DFFE_PP_  (.D(_0511_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[7][9] ),
    .QN(_1798_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0512_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[8][0] ),
    .QN(_1797_));
 DFF_X1 \mem[8][10]$_DFFE_PP_  (.D(_0513_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[8][10] ),
    .QN(_1796_));
 DFF_X1 \mem[8][11]$_DFFE_PP_  (.D(_0514_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[8][11] ),
    .QN(_1795_));
 DFF_X1 \mem[8][12]$_DFFE_PP_  (.D(_0515_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[8][12] ),
    .QN(_1794_));
 DFF_X1 \mem[8][13]$_DFFE_PP_  (.D(_0516_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[8][13] ),
    .QN(_1793_));
 DFF_X1 \mem[8][14]$_DFFE_PP_  (.D(_0517_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[8][14] ),
    .QN(_1792_));
 DFF_X1 \mem[8][15]$_DFFE_PP_  (.D(_0518_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[8][15] ),
    .QN(_1791_));
 DFF_X1 \mem[8][16]$_DFFE_PP_  (.D(_0519_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[8][16] ),
    .QN(_1790_));
 DFF_X1 \mem[8][17]$_DFFE_PP_  (.D(_0520_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[8][17] ),
    .QN(_1789_));
 DFF_X1 \mem[8][18]$_DFFE_PP_  (.D(_0521_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[8][18] ),
    .QN(_1788_));
 DFF_X1 \mem[8][19]$_DFFE_PP_  (.D(_0522_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[8][19] ),
    .QN(_1787_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0523_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[8][1] ),
    .QN(_1786_));
 DFF_X1 \mem[8][20]$_DFFE_PP_  (.D(_0524_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[8][20] ),
    .QN(_1785_));
 DFF_X1 \mem[8][21]$_DFFE_PP_  (.D(_0525_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[8][21] ),
    .QN(_1784_));
 DFF_X1 \mem[8][22]$_DFFE_PP_  (.D(_0526_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[8][22] ),
    .QN(_1783_));
 DFF_X1 \mem[8][23]$_DFFE_PP_  (.D(_0527_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[8][23] ),
    .QN(_1782_));
 DFF_X1 \mem[8][24]$_DFFE_PP_  (.D(_0528_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[8][24] ),
    .QN(_1781_));
 DFF_X1 \mem[8][25]$_DFFE_PP_  (.D(_0529_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[8][25] ),
    .QN(_1780_));
 DFF_X1 \mem[8][26]$_DFFE_PP_  (.D(_0530_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[8][26] ),
    .QN(_1779_));
 DFF_X1 \mem[8][27]$_DFFE_PP_  (.D(_0531_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[8][27] ),
    .QN(_1778_));
 DFF_X1 \mem[8][28]$_DFFE_PP_  (.D(_0532_),
    .CK(clknet_leaf_79_clk),
    .Q(\mem[8][28] ),
    .QN(_1777_));
 DFF_X1 \mem[8][29]$_DFFE_PP_  (.D(_0533_),
    .CK(clknet_leaf_79_clk),
    .Q(\mem[8][29] ),
    .QN(_1776_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0534_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[8][2] ),
    .QN(_1775_));
 DFF_X1 \mem[8][30]$_DFFE_PP_  (.D(_0535_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[8][30] ),
    .QN(_1774_));
 DFF_X1 \mem[8][31]$_DFFE_PP_  (.D(_0536_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[8][31] ),
    .QN(_1773_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0537_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[8][3] ),
    .QN(_1772_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0538_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[8][4] ),
    .QN(_1771_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0539_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[8][5] ),
    .QN(_1770_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0540_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[8][6] ),
    .QN(_1769_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0541_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[8][7] ),
    .QN(_1768_));
 DFF_X1 \mem[8][8]$_DFFE_PP_  (.D(_0542_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[8][8] ),
    .QN(_1767_));
 DFF_X1 \mem[8][9]$_DFFE_PP_  (.D(_0543_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[8][9] ),
    .QN(_1766_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0544_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[9][0] ),
    .QN(_1765_));
 DFF_X1 \mem[9][10]$_DFFE_PP_  (.D(_0545_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[9][10] ),
    .QN(_1764_));
 DFF_X1 \mem[9][11]$_DFFE_PP_  (.D(_0546_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[9][11] ),
    .QN(_1763_));
 DFF_X1 \mem[9][12]$_DFFE_PP_  (.D(_0547_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[9][12] ),
    .QN(_1762_));
 DFF_X1 \mem[9][13]$_DFFE_PP_  (.D(_0548_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[9][13] ),
    .QN(_1761_));
 DFF_X1 \mem[9][14]$_DFFE_PP_  (.D(_0549_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[9][14] ),
    .QN(_1760_));
 DFF_X1 \mem[9][15]$_DFFE_PP_  (.D(_0550_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[9][15] ),
    .QN(_1759_));
 DFF_X1 \mem[9][16]$_DFFE_PP_  (.D(_0551_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[9][16] ),
    .QN(_1758_));
 DFF_X1 \mem[9][17]$_DFFE_PP_  (.D(_0552_),
    .CK(clknet_leaf_43_clk),
    .Q(\mem[9][17] ),
    .QN(_1757_));
 DFF_X1 \mem[9][18]$_DFFE_PP_  (.D(_0553_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[9][18] ),
    .QN(_1756_));
 DFF_X1 \mem[9][19]$_DFFE_PP_  (.D(_0554_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[9][19] ),
    .QN(_1755_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0555_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[9][1] ),
    .QN(_1754_));
 DFF_X1 \mem[9][20]$_DFFE_PP_  (.D(_0556_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[9][20] ),
    .QN(_1753_));
 DFF_X1 \mem[9][21]$_DFFE_PP_  (.D(_0557_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[9][21] ),
    .QN(_1752_));
 DFF_X1 \mem[9][22]$_DFFE_PP_  (.D(_0558_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[9][22] ),
    .QN(_1751_));
 DFF_X1 \mem[9][23]$_DFFE_PP_  (.D(_0559_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[9][23] ),
    .QN(_1750_));
 DFF_X1 \mem[9][24]$_DFFE_PP_  (.D(_0560_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[9][24] ),
    .QN(_1749_));
 DFF_X1 \mem[9][25]$_DFFE_PP_  (.D(_0561_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[9][25] ),
    .QN(_1748_));
 DFF_X1 \mem[9][26]$_DFFE_PP_  (.D(_0562_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[9][26] ),
    .QN(_1747_));
 DFF_X1 \mem[9][27]$_DFFE_PP_  (.D(_0563_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[9][27] ),
    .QN(_1746_));
 DFF_X1 \mem[9][28]$_DFFE_PP_  (.D(_0564_),
    .CK(clknet_leaf_79_clk),
    .Q(\mem[9][28] ),
    .QN(_1745_));
 DFF_X1 \mem[9][29]$_DFFE_PP_  (.D(_0565_),
    .CK(clknet_leaf_79_clk),
    .Q(\mem[9][29] ),
    .QN(_1744_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0566_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[9][2] ),
    .QN(_1743_));
 DFF_X1 \mem[9][30]$_DFFE_PP_  (.D(_0567_),
    .CK(clknet_leaf_78_clk),
    .Q(\mem[9][30] ),
    .QN(_1742_));
 DFF_X1 \mem[9][31]$_DFFE_PP_  (.D(_0568_),
    .CK(clknet_leaf_77_clk),
    .Q(\mem[9][31] ),
    .QN(_1741_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0569_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[9][3] ),
    .QN(_1740_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0570_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[9][4] ),
    .QN(_1739_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0571_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[9][5] ),
    .QN(_1738_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0572_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[9][6] ),
    .QN(_1737_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0573_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[9][7] ),
    .QN(_1736_));
 DFF_X1 \mem[9][8]$_DFFE_PP_  (.D(_0574_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[9][8] ),
    .QN(_1735_));
 DFF_X1 \mem[9][9]$_DFFE_PP_  (.D(_0575_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[9][9] ),
    .QN(_1734_));
 DFF_X2 \rd_ptr[0]$_SDFFE_PN0P_  (.D(_0576_),
    .CK(clknet_leaf_36_clk),
    .Q(\rd_ptr[0] ),
    .QN(_0006_));
 DFF_X1 \rd_ptr[1]$_SDFFE_PN0P_  (.D(_0011_),
    .CK(clknet_leaf_35_clk),
    .Q(\rd_ptr[1] ),
    .QN(_2299_));
 DFF_X1 \rd_ptr[2]$_SDFFE_PN0P_  (.D(_0012_),
    .CK(clknet_leaf_35_clk),
    .Q(\rd_ptr[2] ),
    .QN(_2307_));
 DFF_X1 \rd_ptr[3]$_SDFFE_PN0P_  (.D(_0013_),
    .CK(clknet_leaf_36_clk),
    .Q(\rd_ptr[3] ),
    .QN(_2302_));
 DFF_X1 \rd_ptr[4]$_SDFFE_PN0P_  (.D(_0577_),
    .CK(clknet_leaf_36_clk),
    .Q(\rd_ptr[4] ),
    .QN(_1733_));
 DFF_X2 \wr_ptr[0]$_SDFFE_PN0P_  (.D(_0578_),
    .CK(clknet_leaf_36_clk),
    .Q(\wr_ptr[0] ),
    .QN(_0004_));
 DFF_X2 \wr_ptr[1]$_SDFFE_PN0P_  (.D(_0579_),
    .CK(clknet_leaf_32_clk),
    .Q(\wr_ptr[1] ),
    .QN(_2312_));
 DFF_X1 \wr_ptr[2]$_SDFFE_PN0P_  (.D(_0580_),
    .CK(clknet_leaf_35_clk),
    .Q(\wr_ptr[2] ),
    .QN(_1732_));
 DFF_X1 \wr_ptr[3]$_SDFFE_PN0P_  (.D(_0581_),
    .CK(clknet_leaf_35_clk),
    .Q(\wr_ptr[3] ),
    .QN(_1731_));
 DFF_X1 \wr_ptr[4]$_SDFFE_PN0P_  (.D(_0582_),
    .CK(clknet_leaf_36_clk),
    .Q(\wr_ptr[4] ),
    .QN(_1730_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_135 ();
 BUF_X1 input1 (.A(clear_errors),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(almost_empty));
 BUF_X1 output3 (.A(net3),
    .Z(almost_full));
 BUF_X1 output4 (.A(net4),
    .Z(data_count[0]));
 BUF_X1 output5 (.A(net5),
    .Z(data_count[1]));
 BUF_X1 output6 (.A(net6),
    .Z(data_count[2]));
 BUF_X1 output7 (.A(net7),
    .Z(data_count[3]));
 BUF_X1 output8 (.A(net8),
    .Z(data_count[4]));
 BUF_X1 output9 (.A(net9),
    .Z(empty));
 BUF_X1 output10 (.A(net10),
    .Z(error_count[0]));
 BUF_X1 output11 (.A(net11),
    .Z(error_count[10]));
 BUF_X1 output12 (.A(net12),
    .Z(error_count[11]));
 BUF_X1 output13 (.A(net13),
    .Z(error_count[12]));
 BUF_X1 output14 (.A(net14),
    .Z(error_count[13]));
 BUF_X1 output15 (.A(net15),
    .Z(error_count[14]));
 BUF_X1 output16 (.A(net16),
    .Z(error_count[15]));
 BUF_X1 output17 (.A(net17),
    .Z(error_count[1]));
 BUF_X1 output18 (.A(net18),
    .Z(error_count[2]));
 BUF_X1 output19 (.A(net19),
    .Z(error_count[3]));
 BUF_X1 output20 (.A(net20),
    .Z(error_count[4]));
 BUF_X1 output21 (.A(net21),
    .Z(error_count[5]));
 BUF_X1 output22 (.A(net22),
    .Z(error_count[6]));
 BUF_X1 output23 (.A(net23),
    .Z(error_count[7]));
 BUF_X1 output24 (.A(net24),
    .Z(error_count[8]));
 BUF_X1 output25 (.A(net25),
    .Z(error_count[9]));
 BUF_X1 output26 (.A(net26),
    .Z(error_detected));
 BUF_X1 output27 (.A(net27),
    .Z(full));
 BUF_X1 output28 (.A(net28),
    .Z(overflow_detected));
 BUF_X1 output29 (.A(net29),
    .Z(rd_data[0]));
 BUF_X1 output30 (.A(net30),
    .Z(rd_data[10]));
 BUF_X1 output31 (.A(net31),
    .Z(rd_data[11]));
 BUF_X1 output32 (.A(net32),
    .Z(rd_data[12]));
 BUF_X1 output33 (.A(net33),
    .Z(rd_data[13]));
 BUF_X1 output34 (.A(net34),
    .Z(rd_data[14]));
 BUF_X1 output35 (.A(net35),
    .Z(rd_data[15]));
 BUF_X1 output36 (.A(net36),
    .Z(rd_data[16]));
 BUF_X1 output37 (.A(net37),
    .Z(rd_data[17]));
 BUF_X1 output38 (.A(net38),
    .Z(rd_data[18]));
 BUF_X1 output39 (.A(net39),
    .Z(rd_data[19]));
 BUF_X1 output40 (.A(net40),
    .Z(rd_data[1]));
 BUF_X1 output41 (.A(net41),
    .Z(rd_data[20]));
 BUF_X1 output42 (.A(net42),
    .Z(rd_data[21]));
 BUF_X1 output43 (.A(net43),
    .Z(rd_data[22]));
 BUF_X1 output44 (.A(net44),
    .Z(rd_data[23]));
 BUF_X1 output45 (.A(net45),
    .Z(rd_data[24]));
 BUF_X1 output46 (.A(net46),
    .Z(rd_data[25]));
 BUF_X1 output47 (.A(net47),
    .Z(rd_data[26]));
 BUF_X1 output48 (.A(net48),
    .Z(rd_data[27]));
 BUF_X1 output49 (.A(net49),
    .Z(rd_data[28]));
 BUF_X1 output50 (.A(net50),
    .Z(rd_data[29]));
 BUF_X1 output51 (.A(net51),
    .Z(rd_data[2]));
 BUF_X1 output52 (.A(net52),
    .Z(rd_data[30]));
 BUF_X2 output53 (.A(net53),
    .Z(rd_data[31]));
 BUF_X2 output54 (.A(net54),
    .Z(rd_data[3]));
 BUF_X1 output55 (.A(net55),
    .Z(rd_data[4]));
 BUF_X1 output56 (.A(net56),
    .Z(rd_data[5]));
 BUF_X2 output57 (.A(net57),
    .Z(rd_data[6]));
 BUF_X1 output58 (.A(net58),
    .Z(rd_data[7]));
 BUF_X1 output59 (.A(net59),
    .Z(rd_data[8]));
 BUF_X1 output60 (.A(net60),
    .Z(rd_data[9]));
 BUF_X1 output61 (.A(net61),
    .Z(rd_valid));
 BUF_X1 output62 (.A(net62),
    .Z(underflow_detected));
 BUF_X1 output63 (.A(net63),
    .Z(wr_ready));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 CLKBUF_X3 clkload0 (.A(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkload1 (.A(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkload2 (.A(clknet_3_4__leaf_clk));
 INV_X2 clkload3 (.A(clknet_3_6__leaf_clk));
 INV_X2 clkload4 (.A(clknet_3_7__leaf_clk));
 CLKBUF_X1 clkload5 (.A(clknet_leaf_0_clk));
 INV_X1 clkload6 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload7 (.A(clknet_leaf_72_clk));
 CLKBUF_X1 clkload8 (.A(clknet_leaf_73_clk));
 CLKBUF_X1 clkload9 (.A(clknet_leaf_75_clk));
 INV_X1 clkload10 (.A(clknet_leaf_76_clk));
 CLKBUF_X1 clkload11 (.A(clknet_leaf_77_clk));
 INV_X1 clkload12 (.A(clknet_leaf_79_clk));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_2_clk));
 CLKBUF_X1 clkload14 (.A(clknet_leaf_3_clk));
 INV_X1 clkload15 (.A(clknet_leaf_5_clk));
 INV_X1 clkload16 (.A(clknet_leaf_6_clk));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_7_clk));
 CLKBUF_X1 clkload18 (.A(clknet_leaf_8_clk));
 INV_X2 clkload19 (.A(clknet_leaf_68_clk));
 INV_X1 clkload20 (.A(clknet_leaf_69_clk));
 CLKBUF_X1 clkload21 (.A(clknet_leaf_70_clk));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_56_clk));
 CLKBUF_X1 clkload23 (.A(clknet_leaf_57_clk));
 INV_X1 clkload24 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_59_clk));
 INV_X1 clkload26 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload27 (.A(clknet_leaf_62_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_64_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_65_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_47_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_48_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_49_clk));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_52_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload35 (.A(clknet_leaf_9_clk));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload37 (.A(clknet_leaf_11_clk));
 CLKBUF_X1 clkload38 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload39 (.A(clknet_leaf_13_clk));
 CLKBUF_X1 clkload40 (.A(clknet_leaf_14_clk));
 CLKBUF_X1 clkload41 (.A(clknet_leaf_16_clk));
 CLKBUF_X1 clkload42 (.A(clknet_leaf_28_clk));
 CLKBUF_X1 clkload43 (.A(clknet_leaf_17_clk));
 CLKBUF_X1 clkload44 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload45 (.A(clknet_leaf_23_clk));
 CLKBUF_X1 clkload46 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_26_clk));
 INV_X1 clkload48 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload49 (.A(clknet_leaf_31_clk));
 CLKBUF_X1 clkload50 (.A(clknet_leaf_40_clk));
 INV_X1 clkload51 (.A(clknet_leaf_41_clk));
 INV_X1 clkload52 (.A(clknet_leaf_42_clk));
 CLKBUF_X1 clkload53 (.A(clknet_leaf_43_clk));
 INV_X1 clkload54 (.A(clknet_leaf_45_clk));
 CLKBUF_X1 clkload55 (.A(clknet_leaf_46_clk));
 INV_X1 clkload56 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_34_clk));
 CLKBUF_X1 clkload59 (.A(clknet_leaf_35_clk));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload61 (.A(clknet_leaf_38_clk));
 INV_X1 clkload62 (.A(clknet_leaf_39_clk));
 BUF_X1 rebuffer1 (.A(_2320_),
    .Z(net64));
 BUF_X1 rebuffer2 (.A(\rd_ptr[0] ),
    .Z(net65));
 BUF_X32 clone1 (.A(_0607_),
    .Z(net66));
 BUF_X16 clone2 (.A(_0607_),
    .Z(net67));
 BUF_X16 clone3 (.A(_0606_),
    .Z(net68));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_33 ();
 FILLCELL_X1 FILLER_0_37 ();
 FILLCELL_X2 FILLER_0_42 ();
 FILLCELL_X8 FILLER_0_48 ();
 FILLCELL_X2 FILLER_0_56 ();
 FILLCELL_X16 FILLER_0_75 ();
 FILLCELL_X2 FILLER_0_91 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X8 FILLER_0_113 ();
 FILLCELL_X2 FILLER_0_121 ();
 FILLCELL_X1 FILLER_0_140 ();
 FILLCELL_X16 FILLER_0_144 ();
 FILLCELL_X4 FILLER_0_160 ();
 FILLCELL_X2 FILLER_0_164 ();
 FILLCELL_X1 FILLER_0_166 ();
 FILLCELL_X16 FILLER_0_171 ();
 FILLCELL_X4 FILLER_0_187 ();
 FILLCELL_X2 FILLER_0_191 ();
 FILLCELL_X1 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_198 ();
 FILLCELL_X2 FILLER_0_230 ();
 FILLCELL_X16 FILLER_0_236 ();
 FILLCELL_X8 FILLER_0_252 ();
 FILLCELL_X4 FILLER_0_260 ();
 FILLCELL_X2 FILLER_0_264 ();
 FILLCELL_X1 FILLER_0_266 ();
 FILLCELL_X4 FILLER_0_271 ();
 FILLCELL_X2 FILLER_0_275 ();
 FILLCELL_X1 FILLER_0_277 ();
 FILLCELL_X16 FILLER_0_282 ();
 FILLCELL_X8 FILLER_0_298 ();
 FILLCELL_X1 FILLER_0_306 ();
 FILLCELL_X32 FILLER_0_311 ();
 FILLCELL_X4 FILLER_0_343 ();
 FILLCELL_X2 FILLER_0_347 ();
 FILLCELL_X1 FILLER_0_349 ();
 FILLCELL_X4 FILLER_0_367 ();
 FILLCELL_X16 FILLER_0_374 ();
 FILLCELL_X4 FILLER_0_390 ();
 FILLCELL_X2 FILLER_0_411 ();
 FILLCELL_X32 FILLER_0_420 ();
 FILLCELL_X16 FILLER_0_452 ();
 FILLCELL_X8 FILLER_0_468 ();
 FILLCELL_X4 FILLER_0_476 ();
 FILLCELL_X16 FILLER_0_484 ();
 FILLCELL_X4 FILLER_0_500 ();
 FILLCELL_X1 FILLER_0_504 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_41 ();
 FILLCELL_X1 FILLER_1_45 ();
 FILLCELL_X2 FILLER_1_63 ();
 FILLCELL_X4 FILLER_1_72 ();
 FILLCELL_X4 FILLER_1_93 ();
 FILLCELL_X1 FILLER_1_97 ();
 FILLCELL_X8 FILLER_1_115 ();
 FILLCELL_X2 FILLER_1_123 ();
 FILLCELL_X4 FILLER_1_132 ();
 FILLCELL_X1 FILLER_1_136 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X4 FILLER_1_193 ();
 FILLCELL_X4 FILLER_1_214 ();
 FILLCELL_X2 FILLER_1_218 ();
 FILLCELL_X8 FILLER_1_237 ();
 FILLCELL_X8 FILLER_1_262 ();
 FILLCELL_X4 FILLER_1_270 ();
 FILLCELL_X2 FILLER_1_274 ();
 FILLCELL_X8 FILLER_1_298 ();
 FILLCELL_X1 FILLER_1_306 ();
 FILLCELL_X4 FILLER_1_324 ();
 FILLCELL_X1 FILLER_1_328 ();
 FILLCELL_X2 FILLER_1_360 ();
 FILLCELL_X1 FILLER_1_362 ();
 FILLCELL_X2 FILLER_1_411 ();
 FILLCELL_X1 FILLER_1_413 ();
 FILLCELL_X8 FILLER_1_418 ();
 FILLCELL_X1 FILLER_1_426 ();
 FILLCELL_X32 FILLER_1_448 ();
 FILLCELL_X16 FILLER_1_480 ();
 FILLCELL_X8 FILLER_1_496 ();
 FILLCELL_X1 FILLER_1_504 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X1 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_57 ();
 FILLCELL_X1 FILLER_2_59 ();
 FILLCELL_X1 FILLER_2_74 ();
 FILLCELL_X2 FILLER_2_82 ();
 FILLCELL_X4 FILLER_2_115 ();
 FILLCELL_X2 FILLER_2_119 ();
 FILLCELL_X1 FILLER_2_121 ();
 FILLCELL_X4 FILLER_2_139 ();
 FILLCELL_X2 FILLER_2_143 ();
 FILLCELL_X1 FILLER_2_145 ();
 FILLCELL_X4 FILLER_2_211 ();
 FILLCELL_X1 FILLER_2_215 ();
 FILLCELL_X4 FILLER_2_240 ();
 FILLCELL_X2 FILLER_2_244 ();
 FILLCELL_X4 FILLER_2_270 ();
 FILLCELL_X1 FILLER_2_298 ();
 FILLCELL_X8 FILLER_2_316 ();
 FILLCELL_X8 FILLER_2_352 ();
 FILLCELL_X2 FILLER_2_360 ();
 FILLCELL_X8 FILLER_2_369 ();
 FILLCELL_X2 FILLER_2_377 ();
 FILLCELL_X4 FILLER_2_386 ();
 FILLCELL_X2 FILLER_2_390 ();
 FILLCELL_X1 FILLER_2_392 ();
 FILLCELL_X4 FILLER_2_397 ();
 FILLCELL_X4 FILLER_2_408 ();
 FILLCELL_X2 FILLER_2_412 ();
 FILLCELL_X1 FILLER_2_421 ();
 FILLCELL_X4 FILLER_2_446 ();
 FILLCELL_X1 FILLER_2_450 ();
 FILLCELL_X8 FILLER_2_492 ();
 FILLCELL_X4 FILLER_2_500 ();
 FILLCELL_X1 FILLER_2_504 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_33 ();
 FILLCELL_X2 FILLER_3_58 ();
 FILLCELL_X1 FILLER_3_77 ();
 FILLCELL_X8 FILLER_3_83 ();
 FILLCELL_X1 FILLER_3_91 ();
 FILLCELL_X4 FILLER_3_99 ();
 FILLCELL_X2 FILLER_3_103 ();
 FILLCELL_X1 FILLER_3_105 ();
 FILLCELL_X8 FILLER_3_113 ();
 FILLCELL_X1 FILLER_3_121 ();
 FILLCELL_X8 FILLER_3_136 ();
 FILLCELL_X2 FILLER_3_144 ();
 FILLCELL_X1 FILLER_3_146 ();
 FILLCELL_X1 FILLER_3_154 ();
 FILLCELL_X2 FILLER_3_162 ();
 FILLCELL_X1 FILLER_3_164 ();
 FILLCELL_X4 FILLER_3_179 ();
 FILLCELL_X1 FILLER_3_207 ();
 FILLCELL_X4 FILLER_3_215 ();
 FILLCELL_X2 FILLER_3_219 ();
 FILLCELL_X1 FILLER_3_221 ();
 FILLCELL_X16 FILLER_3_236 ();
 FILLCELL_X8 FILLER_3_266 ();
 FILLCELL_X4 FILLER_3_286 ();
 FILLCELL_X1 FILLER_3_290 ();
 FILLCELL_X1 FILLER_3_298 ();
 FILLCELL_X1 FILLER_3_306 ();
 FILLCELL_X1 FILLER_3_314 ();
 FILLCELL_X1 FILLER_3_322 ();
 FILLCELL_X1 FILLER_3_340 ();
 FILLCELL_X4 FILLER_3_358 ();
 FILLCELL_X1 FILLER_3_362 ();
 FILLCELL_X8 FILLER_3_370 ();
 FILLCELL_X1 FILLER_3_378 ();
 FILLCELL_X8 FILLER_3_396 ();
 FILLCELL_X1 FILLER_3_404 ();
 FILLCELL_X4 FILLER_3_422 ();
 FILLCELL_X1 FILLER_3_426 ();
 FILLCELL_X16 FILLER_3_434 ();
 FILLCELL_X2 FILLER_3_450 ();
 FILLCELL_X1 FILLER_3_452 ();
 FILLCELL_X8 FILLER_3_467 ();
 FILLCELL_X4 FILLER_3_499 ();
 FILLCELL_X2 FILLER_3_503 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X4 FILLER_4_33 ();
 FILLCELL_X2 FILLER_4_37 ();
 FILLCELL_X1 FILLER_4_39 ();
 FILLCELL_X8 FILLER_4_64 ();
 FILLCELL_X16 FILLER_4_89 ();
 FILLCELL_X8 FILLER_4_105 ();
 FILLCELL_X2 FILLER_4_113 ();
 FILLCELL_X1 FILLER_4_115 ();
 FILLCELL_X32 FILLER_4_121 ();
 FILLCELL_X32 FILLER_4_153 ();
 FILLCELL_X4 FILLER_4_185 ();
 FILLCELL_X1 FILLER_4_189 ();
 FILLCELL_X32 FILLER_4_195 ();
 FILLCELL_X16 FILLER_4_227 ();
 FILLCELL_X8 FILLER_4_243 ();
 FILLCELL_X4 FILLER_4_251 ();
 FILLCELL_X1 FILLER_4_255 ();
 FILLCELL_X8 FILLER_4_273 ();
 FILLCELL_X4 FILLER_4_281 ();
 FILLCELL_X2 FILLER_4_285 ();
 FILLCELL_X1 FILLER_4_287 ();
 FILLCELL_X16 FILLER_4_293 ();
 FILLCELL_X4 FILLER_4_309 ();
 FILLCELL_X2 FILLER_4_313 ();
 FILLCELL_X1 FILLER_4_315 ();
 FILLCELL_X8 FILLER_4_323 ();
 FILLCELL_X2 FILLER_4_360 ();
 FILLCELL_X4 FILLER_4_386 ();
 FILLCELL_X1 FILLER_4_390 ();
 FILLCELL_X2 FILLER_4_399 ();
 FILLCELL_X4 FILLER_4_408 ();
 FILLCELL_X2 FILLER_4_412 ();
 FILLCELL_X1 FILLER_4_414 ();
 FILLCELL_X8 FILLER_4_422 ();
 FILLCELL_X16 FILLER_4_444 ();
 FILLCELL_X8 FILLER_4_460 ();
 FILLCELL_X8 FILLER_4_493 ();
 FILLCELL_X4 FILLER_4_501 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_41 ();
 FILLCELL_X2 FILLER_5_45 ();
 FILLCELL_X1 FILLER_5_47 ();
 FILLCELL_X1 FILLER_5_55 ();
 FILLCELL_X4 FILLER_5_63 ();
 FILLCELL_X1 FILLER_5_67 ();
 FILLCELL_X16 FILLER_5_92 ();
 FILLCELL_X2 FILLER_5_108 ();
 FILLCELL_X8 FILLER_5_137 ();
 FILLCELL_X1 FILLER_5_145 ();
 FILLCELL_X1 FILLER_5_187 ();
 FILLCELL_X1 FILLER_5_212 ();
 FILLCELL_X8 FILLER_5_230 ();
 FILLCELL_X8 FILLER_5_246 ();
 FILLCELL_X8 FILLER_5_278 ();
 FILLCELL_X1 FILLER_5_286 ();
 FILLCELL_X8 FILLER_5_304 ();
 FILLCELL_X8 FILLER_5_329 ();
 FILLCELL_X4 FILLER_5_337 ();
 FILLCELL_X1 FILLER_5_341 ();
 FILLCELL_X2 FILLER_5_349 ();
 FILLCELL_X1 FILLER_5_351 ();
 FILLCELL_X16 FILLER_5_359 ();
 FILLCELL_X8 FILLER_5_375 ();
 FILLCELL_X16 FILLER_5_386 ();
 FILLCELL_X2 FILLER_5_419 ();
 FILLCELL_X2 FILLER_5_458 ();
 FILLCELL_X8 FILLER_5_463 ();
 FILLCELL_X16 FILLER_5_485 ();
 FILLCELL_X4 FILLER_5_501 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_33 ();
 FILLCELL_X2 FILLER_6_37 ();
 FILLCELL_X1 FILLER_6_39 ();
 FILLCELL_X4 FILLER_6_71 ();
 FILLCELL_X8 FILLER_6_113 ();
 FILLCELL_X1 FILLER_6_121 ();
 FILLCELL_X2 FILLER_6_139 ();
 FILLCELL_X1 FILLER_6_141 ();
 FILLCELL_X4 FILLER_6_166 ();
 FILLCELL_X2 FILLER_6_170 ();
 FILLCELL_X8 FILLER_6_189 ();
 FILLCELL_X4 FILLER_6_214 ();
 FILLCELL_X16 FILLER_6_242 ();
 FILLCELL_X4 FILLER_6_258 ();
 FILLCELL_X1 FILLER_6_262 ();
 FILLCELL_X2 FILLER_6_270 ();
 FILLCELL_X1 FILLER_6_272 ();
 FILLCELL_X2 FILLER_6_292 ();
 FILLCELL_X4 FILLER_6_318 ();
 FILLCELL_X2 FILLER_6_322 ();
 FILLCELL_X1 FILLER_6_324 ();
 FILLCELL_X16 FILLER_6_332 ();
 FILLCELL_X4 FILLER_6_348 ();
 FILLCELL_X4 FILLER_6_359 ();
 FILLCELL_X2 FILLER_6_363 ();
 FILLCELL_X8 FILLER_6_368 ();
 FILLCELL_X1 FILLER_6_376 ();
 FILLCELL_X2 FILLER_6_408 ();
 FILLCELL_X4 FILLER_6_468 ();
 FILLCELL_X2 FILLER_6_472 ();
 FILLCELL_X1 FILLER_6_474 ();
 FILLCELL_X1 FILLER_6_478 ();
 FILLCELL_X2 FILLER_6_503 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_33 ();
 FILLCELL_X4 FILLER_7_61 ();
 FILLCELL_X1 FILLER_7_65 ();
 FILLCELL_X1 FILLER_7_90 ();
 FILLCELL_X2 FILLER_7_98 ();
 FILLCELL_X4 FILLER_7_117 ();
 FILLCELL_X1 FILLER_7_121 ();
 FILLCELL_X8 FILLER_7_136 ();
 FILLCELL_X4 FILLER_7_144 ();
 FILLCELL_X1 FILLER_7_148 ();
 FILLCELL_X8 FILLER_7_185 ();
 FILLCELL_X4 FILLER_7_193 ();
 FILLCELL_X8 FILLER_7_211 ();
 FILLCELL_X1 FILLER_7_219 ();
 FILLCELL_X8 FILLER_7_234 ();
 FILLCELL_X2 FILLER_7_242 ();
 FILLCELL_X2 FILLER_7_261 ();
 FILLCELL_X16 FILLER_7_268 ();
 FILLCELL_X8 FILLER_7_284 ();
 FILLCELL_X1 FILLER_7_292 ();
 FILLCELL_X2 FILLER_7_317 ();
 FILLCELL_X1 FILLER_7_319 ();
 FILLCELL_X4 FILLER_7_334 ();
 FILLCELL_X2 FILLER_7_338 ();
 FILLCELL_X4 FILLER_7_357 ();
 FILLCELL_X8 FILLER_7_364 ();
 FILLCELL_X1 FILLER_7_372 ();
 FILLCELL_X16 FILLER_7_393 ();
 FILLCELL_X4 FILLER_7_409 ();
 FILLCELL_X2 FILLER_7_413 ();
 FILLCELL_X2 FILLER_7_422 ();
 FILLCELL_X1 FILLER_7_424 ();
 FILLCELL_X8 FILLER_7_432 ();
 FILLCELL_X2 FILLER_7_443 ();
 FILLCELL_X2 FILLER_7_452 ();
 FILLCELL_X1 FILLER_7_454 ();
 FILLCELL_X2 FILLER_7_462 ();
 FILLCELL_X1 FILLER_7_464 ();
 FILLCELL_X4 FILLER_7_492 ();
 FILLCELL_X2 FILLER_7_496 ();
 FILLCELL_X1 FILLER_7_498 ();
 FILLCELL_X2 FILLER_7_502 ();
 FILLCELL_X1 FILLER_7_504 ();
 FILLCELL_X8 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_9 ();
 FILLCELL_X1 FILLER_8_11 ();
 FILLCELL_X8 FILLER_8_29 ();
 FILLCELL_X4 FILLER_8_37 ();
 FILLCELL_X2 FILLER_8_41 ();
 FILLCELL_X8 FILLER_8_74 ();
 FILLCELL_X4 FILLER_8_82 ();
 FILLCELL_X2 FILLER_8_86 ();
 FILLCELL_X8 FILLER_8_91 ();
 FILLCELL_X4 FILLER_8_99 ();
 FILLCELL_X16 FILLER_8_110 ();
 FILLCELL_X4 FILLER_8_126 ();
 FILLCELL_X2 FILLER_8_130 ();
 FILLCELL_X1 FILLER_8_132 ();
 FILLCELL_X16 FILLER_8_136 ();
 FILLCELL_X8 FILLER_8_152 ();
 FILLCELL_X1 FILLER_8_160 ();
 FILLCELL_X8 FILLER_8_167 ();
 FILLCELL_X2 FILLER_8_175 ();
 FILLCELL_X1 FILLER_8_177 ();
 FILLCELL_X16 FILLER_8_181 ();
 FILLCELL_X8 FILLER_8_197 ();
 FILLCELL_X2 FILLER_8_205 ();
 FILLCELL_X1 FILLER_8_207 ();
 FILLCELL_X8 FILLER_8_211 ();
 FILLCELL_X4 FILLER_8_219 ();
 FILLCELL_X2 FILLER_8_223 ();
 FILLCELL_X1 FILLER_8_225 ();
 FILLCELL_X8 FILLER_8_229 ();
 FILLCELL_X4 FILLER_8_237 ();
 FILLCELL_X1 FILLER_8_241 ();
 FILLCELL_X4 FILLER_8_259 ();
 FILLCELL_X2 FILLER_8_263 ();
 FILLCELL_X32 FILLER_8_268 ();
 FILLCELL_X16 FILLER_8_300 ();
 FILLCELL_X8 FILLER_8_316 ();
 FILLCELL_X4 FILLER_8_324 ();
 FILLCELL_X2 FILLER_8_328 ();
 FILLCELL_X4 FILLER_8_337 ();
 FILLCELL_X1 FILLER_8_341 ();
 FILLCELL_X2 FILLER_8_359 ();
 FILLCELL_X8 FILLER_8_368 ();
 FILLCELL_X2 FILLER_8_376 ();
 FILLCELL_X16 FILLER_8_392 ();
 FILLCELL_X4 FILLER_8_408 ();
 FILLCELL_X2 FILLER_8_412 ();
 FILLCELL_X32 FILLER_8_421 ();
 FILLCELL_X4 FILLER_8_453 ();
 FILLCELL_X2 FILLER_8_457 ();
 FILLCELL_X8 FILLER_8_462 ();
 FILLCELL_X4 FILLER_8_470 ();
 FILLCELL_X8 FILLER_8_491 ();
 FILLCELL_X4 FILLER_8_499 ();
 FILLCELL_X2 FILLER_8_503 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X4 FILLER_9_57 ();
 FILLCELL_X2 FILLER_9_61 ();
 FILLCELL_X1 FILLER_9_63 ();
 FILLCELL_X8 FILLER_9_67 ();
 FILLCELL_X8 FILLER_9_78 ();
 FILLCELL_X2 FILLER_9_86 ();
 FILLCELL_X8 FILLER_9_91 ();
 FILLCELL_X4 FILLER_9_99 ();
 FILLCELL_X2 FILLER_9_103 ();
 FILLCELL_X1 FILLER_9_105 ();
 FILLCELL_X2 FILLER_9_129 ();
 FILLCELL_X16 FILLER_9_151 ();
 FILLCELL_X8 FILLER_9_167 ();
 FILLCELL_X2 FILLER_9_175 ();
 FILLCELL_X1 FILLER_9_177 ();
 FILLCELL_X2 FILLER_9_195 ();
 FILLCELL_X4 FILLER_9_204 ();
 FILLCELL_X2 FILLER_9_208 ();
 FILLCELL_X2 FILLER_9_237 ();
 FILLCELL_X1 FILLER_9_239 ();
 FILLCELL_X2 FILLER_9_258 ();
 FILLCELL_X8 FILLER_9_267 ();
 FILLCELL_X2 FILLER_9_275 ();
 FILLCELL_X1 FILLER_9_277 ();
 FILLCELL_X1 FILLER_9_295 ();
 FILLCELL_X2 FILLER_9_313 ();
 FILLCELL_X1 FILLER_9_315 ();
 FILLCELL_X2 FILLER_9_333 ();
 FILLCELL_X4 FILLER_9_342 ();
 FILLCELL_X1 FILLER_9_355 ();
 FILLCELL_X32 FILLER_9_373 ();
 FILLCELL_X4 FILLER_9_405 ();
 FILLCELL_X16 FILLER_9_426 ();
 FILLCELL_X4 FILLER_9_442 ();
 FILLCELL_X2 FILLER_9_453 ();
 FILLCELL_X8 FILLER_9_462 ();
 FILLCELL_X4 FILLER_9_470 ();
 FILLCELL_X2 FILLER_9_474 ();
 FILLCELL_X1 FILLER_9_476 ();
 FILLCELL_X2 FILLER_9_484 ();
 FILLCELL_X2 FILLER_9_503 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_9 ();
 FILLCELL_X2 FILLER_10_13 ();
 FILLCELL_X16 FILLER_10_29 ();
 FILLCELL_X4 FILLER_10_45 ();
 FILLCELL_X4 FILLER_10_52 ();
 FILLCELL_X1 FILLER_10_56 ();
 FILLCELL_X8 FILLER_10_64 ();
 FILLCELL_X4 FILLER_10_72 ();
 FILLCELL_X8 FILLER_10_89 ();
 FILLCELL_X1 FILLER_10_97 ();
 FILLCELL_X1 FILLER_10_129 ();
 FILLCELL_X4 FILLER_10_137 ();
 FILLCELL_X1 FILLER_10_141 ();
 FILLCELL_X1 FILLER_10_156 ();
 FILLCELL_X1 FILLER_10_180 ();
 FILLCELL_X1 FILLER_10_198 ();
 FILLCELL_X2 FILLER_10_233 ();
 FILLCELL_X4 FILLER_10_238 ();
 FILLCELL_X4 FILLER_10_259 ();
 FILLCELL_X2 FILLER_10_263 ();
 FILLCELL_X1 FILLER_10_265 ();
 FILLCELL_X8 FILLER_10_269 ();
 FILLCELL_X4 FILLER_10_277 ();
 FILLCELL_X16 FILLER_10_302 ();
 FILLCELL_X2 FILLER_10_318 ();
 FILLCELL_X1 FILLER_10_320 ();
 FILLCELL_X4 FILLER_10_338 ();
 FILLCELL_X1 FILLER_10_342 ();
 FILLCELL_X16 FILLER_10_362 ();
 FILLCELL_X1 FILLER_10_378 ();
 FILLCELL_X8 FILLER_10_413 ();
 FILLCELL_X4 FILLER_10_421 ();
 FILLCELL_X2 FILLER_10_425 ();
 FILLCELL_X8 FILLER_10_434 ();
 FILLCELL_X8 FILLER_10_466 ();
 FILLCELL_X2 FILLER_10_474 ();
 FILLCELL_X4 FILLER_10_500 ();
 FILLCELL_X1 FILLER_10_504 ();
 FILLCELL_X16 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_17 ();
 FILLCELL_X2 FILLER_11_25 ();
 FILLCELL_X2 FILLER_11_75 ();
 FILLCELL_X2 FILLER_11_97 ();
 FILLCELL_X16 FILLER_11_109 ();
 FILLCELL_X2 FILLER_11_132 ();
 FILLCELL_X8 FILLER_11_137 ();
 FILLCELL_X4 FILLER_11_145 ();
 FILLCELL_X2 FILLER_11_149 ();
 FILLCELL_X1 FILLER_11_151 ();
 FILLCELL_X16 FILLER_11_166 ();
 FILLCELL_X8 FILLER_11_182 ();
 FILLCELL_X1 FILLER_11_190 ();
 FILLCELL_X2 FILLER_11_198 ();
 FILLCELL_X1 FILLER_11_200 ();
 FILLCELL_X8 FILLER_11_212 ();
 FILLCELL_X2 FILLER_11_220 ();
 FILLCELL_X1 FILLER_11_222 ();
 FILLCELL_X2 FILLER_11_233 ();
 FILLCELL_X4 FILLER_11_257 ();
 FILLCELL_X2 FILLER_11_261 ();
 FILLCELL_X4 FILLER_11_275 ();
 FILLCELL_X2 FILLER_11_279 ();
 FILLCELL_X16 FILLER_11_284 ();
 FILLCELL_X1 FILLER_11_300 ();
 FILLCELL_X1 FILLER_11_304 ();
 FILLCELL_X8 FILLER_11_329 ();
 FILLCELL_X2 FILLER_11_337 ();
 FILLCELL_X1 FILLER_11_339 ();
 FILLCELL_X1 FILLER_11_343 ();
 FILLCELL_X1 FILLER_11_364 ();
 FILLCELL_X4 FILLER_11_368 ();
 FILLCELL_X1 FILLER_11_372 ();
 FILLCELL_X2 FILLER_11_390 ();
 FILLCELL_X1 FILLER_11_392 ();
 FILLCELL_X1 FILLER_11_400 ();
 FILLCELL_X4 FILLER_11_408 ();
 FILLCELL_X4 FILLER_11_422 ();
 FILLCELL_X8 FILLER_11_443 ();
 FILLCELL_X1 FILLER_11_451 ();
 FILLCELL_X8 FILLER_11_469 ();
 FILLCELL_X4 FILLER_11_477 ();
 FILLCELL_X2 FILLER_11_481 ();
 FILLCELL_X8 FILLER_11_490 ();
 FILLCELL_X4 FILLER_11_498 ();
 FILLCELL_X2 FILLER_11_502 ();
 FILLCELL_X1 FILLER_11_504 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_46 ();
 FILLCELL_X4 FILLER_12_54 ();
 FILLCELL_X2 FILLER_12_58 ();
 FILLCELL_X1 FILLER_12_60 ();
 FILLCELL_X4 FILLER_12_68 ();
 FILLCELL_X4 FILLER_12_86 ();
 FILLCELL_X1 FILLER_12_90 ();
 FILLCELL_X16 FILLER_12_98 ();
 FILLCELL_X8 FILLER_12_114 ();
 FILLCELL_X2 FILLER_12_122 ();
 FILLCELL_X1 FILLER_12_124 ();
 FILLCELL_X1 FILLER_12_128 ();
 FILLCELL_X8 FILLER_12_134 ();
 FILLCELL_X16 FILLER_12_149 ();
 FILLCELL_X8 FILLER_12_165 ();
 FILLCELL_X32 FILLER_12_183 ();
 FILLCELL_X8 FILLER_12_215 ();
 FILLCELL_X4 FILLER_12_223 ();
 FILLCELL_X1 FILLER_12_239 ();
 FILLCELL_X4 FILLER_12_261 ();
 FILLCELL_X2 FILLER_12_265 ();
 FILLCELL_X16 FILLER_12_270 ();
 FILLCELL_X1 FILLER_12_286 ();
 FILLCELL_X16 FILLER_12_295 ();
 FILLCELL_X1 FILLER_12_311 ();
 FILLCELL_X4 FILLER_12_326 ();
 FILLCELL_X2 FILLER_12_330 ();
 FILLCELL_X1 FILLER_12_332 ();
 FILLCELL_X2 FILLER_12_336 ();
 FILLCELL_X1 FILLER_12_338 ();
 FILLCELL_X8 FILLER_12_342 ();
 FILLCELL_X8 FILLER_12_367 ();
 FILLCELL_X1 FILLER_12_375 ();
 FILLCELL_X2 FILLER_12_388 ();
 FILLCELL_X2 FILLER_12_400 ();
 FILLCELL_X1 FILLER_12_402 ();
 FILLCELL_X32 FILLER_12_423 ();
 FILLCELL_X16 FILLER_12_455 ();
 FILLCELL_X4 FILLER_12_471 ();
 FILLCELL_X2 FILLER_12_475 ();
 FILLCELL_X1 FILLER_12_485 ();
 FILLCELL_X8 FILLER_12_493 ();
 FILLCELL_X4 FILLER_12_501 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_3 ();
 FILLCELL_X2 FILLER_13_36 ();
 FILLCELL_X1 FILLER_13_38 ();
 FILLCELL_X8 FILLER_13_49 ();
 FILLCELL_X2 FILLER_13_57 ();
 FILLCELL_X1 FILLER_13_59 ();
 FILLCELL_X4 FILLER_13_87 ();
 FILLCELL_X2 FILLER_13_91 ();
 FILLCELL_X1 FILLER_13_93 ();
 FILLCELL_X4 FILLER_13_118 ();
 FILLCELL_X2 FILLER_13_129 ();
 FILLCELL_X1 FILLER_13_155 ();
 FILLCELL_X4 FILLER_13_159 ();
 FILLCELL_X1 FILLER_13_190 ();
 FILLCELL_X2 FILLER_13_208 ();
 FILLCELL_X1 FILLER_13_210 ();
 FILLCELL_X4 FILLER_13_214 ();
 FILLCELL_X32 FILLER_13_238 ();
 FILLCELL_X4 FILLER_13_294 ();
 FILLCELL_X2 FILLER_13_301 ();
 FILLCELL_X2 FILLER_13_306 ();
 FILLCELL_X1 FILLER_13_308 ();
 FILLCELL_X4 FILLER_13_329 ();
 FILLCELL_X2 FILLER_13_333 ();
 FILLCELL_X2 FILLER_13_359 ();
 FILLCELL_X1 FILLER_13_368 ();
 FILLCELL_X2 FILLER_13_394 ();
 FILLCELL_X1 FILLER_13_396 ();
 FILLCELL_X2 FILLER_13_411 ();
 FILLCELL_X4 FILLER_13_420 ();
 FILLCELL_X2 FILLER_13_424 ();
 FILLCELL_X8 FILLER_13_450 ();
 FILLCELL_X8 FILLER_13_475 ();
 FILLCELL_X2 FILLER_13_483 ();
 FILLCELL_X2 FILLER_13_502 ();
 FILLCELL_X1 FILLER_13_504 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X16 FILLER_14_27 ();
 FILLCELL_X8 FILLER_14_43 ();
 FILLCELL_X16 FILLER_14_54 ();
 FILLCELL_X1 FILLER_14_70 ();
 FILLCELL_X4 FILLER_14_92 ();
 FILLCELL_X1 FILLER_14_96 ();
 FILLCELL_X1 FILLER_14_128 ();
 FILLCELL_X4 FILLER_14_146 ();
 FILLCELL_X2 FILLER_14_164 ();
 FILLCELL_X1 FILLER_14_173 ();
 FILLCELL_X8 FILLER_14_181 ();
 FILLCELL_X4 FILLER_14_189 ();
 FILLCELL_X1 FILLER_14_210 ();
 FILLCELL_X2 FILLER_14_228 ();
 FILLCELL_X1 FILLER_14_230 ();
 FILLCELL_X4 FILLER_14_238 ();
 FILLCELL_X2 FILLER_14_242 ();
 FILLCELL_X1 FILLER_14_244 ();
 FILLCELL_X1 FILLER_14_269 ();
 FILLCELL_X4 FILLER_14_295 ();
 FILLCELL_X1 FILLER_14_306 ();
 FILLCELL_X8 FILLER_14_331 ();
 FILLCELL_X4 FILLER_14_339 ();
 FILLCELL_X1 FILLER_14_343 ();
 FILLCELL_X2 FILLER_14_351 ();
 FILLCELL_X1 FILLER_14_353 ();
 FILLCELL_X2 FILLER_14_364 ();
 FILLCELL_X2 FILLER_14_383 ();
 FILLCELL_X4 FILLER_14_392 ();
 FILLCELL_X8 FILLER_14_416 ();
 FILLCELL_X1 FILLER_14_424 ();
 FILLCELL_X8 FILLER_14_432 ();
 FILLCELL_X1 FILLER_14_440 ();
 FILLCELL_X8 FILLER_14_469 ();
 FILLCELL_X2 FILLER_14_477 ();
 FILLCELL_X2 FILLER_14_482 ();
 FILLCELL_X4 FILLER_14_501 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_5 ();
 FILLCELL_X2 FILLER_15_23 ();
 FILLCELL_X4 FILLER_15_32 ();
 FILLCELL_X8 FILLER_15_67 ();
 FILLCELL_X2 FILLER_15_75 ();
 FILLCELL_X4 FILLER_15_84 ();
 FILLCELL_X8 FILLER_15_105 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X1 FILLER_15_117 ();
 FILLCELL_X2 FILLER_15_125 ();
 FILLCELL_X1 FILLER_15_127 ();
 FILLCELL_X4 FILLER_15_135 ();
 FILLCELL_X2 FILLER_15_139 ();
 FILLCELL_X2 FILLER_15_158 ();
 FILLCELL_X1 FILLER_15_160 ();
 FILLCELL_X1 FILLER_15_168 ();
 FILLCELL_X4 FILLER_15_212 ();
 FILLCELL_X2 FILLER_15_216 ();
 FILLCELL_X1 FILLER_15_218 ();
 FILLCELL_X4 FILLER_15_236 ();
 FILLCELL_X1 FILLER_15_240 ();
 FILLCELL_X1 FILLER_15_272 ();
 FILLCELL_X1 FILLER_15_287 ();
 FILLCELL_X2 FILLER_15_295 ();
 FILLCELL_X8 FILLER_15_302 ();
 FILLCELL_X2 FILLER_15_310 ();
 FILLCELL_X4 FILLER_15_329 ();
 FILLCELL_X1 FILLER_15_333 ();
 FILLCELL_X2 FILLER_15_337 ();
 FILLCELL_X1 FILLER_15_339 ();
 FILLCELL_X8 FILLER_15_364 ();
 FILLCELL_X2 FILLER_15_372 ();
 FILLCELL_X1 FILLER_15_388 ();
 FILLCELL_X1 FILLER_15_392 ();
 FILLCELL_X1 FILLER_15_400 ();
 FILLCELL_X2 FILLER_15_418 ();
 FILLCELL_X4 FILLER_15_456 ();
 FILLCELL_X2 FILLER_15_460 ();
 FILLCELL_X1 FILLER_15_462 ();
 FILLCELL_X4 FILLER_15_473 ();
 FILLCELL_X2 FILLER_15_477 ();
 FILLCELL_X1 FILLER_15_479 ();
 FILLCELL_X2 FILLER_15_483 ();
 FILLCELL_X1 FILLER_15_485 ();
 FILLCELL_X4 FILLER_15_500 ();
 FILLCELL_X1 FILLER_15_504 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X2 FILLER_16_13 ();
 FILLCELL_X2 FILLER_16_22 ();
 FILLCELL_X1 FILLER_16_24 ();
 FILLCELL_X8 FILLER_16_32 ();
 FILLCELL_X2 FILLER_16_40 ();
 FILLCELL_X4 FILLER_16_69 ();
 FILLCELL_X2 FILLER_16_73 ();
 FILLCELL_X16 FILLER_16_92 ();
 FILLCELL_X2 FILLER_16_108 ();
 FILLCELL_X1 FILLER_16_110 ();
 FILLCELL_X32 FILLER_16_128 ();
 FILLCELL_X1 FILLER_16_160 ();
 FILLCELL_X32 FILLER_16_178 ();
 FILLCELL_X2 FILLER_16_210 ();
 FILLCELL_X1 FILLER_16_212 ();
 FILLCELL_X8 FILLER_16_224 ();
 FILLCELL_X4 FILLER_16_232 ();
 FILLCELL_X2 FILLER_16_236 ();
 FILLCELL_X4 FILLER_16_243 ();
 FILLCELL_X1 FILLER_16_247 ();
 FILLCELL_X2 FILLER_16_255 ();
 FILLCELL_X1 FILLER_16_257 ();
 FILLCELL_X4 FILLER_16_275 ();
 FILLCELL_X2 FILLER_16_279 ();
 FILLCELL_X2 FILLER_16_285 ();
 FILLCELL_X1 FILLER_16_287 ();
 FILLCELL_X8 FILLER_16_295 ();
 FILLCELL_X4 FILLER_16_303 ();
 FILLCELL_X8 FILLER_16_310 ();
 FILLCELL_X4 FILLER_16_328 ();
 FILLCELL_X2 FILLER_16_332 ();
 FILLCELL_X1 FILLER_16_334 ();
 FILLCELL_X16 FILLER_16_338 ();
 FILLCELL_X1 FILLER_16_354 ();
 FILLCELL_X2 FILLER_16_372 ();
 FILLCELL_X1 FILLER_16_388 ();
 FILLCELL_X32 FILLER_16_416 ();
 FILLCELL_X1 FILLER_16_448 ();
 FILLCELL_X16 FILLER_16_452 ();
 FILLCELL_X4 FILLER_16_468 ();
 FILLCELL_X2 FILLER_16_472 ();
 FILLCELL_X16 FILLER_16_481 ();
 FILLCELL_X8 FILLER_16_497 ();
 FILLCELL_X1 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_10 ();
 FILLCELL_X16 FILLER_17_29 ();
 FILLCELL_X8 FILLER_17_45 ();
 FILLCELL_X2 FILLER_17_53 ();
 FILLCELL_X1 FILLER_17_55 ();
 FILLCELL_X16 FILLER_17_63 ();
 FILLCELL_X8 FILLER_17_79 ();
 FILLCELL_X8 FILLER_17_98 ();
 FILLCELL_X2 FILLER_17_106 ();
 FILLCELL_X1 FILLER_17_108 ();
 FILLCELL_X8 FILLER_17_133 ();
 FILLCELL_X4 FILLER_17_141 ();
 FILLCELL_X1 FILLER_17_145 ();
 FILLCELL_X16 FILLER_17_150 ();
 FILLCELL_X16 FILLER_17_190 ();
 FILLCELL_X8 FILLER_17_206 ();
 FILLCELL_X4 FILLER_17_214 ();
 FILLCELL_X1 FILLER_17_218 ();
 FILLCELL_X4 FILLER_17_236 ();
 FILLCELL_X2 FILLER_17_240 ();
 FILLCELL_X1 FILLER_17_242 ();
 FILLCELL_X32 FILLER_17_250 ();
 FILLCELL_X1 FILLER_17_282 ();
 FILLCELL_X8 FILLER_17_307 ();
 FILLCELL_X4 FILLER_17_315 ();
 FILLCELL_X1 FILLER_17_319 ();
 FILLCELL_X16 FILLER_17_349 ();
 FILLCELL_X4 FILLER_17_365 ();
 FILLCELL_X32 FILLER_17_393 ();
 FILLCELL_X8 FILLER_17_425 ();
 FILLCELL_X2 FILLER_17_440 ();
 FILLCELL_X1 FILLER_17_442 ();
 FILLCELL_X8 FILLER_17_457 ();
 FILLCELL_X1 FILLER_17_465 ();
 FILLCELL_X2 FILLER_17_483 ();
 FILLCELL_X1 FILLER_17_485 ();
 FILLCELL_X2 FILLER_17_503 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_9 ();
 FILLCELL_X2 FILLER_18_13 ();
 FILLCELL_X4 FILLER_18_26 ();
 FILLCELL_X2 FILLER_18_30 ();
 FILLCELL_X1 FILLER_18_32 ();
 FILLCELL_X1 FILLER_18_37 ();
 FILLCELL_X8 FILLER_18_52 ();
 FILLCELL_X4 FILLER_18_60 ();
 FILLCELL_X2 FILLER_18_64 ();
 FILLCELL_X1 FILLER_18_66 ();
 FILLCELL_X8 FILLER_18_74 ();
 FILLCELL_X4 FILLER_18_82 ();
 FILLCELL_X1 FILLER_18_86 ();
 FILLCELL_X2 FILLER_18_104 ();
 FILLCELL_X2 FILLER_18_137 ();
 FILLCELL_X1 FILLER_18_139 ();
 FILLCELL_X16 FILLER_18_181 ();
 FILLCELL_X8 FILLER_18_197 ();
 FILLCELL_X2 FILLER_18_205 ();
 FILLCELL_X1 FILLER_18_207 ();
 FILLCELL_X2 FILLER_18_215 ();
 FILLCELL_X1 FILLER_18_217 ();
 FILLCELL_X2 FILLER_18_242 ();
 FILLCELL_X1 FILLER_18_251 ();
 FILLCELL_X8 FILLER_18_269 ();
 FILLCELL_X4 FILLER_18_277 ();
 FILLCELL_X32 FILLER_18_326 ();
 FILLCELL_X16 FILLER_18_358 ();
 FILLCELL_X8 FILLER_18_391 ();
 FILLCELL_X2 FILLER_18_399 ();
 FILLCELL_X1 FILLER_18_401 ();
 FILLCELL_X8 FILLER_18_419 ();
 FILLCELL_X4 FILLER_18_427 ();
 FILLCELL_X2 FILLER_18_431 ();
 FILLCELL_X1 FILLER_18_433 ();
 FILLCELL_X2 FILLER_18_451 ();
 FILLCELL_X4 FILLER_18_470 ();
 FILLCELL_X4 FILLER_18_481 ();
 FILLCELL_X4 FILLER_18_492 ();
 FILLCELL_X2 FILLER_18_503 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_22 ();
 FILLCELL_X2 FILLER_19_40 ();
 FILLCELL_X8 FILLER_19_59 ();
 FILLCELL_X2 FILLER_19_67 ();
 FILLCELL_X4 FILLER_19_119 ();
 FILLCELL_X1 FILLER_19_123 ();
 FILLCELL_X4 FILLER_19_131 ();
 FILLCELL_X1 FILLER_19_135 ();
 FILLCELL_X2 FILLER_19_143 ();
 FILLCELL_X4 FILLER_19_152 ();
 FILLCELL_X1 FILLER_19_156 ();
 FILLCELL_X8 FILLER_19_164 ();
 FILLCELL_X2 FILLER_19_172 ();
 FILLCELL_X1 FILLER_19_174 ();
 FILLCELL_X4 FILLER_19_182 ();
 FILLCELL_X1 FILLER_19_193 ();
 FILLCELL_X8 FILLER_19_211 ();
 FILLCELL_X2 FILLER_19_219 ();
 FILLCELL_X1 FILLER_19_221 ();
 FILLCELL_X2 FILLER_19_229 ();
 FILLCELL_X1 FILLER_19_231 ();
 FILLCELL_X16 FILLER_19_239 ();
 FILLCELL_X1 FILLER_19_255 ();
 FILLCELL_X32 FILLER_19_277 ();
 FILLCELL_X2 FILLER_19_309 ();
 FILLCELL_X1 FILLER_19_311 ();
 FILLCELL_X8 FILLER_19_329 ();
 FILLCELL_X16 FILLER_19_378 ();
 FILLCELL_X1 FILLER_19_394 ();
 FILLCELL_X8 FILLER_19_419 ();
 FILLCELL_X4 FILLER_19_427 ();
 FILLCELL_X16 FILLER_19_453 ();
 FILLCELL_X4 FILLER_19_469 ();
 FILLCELL_X2 FILLER_19_473 ();
 FILLCELL_X8 FILLER_19_478 ();
 FILLCELL_X2 FILLER_19_503 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_9 ();
 FILLCELL_X1 FILLER_20_13 ();
 FILLCELL_X1 FILLER_20_46 ();
 FILLCELL_X4 FILLER_20_64 ();
 FILLCELL_X1 FILLER_20_75 ();
 FILLCELL_X8 FILLER_20_83 ();
 FILLCELL_X4 FILLER_20_91 ();
 FILLCELL_X2 FILLER_20_95 ();
 FILLCELL_X2 FILLER_20_107 ();
 FILLCELL_X16 FILLER_20_116 ();
 FILLCELL_X8 FILLER_20_132 ();
 FILLCELL_X4 FILLER_20_140 ();
 FILLCELL_X2 FILLER_20_144 ();
 FILLCELL_X1 FILLER_20_146 ();
 FILLCELL_X2 FILLER_20_164 ();
 FILLCELL_X1 FILLER_20_166 ();
 FILLCELL_X8 FILLER_20_178 ();
 FILLCELL_X2 FILLER_20_186 ();
 FILLCELL_X1 FILLER_20_188 ();
 FILLCELL_X4 FILLER_20_213 ();
 FILLCELL_X2 FILLER_20_217 ();
 FILLCELL_X1 FILLER_20_219 ();
 FILLCELL_X2 FILLER_20_227 ();
 FILLCELL_X1 FILLER_20_236 ();
 FILLCELL_X16 FILLER_20_240 ();
 FILLCELL_X2 FILLER_20_263 ();
 FILLCELL_X1 FILLER_20_265 ();
 FILLCELL_X2 FILLER_20_283 ();
 FILLCELL_X1 FILLER_20_285 ();
 FILLCELL_X32 FILLER_20_291 ();
 FILLCELL_X16 FILLER_20_323 ();
 FILLCELL_X4 FILLER_20_339 ();
 FILLCELL_X2 FILLER_20_343 ();
 FILLCELL_X1 FILLER_20_345 ();
 FILLCELL_X4 FILLER_20_360 ();
 FILLCELL_X8 FILLER_20_391 ();
 FILLCELL_X8 FILLER_20_420 ();
 FILLCELL_X1 FILLER_20_435 ();
 FILLCELL_X1 FILLER_20_491 ();
 FILLCELL_X4 FILLER_20_499 ();
 FILLCELL_X2 FILLER_20_503 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X8 FILLER_21_65 ();
 FILLCELL_X2 FILLER_21_73 ();
 FILLCELL_X1 FILLER_21_75 ();
 FILLCELL_X16 FILLER_21_93 ();
 FILLCELL_X8 FILLER_21_126 ();
 FILLCELL_X4 FILLER_21_134 ();
 FILLCELL_X2 FILLER_21_138 ();
 FILLCELL_X1 FILLER_21_147 ();
 FILLCELL_X8 FILLER_21_155 ();
 FILLCELL_X4 FILLER_21_163 ();
 FILLCELL_X16 FILLER_21_206 ();
 FILLCELL_X2 FILLER_21_222 ();
 FILLCELL_X1 FILLER_21_224 ();
 FILLCELL_X8 FILLER_21_242 ();
 FILLCELL_X2 FILLER_21_250 ();
 FILLCELL_X1 FILLER_21_252 ();
 FILLCELL_X4 FILLER_21_275 ();
 FILLCELL_X1 FILLER_21_279 ();
 FILLCELL_X4 FILLER_21_297 ();
 FILLCELL_X1 FILLER_21_301 ();
 FILLCELL_X1 FILLER_21_306 ();
 FILLCELL_X16 FILLER_21_324 ();
 FILLCELL_X4 FILLER_21_340 ();
 FILLCELL_X1 FILLER_21_344 ();
 FILLCELL_X4 FILLER_21_352 ();
 FILLCELL_X2 FILLER_21_356 ();
 FILLCELL_X1 FILLER_21_358 ();
 FILLCELL_X2 FILLER_21_381 ();
 FILLCELL_X2 FILLER_21_388 ();
 FILLCELL_X8 FILLER_21_407 ();
 FILLCELL_X2 FILLER_21_415 ();
 FILLCELL_X2 FILLER_21_424 ();
 FILLCELL_X1 FILLER_21_433 ();
 FILLCELL_X16 FILLER_21_451 ();
 FILLCELL_X2 FILLER_21_467 ();
 FILLCELL_X1 FILLER_21_469 ();
 FILLCELL_X2 FILLER_21_477 ();
 FILLCELL_X2 FILLER_21_484 ();
 FILLCELL_X8 FILLER_21_493 ();
 FILLCELL_X4 FILLER_21_501 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_9 ();
 FILLCELL_X4 FILLER_22_20 ();
 FILLCELL_X1 FILLER_22_24 ();
 FILLCELL_X8 FILLER_22_32 ();
 FILLCELL_X4 FILLER_22_47 ();
 FILLCELL_X2 FILLER_22_51 ();
 FILLCELL_X1 FILLER_22_53 ();
 FILLCELL_X16 FILLER_22_88 ();
 FILLCELL_X2 FILLER_22_104 ();
 FILLCELL_X1 FILLER_22_106 ();
 FILLCELL_X1 FILLER_22_124 ();
 FILLCELL_X1 FILLER_22_152 ();
 FILLCELL_X16 FILLER_22_170 ();
 FILLCELL_X8 FILLER_22_186 ();
 FILLCELL_X2 FILLER_22_194 ();
 FILLCELL_X2 FILLER_22_213 ();
 FILLCELL_X8 FILLER_22_248 ();
 FILLCELL_X4 FILLER_22_256 ();
 FILLCELL_X2 FILLER_22_260 ();
 FILLCELL_X8 FILLER_22_267 ();
 FILLCELL_X4 FILLER_22_299 ();
 FILLCELL_X4 FILLER_22_310 ();
 FILLCELL_X2 FILLER_22_314 ();
 FILLCELL_X4 FILLER_22_323 ();
 FILLCELL_X2 FILLER_22_327 ();
 FILLCELL_X1 FILLER_22_329 ();
 FILLCELL_X2 FILLER_22_347 ();
 FILLCELL_X1 FILLER_22_356 ();
 FILLCELL_X1 FILLER_22_388 ();
 FILLCELL_X2 FILLER_22_396 ();
 FILLCELL_X1 FILLER_22_398 ();
 FILLCELL_X2 FILLER_22_406 ();
 FILLCELL_X1 FILLER_22_408 ();
 FILLCELL_X4 FILLER_22_440 ();
 FILLCELL_X2 FILLER_22_468 ();
 FILLCELL_X1 FILLER_22_470 ();
 FILLCELL_X4 FILLER_22_474 ();
 FILLCELL_X2 FILLER_22_478 ();
 FILLCELL_X16 FILLER_22_483 ();
 FILLCELL_X4 FILLER_22_499 ();
 FILLCELL_X2 FILLER_22_503 ();
 FILLCELL_X1 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_19 ();
 FILLCELL_X1 FILLER_23_37 ();
 FILLCELL_X1 FILLER_23_55 ();
 FILLCELL_X16 FILLER_23_94 ();
 FILLCELL_X4 FILLER_23_110 ();
 FILLCELL_X2 FILLER_23_114 ();
 FILLCELL_X1 FILLER_23_116 ();
 FILLCELL_X1 FILLER_23_131 ();
 FILLCELL_X1 FILLER_23_163 ();
 FILLCELL_X1 FILLER_23_171 ();
 FILLCELL_X2 FILLER_23_179 ();
 FILLCELL_X16 FILLER_23_198 ();
 FILLCELL_X8 FILLER_23_214 ();
 FILLCELL_X2 FILLER_23_222 ();
 FILLCELL_X1 FILLER_23_224 ();
 FILLCELL_X16 FILLER_23_230 ();
 FILLCELL_X1 FILLER_23_246 ();
 FILLCELL_X4 FILLER_23_254 ();
 FILLCELL_X1 FILLER_23_258 ();
 FILLCELL_X4 FILLER_23_271 ();
 FILLCELL_X2 FILLER_23_275 ();
 FILLCELL_X1 FILLER_23_277 ();
 FILLCELL_X4 FILLER_23_295 ();
 FILLCELL_X8 FILLER_23_323 ();
 FILLCELL_X1 FILLER_23_331 ();
 FILLCELL_X1 FILLER_23_363 ();
 FILLCELL_X16 FILLER_23_371 ();
 FILLCELL_X1 FILLER_23_407 ();
 FILLCELL_X16 FILLER_23_411 ();
 FILLCELL_X8 FILLER_23_427 ();
 FILLCELL_X4 FILLER_23_435 ();
 FILLCELL_X2 FILLER_23_439 ();
 FILLCELL_X1 FILLER_23_441 ();
 FILLCELL_X8 FILLER_23_497 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X4 FILLER_24_9 ();
 FILLCELL_X2 FILLER_24_13 ();
 FILLCELL_X8 FILLER_24_22 ();
 FILLCELL_X1 FILLER_24_37 ();
 FILLCELL_X4 FILLER_24_45 ();
 FILLCELL_X1 FILLER_24_49 ();
 FILLCELL_X4 FILLER_24_57 ();
 FILLCELL_X2 FILLER_24_75 ();
 FILLCELL_X2 FILLER_24_84 ();
 FILLCELL_X8 FILLER_24_89 ();
 FILLCELL_X8 FILLER_24_121 ();
 FILLCELL_X4 FILLER_24_129 ();
 FILLCELL_X16 FILLER_24_141 ();
 FILLCELL_X1 FILLER_24_157 ();
 FILLCELL_X8 FILLER_24_164 ();
 FILLCELL_X4 FILLER_24_172 ();
 FILLCELL_X1 FILLER_24_176 ();
 FILLCELL_X2 FILLER_24_183 ();
 FILLCELL_X4 FILLER_24_199 ();
 FILLCELL_X2 FILLER_24_203 ();
 FILLCELL_X8 FILLER_24_212 ();
 FILLCELL_X2 FILLER_24_220 ();
 FILLCELL_X8 FILLER_24_239 ();
 FILLCELL_X1 FILLER_24_247 ();
 FILLCELL_X4 FILLER_24_265 ();
 FILLCELL_X1 FILLER_24_269 ();
 FILLCELL_X4 FILLER_24_273 ();
 FILLCELL_X1 FILLER_24_277 ();
 FILLCELL_X4 FILLER_24_288 ();
 FILLCELL_X4 FILLER_24_299 ();
 FILLCELL_X2 FILLER_24_303 ();
 FILLCELL_X8 FILLER_24_312 ();
 FILLCELL_X2 FILLER_24_320 ();
 FILLCELL_X16 FILLER_24_325 ();
 FILLCELL_X8 FILLER_24_341 ();
 FILLCELL_X4 FILLER_24_349 ();
 FILLCELL_X1 FILLER_24_353 ();
 FILLCELL_X2 FILLER_24_371 ();
 FILLCELL_X1 FILLER_24_373 ();
 FILLCELL_X8 FILLER_24_384 ();
 FILLCELL_X1 FILLER_24_392 ();
 FILLCELL_X4 FILLER_24_398 ();
 FILLCELL_X2 FILLER_24_402 ();
 FILLCELL_X32 FILLER_24_411 ();
 FILLCELL_X16 FILLER_24_443 ();
 FILLCELL_X8 FILLER_24_459 ();
 FILLCELL_X2 FILLER_24_467 ();
 FILLCELL_X1 FILLER_24_504 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_9 ();
 FILLCELL_X32 FILLER_25_40 ();
 FILLCELL_X4 FILLER_25_72 ();
 FILLCELL_X2 FILLER_25_76 ();
 FILLCELL_X2 FILLER_25_90 ();
 FILLCELL_X8 FILLER_25_98 ();
 FILLCELL_X4 FILLER_25_123 ();
 FILLCELL_X2 FILLER_25_127 ();
 FILLCELL_X1 FILLER_25_129 ();
 FILLCELL_X2 FILLER_25_133 ();
 FILLCELL_X16 FILLER_25_162 ();
 FILLCELL_X8 FILLER_25_195 ();
 FILLCELL_X4 FILLER_25_220 ();
 FILLCELL_X1 FILLER_25_224 ();
 FILLCELL_X2 FILLER_25_232 ();
 FILLCELL_X8 FILLER_25_237 ();
 FILLCELL_X1 FILLER_25_245 ();
 FILLCELL_X2 FILLER_25_249 ();
 FILLCELL_X8 FILLER_25_256 ();
 FILLCELL_X4 FILLER_25_264 ();
 FILLCELL_X1 FILLER_25_324 ();
 FILLCELL_X32 FILLER_25_332 ();
 FILLCELL_X4 FILLER_25_364 ();
 FILLCELL_X2 FILLER_25_399 ();
 FILLCELL_X1 FILLER_25_401 ();
 FILLCELL_X2 FILLER_25_412 ();
 FILLCELL_X8 FILLER_25_421 ();
 FILLCELL_X2 FILLER_25_429 ();
 FILLCELL_X8 FILLER_25_438 ();
 FILLCELL_X2 FILLER_25_446 ();
 FILLCELL_X4 FILLER_25_465 ();
 FILLCELL_X1 FILLER_25_469 ();
 FILLCELL_X4 FILLER_25_473 ();
 FILLCELL_X2 FILLER_25_477 ();
 FILLCELL_X16 FILLER_25_482 ();
 FILLCELL_X4 FILLER_25_498 ();
 FILLCELL_X2 FILLER_25_502 ();
 FILLCELL_X1 FILLER_25_504 ();
 FILLCELL_X2 FILLER_26_1 ();
 FILLCELL_X8 FILLER_26_44 ();
 FILLCELL_X2 FILLER_26_76 ();
 FILLCELL_X2 FILLER_26_91 ();
 FILLCELL_X1 FILLER_26_93 ();
 FILLCELL_X8 FILLER_26_97 ();
 FILLCELL_X2 FILLER_26_105 ();
 FILLCELL_X1 FILLER_26_107 ();
 FILLCELL_X4 FILLER_26_125 ();
 FILLCELL_X1 FILLER_26_136 ();
 FILLCELL_X2 FILLER_26_144 ();
 FILLCELL_X4 FILLER_26_153 ();
 FILLCELL_X1 FILLER_26_157 ();
 FILLCELL_X2 FILLER_26_172 ();
 FILLCELL_X2 FILLER_26_195 ();
 FILLCELL_X1 FILLER_26_197 ();
 FILLCELL_X8 FILLER_26_215 ();
 FILLCELL_X1 FILLER_26_230 ();
 FILLCELL_X1 FILLER_26_238 ();
 FILLCELL_X2 FILLER_26_273 ();
 FILLCELL_X4 FILLER_26_299 ();
 FILLCELL_X2 FILLER_26_303 ();
 FILLCELL_X4 FILLER_26_319 ();
 FILLCELL_X2 FILLER_26_323 ();
 FILLCELL_X1 FILLER_26_325 ();
 FILLCELL_X16 FILLER_26_350 ();
 FILLCELL_X8 FILLER_26_366 ();
 FILLCELL_X8 FILLER_26_381 ();
 FILLCELL_X4 FILLER_26_389 ();
 FILLCELL_X1 FILLER_26_393 ();
 FILLCELL_X8 FILLER_26_406 ();
 FILLCELL_X2 FILLER_26_462 ();
 FILLCELL_X1 FILLER_26_464 ();
 FILLCELL_X2 FILLER_26_479 ();
 FILLCELL_X2 FILLER_26_484 ();
 FILLCELL_X2 FILLER_26_503 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_5 ();
 FILLCELL_X4 FILLER_27_24 ();
 FILLCELL_X2 FILLER_27_28 ();
 FILLCELL_X4 FILLER_27_54 ();
 FILLCELL_X1 FILLER_27_58 ();
 FILLCELL_X4 FILLER_27_66 ();
 FILLCELL_X1 FILLER_27_70 ();
 FILLCELL_X1 FILLER_27_78 ();
 FILLCELL_X1 FILLER_27_82 ();
 FILLCELL_X16 FILLER_27_104 ();
 FILLCELL_X8 FILLER_27_120 ();
 FILLCELL_X2 FILLER_27_128 ();
 FILLCELL_X8 FILLER_27_184 ();
 FILLCELL_X1 FILLER_27_192 ();
 FILLCELL_X8 FILLER_27_196 ();
 FILLCELL_X2 FILLER_27_204 ();
 FILLCELL_X4 FILLER_27_223 ();
 FILLCELL_X2 FILLER_27_227 ();
 FILLCELL_X1 FILLER_27_229 ();
 FILLCELL_X16 FILLER_27_233 ();
 FILLCELL_X8 FILLER_27_266 ();
 FILLCELL_X1 FILLER_27_274 ();
 FILLCELL_X1 FILLER_27_282 ();
 FILLCELL_X8 FILLER_27_288 ();
 FILLCELL_X4 FILLER_27_299 ();
 FILLCELL_X1 FILLER_27_320 ();
 FILLCELL_X4 FILLER_27_324 ();
 FILLCELL_X4 FILLER_27_335 ();
 FILLCELL_X2 FILLER_27_339 ();
 FILLCELL_X4 FILLER_27_348 ();
 FILLCELL_X4 FILLER_27_362 ();
 FILLCELL_X4 FILLER_27_390 ();
 FILLCELL_X2 FILLER_27_411 ();
 FILLCELL_X1 FILLER_27_413 ();
 FILLCELL_X4 FILLER_27_421 ();
 FILLCELL_X1 FILLER_27_425 ();
 FILLCELL_X8 FILLER_27_433 ();
 FILLCELL_X4 FILLER_27_441 ();
 FILLCELL_X2 FILLER_27_445 ();
 FILLCELL_X4 FILLER_27_450 ();
 FILLCELL_X1 FILLER_27_454 ();
 FILLCELL_X2 FILLER_27_472 ();
 FILLCELL_X2 FILLER_27_481 ();
 FILLCELL_X1 FILLER_27_483 ();
 FILLCELL_X8 FILLER_27_491 ();
 FILLCELL_X4 FILLER_27_499 ();
 FILLCELL_X2 FILLER_27_503 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_17 ();
 FILLCELL_X8 FILLER_28_49 ();
 FILLCELL_X2 FILLER_28_57 ();
 FILLCELL_X1 FILLER_28_76 ();
 FILLCELL_X2 FILLER_28_80 ();
 FILLCELL_X2 FILLER_28_89 ();
 FILLCELL_X2 FILLER_28_108 ();
 FILLCELL_X16 FILLER_28_127 ();
 FILLCELL_X8 FILLER_28_143 ();
 FILLCELL_X2 FILLER_28_151 ();
 FILLCELL_X1 FILLER_28_153 ();
 FILLCELL_X16 FILLER_28_181 ();
 FILLCELL_X2 FILLER_28_197 ();
 FILLCELL_X4 FILLER_28_209 ();
 FILLCELL_X2 FILLER_28_213 ();
 FILLCELL_X16 FILLER_28_229 ();
 FILLCELL_X2 FILLER_28_245 ();
 FILLCELL_X1 FILLER_28_247 ();
 FILLCELL_X2 FILLER_28_255 ();
 FILLCELL_X16 FILLER_28_264 ();
 FILLCELL_X8 FILLER_28_280 ();
 FILLCELL_X16 FILLER_28_295 ();
 FILLCELL_X4 FILLER_28_311 ();
 FILLCELL_X1 FILLER_28_315 ();
 FILLCELL_X4 FILLER_28_323 ();
 FILLCELL_X2 FILLER_28_327 ();
 FILLCELL_X1 FILLER_28_329 ();
 FILLCELL_X2 FILLER_28_347 ();
 FILLCELL_X1 FILLER_28_349 ();
 FILLCELL_X16 FILLER_28_374 ();
 FILLCELL_X4 FILLER_28_390 ();
 FILLCELL_X4 FILLER_28_411 ();
 FILLCELL_X4 FILLER_28_432 ();
 FILLCELL_X2 FILLER_28_436 ();
 FILLCELL_X4 FILLER_28_442 ();
 FILLCELL_X2 FILLER_28_446 ();
 FILLCELL_X2 FILLER_28_452 ();
 FILLCELL_X1 FILLER_28_454 ();
 FILLCELL_X16 FILLER_28_459 ();
 FILLCELL_X2 FILLER_28_475 ();
 FILLCELL_X4 FILLER_28_501 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_9 ();
 FILLCELL_X2 FILLER_29_13 ();
 FILLCELL_X1 FILLER_29_15 ();
 FILLCELL_X32 FILLER_29_40 ();
 FILLCELL_X8 FILLER_29_72 ();
 FILLCELL_X4 FILLER_29_80 ();
 FILLCELL_X1 FILLER_29_84 ();
 FILLCELL_X2 FILLER_29_102 ();
 FILLCELL_X1 FILLER_29_104 ();
 FILLCELL_X4 FILLER_29_119 ();
 FILLCELL_X2 FILLER_29_123 ();
 FILLCELL_X8 FILLER_29_132 ();
 FILLCELL_X1 FILLER_29_147 ();
 FILLCELL_X1 FILLER_29_165 ();
 FILLCELL_X8 FILLER_29_174 ();
 FILLCELL_X4 FILLER_29_182 ();
 FILLCELL_X1 FILLER_29_193 ();
 FILLCELL_X1 FILLER_29_197 ();
 FILLCELL_X8 FILLER_29_201 ();
 FILLCELL_X4 FILLER_29_209 ();
 FILLCELL_X1 FILLER_29_213 ();
 FILLCELL_X16 FILLER_29_265 ();
 FILLCELL_X4 FILLER_29_281 ();
 FILLCELL_X1 FILLER_29_285 ();
 FILLCELL_X2 FILLER_29_291 ();
 FILLCELL_X1 FILLER_29_293 ();
 FILLCELL_X2 FILLER_29_301 ();
 FILLCELL_X1 FILLER_29_303 ();
 FILLCELL_X1 FILLER_29_328 ();
 FILLCELL_X2 FILLER_29_358 ();
 FILLCELL_X2 FILLER_29_367 ();
 FILLCELL_X1 FILLER_29_369 ();
 FILLCELL_X4 FILLER_29_373 ();
 FILLCELL_X1 FILLER_29_377 ();
 FILLCELL_X16 FILLER_29_402 ();
 FILLCELL_X2 FILLER_29_418 ();
 FILLCELL_X1 FILLER_29_451 ();
 FILLCELL_X8 FILLER_29_469 ();
 FILLCELL_X2 FILLER_29_502 ();
 FILLCELL_X1 FILLER_29_504 ();
 FILLCELL_X16 FILLER_30_1 ();
 FILLCELL_X8 FILLER_30_17 ();
 FILLCELL_X2 FILLER_30_25 ();
 FILLCELL_X1 FILLER_30_27 ();
 FILLCELL_X8 FILLER_30_42 ();
 FILLCELL_X4 FILLER_30_50 ();
 FILLCELL_X1 FILLER_30_54 ();
 FILLCELL_X1 FILLER_30_82 ();
 FILLCELL_X8 FILLER_30_90 ();
 FILLCELL_X4 FILLER_30_98 ();
 FILLCELL_X2 FILLER_30_102 ();
 FILLCELL_X1 FILLER_30_104 ();
 FILLCELL_X2 FILLER_30_112 ();
 FILLCELL_X1 FILLER_30_114 ();
 FILLCELL_X1 FILLER_30_149 ();
 FILLCELL_X8 FILLER_30_167 ();
 FILLCELL_X2 FILLER_30_175 ();
 FILLCELL_X1 FILLER_30_177 ();
 FILLCELL_X1 FILLER_30_205 ();
 FILLCELL_X16 FILLER_30_213 ();
 FILLCELL_X4 FILLER_30_229 ();
 FILLCELL_X2 FILLER_30_233 ();
 FILLCELL_X1 FILLER_30_235 ();
 FILLCELL_X2 FILLER_30_265 ();
 FILLCELL_X8 FILLER_30_284 ();
 FILLCELL_X8 FILLER_30_316 ();
 FILLCELL_X1 FILLER_30_341 ();
 FILLCELL_X8 FILLER_30_373 ();
 FILLCELL_X2 FILLER_30_381 ();
 FILLCELL_X8 FILLER_30_397 ();
 FILLCELL_X4 FILLER_30_405 ();
 FILLCELL_X2 FILLER_30_409 ();
 FILLCELL_X1 FILLER_30_411 ();
 FILLCELL_X1 FILLER_30_415 ();
 FILLCELL_X2 FILLER_30_440 ();
 FILLCELL_X1 FILLER_30_442 ();
 FILLCELL_X2 FILLER_30_467 ();
 FILLCELL_X1 FILLER_30_469 ();
 FILLCELL_X4 FILLER_30_484 ();
 FILLCELL_X2 FILLER_30_488 ();
 FILLCELL_X8 FILLER_30_497 ();
 FILLCELL_X8 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_9 ();
 FILLCELL_X1 FILLER_31_11 ();
 FILLCELL_X2 FILLER_31_19 ();
 FILLCELL_X8 FILLER_31_38 ();
 FILLCELL_X2 FILLER_31_46 ();
 FILLCELL_X1 FILLER_31_48 ();
 FILLCELL_X1 FILLER_31_80 ();
 FILLCELL_X8 FILLER_31_84 ();
 FILLCELL_X4 FILLER_31_92 ();
 FILLCELL_X2 FILLER_31_105 ();
 FILLCELL_X1 FILLER_31_107 ();
 FILLCELL_X8 FILLER_31_111 ();
 FILLCELL_X4 FILLER_31_119 ();
 FILLCELL_X1 FILLER_31_123 ();
 FILLCELL_X16 FILLER_31_131 ();
 FILLCELL_X8 FILLER_31_147 ();
 FILLCELL_X4 FILLER_31_155 ();
 FILLCELL_X2 FILLER_31_159 ();
 FILLCELL_X4 FILLER_31_168 ();
 FILLCELL_X2 FILLER_31_172 ();
 FILLCELL_X1 FILLER_31_174 ();
 FILLCELL_X2 FILLER_31_199 ();
 FILLCELL_X1 FILLER_31_208 ();
 FILLCELL_X2 FILLER_31_233 ();
 FILLCELL_X2 FILLER_31_242 ();
 FILLCELL_X8 FILLER_31_254 ();
 FILLCELL_X2 FILLER_31_262 ();
 FILLCELL_X8 FILLER_31_288 ();
 FILLCELL_X1 FILLER_31_296 ();
 FILLCELL_X2 FILLER_31_314 ();
 FILLCELL_X1 FILLER_31_316 ();
 FILLCELL_X16 FILLER_31_320 ();
 FILLCELL_X8 FILLER_31_336 ();
 FILLCELL_X1 FILLER_31_357 ();
 FILLCELL_X1 FILLER_31_365 ();
 FILLCELL_X16 FILLER_31_369 ();
 FILLCELL_X4 FILLER_31_385 ();
 FILLCELL_X2 FILLER_31_389 ();
 FILLCELL_X2 FILLER_31_401 ();
 FILLCELL_X8 FILLER_31_413 ();
 FILLCELL_X2 FILLER_31_421 ();
 FILLCELL_X4 FILLER_31_430 ();
 FILLCELL_X8 FILLER_31_439 ();
 FILLCELL_X4 FILLER_31_461 ();
 FILLCELL_X2 FILLER_31_465 ();
 FILLCELL_X1 FILLER_31_467 ();
 FILLCELL_X4 FILLER_31_471 ();
 FILLCELL_X1 FILLER_31_478 ();
 FILLCELL_X4 FILLER_31_496 ();
 FILLCELL_X1 FILLER_31_504 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X4 FILLER_32_27 ();
 FILLCELL_X1 FILLER_32_31 ();
 FILLCELL_X1 FILLER_32_46 ();
 FILLCELL_X8 FILLER_32_71 ();
 FILLCELL_X2 FILLER_32_89 ();
 FILLCELL_X8 FILLER_32_120 ();
 FILLCELL_X2 FILLER_32_128 ();
 FILLCELL_X32 FILLER_32_139 ();
 FILLCELL_X4 FILLER_32_171 ();
 FILLCELL_X2 FILLER_32_175 ();
 FILLCELL_X1 FILLER_32_177 ();
 FILLCELL_X1 FILLER_32_181 ();
 FILLCELL_X2 FILLER_32_206 ();
 FILLCELL_X1 FILLER_32_208 ();
 FILLCELL_X16 FILLER_32_216 ();
 FILLCELL_X4 FILLER_32_232 ();
 FILLCELL_X2 FILLER_32_236 ();
 FILLCELL_X2 FILLER_32_262 ();
 FILLCELL_X4 FILLER_32_283 ();
 FILLCELL_X4 FILLER_32_297 ();
 FILLCELL_X4 FILLER_32_306 ();
 FILLCELL_X1 FILLER_32_310 ();
 FILLCELL_X16 FILLER_32_325 ();
 FILLCELL_X4 FILLER_32_341 ();
 FILLCELL_X1 FILLER_32_345 ();
 FILLCELL_X4 FILLER_32_370 ();
 FILLCELL_X1 FILLER_32_374 ();
 FILLCELL_X8 FILLER_32_382 ();
 FILLCELL_X4 FILLER_32_414 ();
 FILLCELL_X2 FILLER_32_418 ();
 FILLCELL_X1 FILLER_32_420 ();
 FILLCELL_X32 FILLER_32_438 ();
 FILLCELL_X32 FILLER_32_470 ();
 FILLCELL_X2 FILLER_32_502 ();
 FILLCELL_X1 FILLER_32_504 ();
 FILLCELL_X8 FILLER_33_1 ();
 FILLCELL_X4 FILLER_33_9 ();
 FILLCELL_X2 FILLER_33_13 ();
 FILLCELL_X1 FILLER_33_15 ();
 FILLCELL_X16 FILLER_33_40 ();
 FILLCELL_X4 FILLER_33_56 ();
 FILLCELL_X2 FILLER_33_67 ();
 FILLCELL_X2 FILLER_33_76 ();
 FILLCELL_X1 FILLER_33_78 ();
 FILLCELL_X4 FILLER_33_82 ();
 FILLCELL_X2 FILLER_33_86 ();
 FILLCELL_X1 FILLER_33_97 ();
 FILLCELL_X1 FILLER_33_110 ();
 FILLCELL_X2 FILLER_33_144 ();
 FILLCELL_X4 FILLER_33_149 ();
 FILLCELL_X4 FILLER_33_198 ();
 FILLCELL_X1 FILLER_33_202 ();
 FILLCELL_X4 FILLER_33_210 ();
 FILLCELL_X8 FILLER_33_234 ();
 FILLCELL_X4 FILLER_33_242 ();
 FILLCELL_X2 FILLER_33_253 ();
 FILLCELL_X1 FILLER_33_269 ();
 FILLCELL_X4 FILLER_33_277 ();
 FILLCELL_X1 FILLER_33_281 ();
 FILLCELL_X4 FILLER_33_292 ();
 FILLCELL_X2 FILLER_33_296 ();
 FILLCELL_X1 FILLER_33_298 ();
 FILLCELL_X2 FILLER_33_313 ();
 FILLCELL_X1 FILLER_33_315 ();
 FILLCELL_X4 FILLER_33_319 ();
 FILLCELL_X1 FILLER_33_323 ();
 FILLCELL_X8 FILLER_33_331 ();
 FILLCELL_X1 FILLER_33_339 ();
 FILLCELL_X16 FILLER_33_347 ();
 FILLCELL_X2 FILLER_33_363 ();
 FILLCELL_X16 FILLER_33_399 ();
 FILLCELL_X4 FILLER_33_415 ();
 FILLCELL_X16 FILLER_33_426 ();
 FILLCELL_X8 FILLER_33_460 ();
 FILLCELL_X4 FILLER_33_468 ();
 FILLCELL_X2 FILLER_33_472 ();
 FILLCELL_X1 FILLER_33_474 ();
 FILLCELL_X1 FILLER_33_481 ();
 FILLCELL_X8 FILLER_34_1 ();
 FILLCELL_X2 FILLER_34_9 ();
 FILLCELL_X32 FILLER_34_25 ();
 FILLCELL_X2 FILLER_34_57 ();
 FILLCELL_X4 FILLER_34_76 ();
 FILLCELL_X1 FILLER_34_80 ();
 FILLCELL_X1 FILLER_34_104 ();
 FILLCELL_X1 FILLER_34_114 ();
 FILLCELL_X2 FILLER_34_118 ();
 FILLCELL_X2 FILLER_34_126 ();
 FILLCELL_X2 FILLER_34_134 ();
 FILLCELL_X2 FILLER_34_187 ();
 FILLCELL_X2 FILLER_34_202 ();
 FILLCELL_X1 FILLER_34_204 ();
 FILLCELL_X4 FILLER_34_238 ();
 FILLCELL_X2 FILLER_34_242 ();
 FILLCELL_X4 FILLER_34_251 ();
 FILLCELL_X1 FILLER_34_260 ();
 FILLCELL_X8 FILLER_34_278 ();
 FILLCELL_X4 FILLER_34_286 ();
 FILLCELL_X2 FILLER_34_290 ();
 FILLCELL_X1 FILLER_34_292 ();
 FILLCELL_X1 FILLER_34_317 ();
 FILLCELL_X2 FILLER_34_325 ();
 FILLCELL_X1 FILLER_34_351 ();
 FILLCELL_X8 FILLER_34_373 ();
 FILLCELL_X4 FILLER_34_381 ();
 FILLCELL_X8 FILLER_34_402 ();
 FILLCELL_X4 FILLER_34_410 ();
 FILLCELL_X2 FILLER_34_414 ();
 FILLCELL_X8 FILLER_34_433 ();
 FILLCELL_X2 FILLER_34_441 ();
 FILLCELL_X1 FILLER_34_443 ();
 FILLCELL_X2 FILLER_34_464 ();
 FILLCELL_X2 FILLER_34_495 ();
 FILLCELL_X1 FILLER_34_497 ();
 FILLCELL_X1 FILLER_34_504 ();
 FILLCELL_X4 FILLER_35_1 ();
 FILLCELL_X8 FILLER_35_22 ();
 FILLCELL_X2 FILLER_35_30 ();
 FILLCELL_X16 FILLER_35_59 ();
 FILLCELL_X4 FILLER_35_115 ();
 FILLCELL_X1 FILLER_35_136 ();
 FILLCELL_X16 FILLER_35_143 ();
 FILLCELL_X4 FILLER_35_162 ();
 FILLCELL_X2 FILLER_35_166 ();
 FILLCELL_X1 FILLER_35_191 ();
 FILLCELL_X1 FILLER_35_239 ();
 FILLCELL_X8 FILLER_35_254 ();
 FILLCELL_X2 FILLER_35_262 ();
 FILLCELL_X1 FILLER_35_271 ();
 FILLCELL_X2 FILLER_35_296 ();
 FILLCELL_X4 FILLER_35_322 ();
 FILLCELL_X2 FILLER_35_326 ();
 FILLCELL_X1 FILLER_35_328 ();
 FILLCELL_X4 FILLER_35_357 ();
 FILLCELL_X32 FILLER_35_367 ();
 FILLCELL_X2 FILLER_35_399 ();
 FILLCELL_X1 FILLER_35_431 ();
 FILLCELL_X16 FILLER_35_446 ();
 FILLCELL_X1 FILLER_35_471 ();
 FILLCELL_X1 FILLER_35_486 ();
 FILLCELL_X1 FILLER_35_490 ();
 FILLCELL_X1 FILLER_36_4 ();
 FILLCELL_X2 FILLER_36_39 ();
 FILLCELL_X4 FILLER_36_58 ();
 FILLCELL_X8 FILLER_36_79 ();
 FILLCELL_X4 FILLER_36_87 ();
 FILLCELL_X2 FILLER_36_104 ();
 FILLCELL_X32 FILLER_36_118 ();
 FILLCELL_X16 FILLER_36_150 ();
 FILLCELL_X4 FILLER_36_166 ();
 FILLCELL_X2 FILLER_36_170 ();
 FILLCELL_X1 FILLER_36_265 ();
 FILLCELL_X1 FILLER_36_278 ();
 FILLCELL_X8 FILLER_36_303 ();
 FILLCELL_X1 FILLER_36_311 ();
 FILLCELL_X8 FILLER_36_326 ();
 FILLCELL_X1 FILLER_36_334 ();
 FILLCELL_X2 FILLER_36_354 ();
 FILLCELL_X1 FILLER_36_356 ();
 FILLCELL_X16 FILLER_36_365 ();
 FILLCELL_X8 FILLER_36_405 ();
 FILLCELL_X16 FILLER_36_447 ();
 FILLCELL_X2 FILLER_36_463 ();
 FILLCELL_X1 FILLER_36_465 ();
 FILLCELL_X4 FILLER_36_477 ();
 FILLCELL_X2 FILLER_36_481 ();
 FILLCELL_X1 FILLER_36_483 ();
 FILLCELL_X8 FILLER_36_488 ();
 FILLCELL_X8 FILLER_37_1 ();
 FILLCELL_X2 FILLER_37_9 ();
 FILLCELL_X1 FILLER_37_11 ();
 FILLCELL_X2 FILLER_37_26 ();
 FILLCELL_X1 FILLER_37_28 ();
 FILLCELL_X2 FILLER_37_36 ();
 FILLCELL_X1 FILLER_37_38 ();
 FILLCELL_X4 FILLER_37_46 ();
 FILLCELL_X1 FILLER_37_50 ();
 FILLCELL_X4 FILLER_37_54 ();
 FILLCELL_X1 FILLER_37_58 ();
 FILLCELL_X2 FILLER_37_84 ();
 FILLCELL_X4 FILLER_37_121 ();
 FILLCELL_X1 FILLER_37_125 ();
 FILLCELL_X8 FILLER_37_167 ();
 FILLCELL_X1 FILLER_37_175 ();
 FILLCELL_X1 FILLER_37_183 ();
 FILLCELL_X1 FILLER_37_246 ();
 FILLCELL_X4 FILLER_37_264 ();
 FILLCELL_X2 FILLER_37_279 ();
 FILLCELL_X1 FILLER_37_281 ();
 FILLCELL_X8 FILLER_37_299 ();
 FILLCELL_X2 FILLER_37_307 ();
 FILLCELL_X1 FILLER_37_329 ();
 FILLCELL_X8 FILLER_37_349 ();
 FILLCELL_X2 FILLER_37_357 ();
 FILLCELL_X1 FILLER_37_359 ();
 FILLCELL_X8 FILLER_37_367 ();
 FILLCELL_X4 FILLER_37_375 ();
 FILLCELL_X2 FILLER_37_379 ();
 FILLCELL_X1 FILLER_37_381 ();
 FILLCELL_X8 FILLER_37_389 ();
 FILLCELL_X2 FILLER_37_397 ();
 FILLCELL_X1 FILLER_37_406 ();
 FILLCELL_X1 FILLER_37_424 ();
 FILLCELL_X1 FILLER_37_437 ();
 FILLCELL_X8 FILLER_37_449 ();
 FILLCELL_X4 FILLER_37_457 ();
 FILLCELL_X1 FILLER_37_461 ();
 FILLCELL_X4 FILLER_37_466 ();
 FILLCELL_X1 FILLER_37_470 ();
 FILLCELL_X2 FILLER_37_486 ();
 FILLCELL_X1 FILLER_37_498 ();
 FILLCELL_X8 FILLER_38_1 ();
 FILLCELL_X4 FILLER_38_9 ();
 FILLCELL_X1 FILLER_38_13 ();
 FILLCELL_X8 FILLER_38_17 ();
 FILLCELL_X4 FILLER_38_25 ();
 FILLCELL_X1 FILLER_38_29 ();
 FILLCELL_X16 FILLER_38_34 ();
 FILLCELL_X4 FILLER_38_50 ();
 FILLCELL_X4 FILLER_38_61 ();
 FILLCELL_X2 FILLER_38_65 ();
 FILLCELL_X1 FILLER_38_67 ();
 FILLCELL_X4 FILLER_38_92 ();
 FILLCELL_X1 FILLER_38_96 ();
 FILLCELL_X8 FILLER_38_117 ();
 FILLCELL_X4 FILLER_38_125 ();
 FILLCELL_X1 FILLER_38_136 ();
 FILLCELL_X2 FILLER_38_144 ();
 FILLCELL_X4 FILLER_38_162 ();
 FILLCELL_X1 FILLER_38_166 ();
 FILLCELL_X2 FILLER_38_204 ();
 FILLCELL_X1 FILLER_38_291 ();
 FILLCELL_X4 FILLER_38_355 ();
 FILLCELL_X1 FILLER_38_359 ();
 FILLCELL_X2 FILLER_38_377 ();
 FILLCELL_X1 FILLER_38_379 ();
 FILLCELL_X4 FILLER_38_404 ();
 FILLCELL_X1 FILLER_38_408 ();
 FILLCELL_X1 FILLER_38_429 ();
 FILLCELL_X8 FILLER_38_433 ();
 FILLCELL_X1 FILLER_38_441 ();
 FILLCELL_X1 FILLER_38_465 ();
 FILLCELL_X1 FILLER_38_483 ();
 FILLCELL_X4 FILLER_38_489 ();
 FILLCELL_X2 FILLER_38_493 ();
 FILLCELL_X4 FILLER_38_498 ();
 FILLCELL_X2 FILLER_38_502 ();
 FILLCELL_X1 FILLER_38_504 ();
 FILLCELL_X2 FILLER_39_1 ();
 FILLCELL_X2 FILLER_39_20 ();
 FILLCELL_X1 FILLER_39_22 ();
 FILLCELL_X2 FILLER_39_30 ();
 FILLCELL_X1 FILLER_39_32 ();
 FILLCELL_X32 FILLER_39_53 ();
 FILLCELL_X16 FILLER_39_85 ();
 FILLCELL_X8 FILLER_39_101 ();
 FILLCELL_X4 FILLER_39_109 ();
 FILLCELL_X1 FILLER_39_113 ();
 FILLCELL_X4 FILLER_39_131 ();
 FILLCELL_X2 FILLER_39_135 ();
 FILLCELL_X1 FILLER_39_137 ();
 FILLCELL_X4 FILLER_39_187 ();
 FILLCELL_X2 FILLER_39_191 ();
 FILLCELL_X1 FILLER_39_193 ();
 FILLCELL_X2 FILLER_39_221 ();
 FILLCELL_X1 FILLER_39_240 ();
 FILLCELL_X4 FILLER_39_262 ();
 FILLCELL_X2 FILLER_39_266 ();
 FILLCELL_X4 FILLER_39_275 ();
 FILLCELL_X2 FILLER_39_279 ();
 FILLCELL_X1 FILLER_39_312 ();
 FILLCELL_X1 FILLER_39_321 ();
 FILLCELL_X2 FILLER_39_336 ();
 FILLCELL_X1 FILLER_39_338 ();
 FILLCELL_X4 FILLER_39_366 ();
 FILLCELL_X2 FILLER_39_370 ();
 FILLCELL_X1 FILLER_39_372 ();
 FILLCELL_X8 FILLER_39_395 ();
 FILLCELL_X2 FILLER_39_403 ();
 FILLCELL_X4 FILLER_39_408 ();
 FILLCELL_X2 FILLER_39_412 ();
 FILLCELL_X1 FILLER_39_414 ();
 FILLCELL_X16 FILLER_39_427 ();
 FILLCELL_X2 FILLER_39_443 ();
 FILLCELL_X1 FILLER_39_445 ();
 FILLCELL_X4 FILLER_39_458 ();
 FILLCELL_X2 FILLER_39_462 ();
 FILLCELL_X1 FILLER_39_464 ();
 FILLCELL_X1 FILLER_39_476 ();
 FILLCELL_X1 FILLER_39_483 ();
 FILLCELL_X1 FILLER_39_488 ();
 FILLCELL_X1 FILLER_39_492 ();
 FILLCELL_X2 FILLER_39_500 ();
 FILLCELL_X8 FILLER_40_1 ();
 FILLCELL_X4 FILLER_40_9 ();
 FILLCELL_X1 FILLER_40_13 ();
 FILLCELL_X2 FILLER_40_21 ();
 FILLCELL_X1 FILLER_40_23 ();
 FILLCELL_X2 FILLER_40_31 ();
 FILLCELL_X1 FILLER_40_43 ();
 FILLCELL_X4 FILLER_40_51 ();
 FILLCELL_X16 FILLER_40_62 ();
 FILLCELL_X2 FILLER_40_78 ();
 FILLCELL_X8 FILLER_40_97 ();
 FILLCELL_X4 FILLER_40_105 ();
 FILLCELL_X2 FILLER_40_109 ();
 FILLCELL_X2 FILLER_40_118 ();
 FILLCELL_X1 FILLER_40_130 ();
 FILLCELL_X1 FILLER_40_138 ();
 FILLCELL_X2 FILLER_40_142 ();
 FILLCELL_X16 FILLER_40_175 ();
 FILLCELL_X4 FILLER_40_191 ();
 FILLCELL_X2 FILLER_40_195 ();
 FILLCELL_X1 FILLER_40_197 ();
 FILLCELL_X1 FILLER_40_229 ();
 FILLCELL_X4 FILLER_40_251 ();
 FILLCELL_X2 FILLER_40_262 ();
 FILLCELL_X1 FILLER_40_264 ();
 FILLCELL_X4 FILLER_40_272 ();
 FILLCELL_X1 FILLER_40_276 ();
 FILLCELL_X2 FILLER_40_284 ();
 FILLCELL_X1 FILLER_40_307 ();
 FILLCELL_X32 FILLER_40_343 ();
 FILLCELL_X2 FILLER_40_375 ();
 FILLCELL_X4 FILLER_40_384 ();
 FILLCELL_X2 FILLER_40_388 ();
 FILLCELL_X16 FILLER_40_407 ();
 FILLCELL_X4 FILLER_40_423 ();
 FILLCELL_X2 FILLER_40_427 ();
 FILLCELL_X1 FILLER_40_429 ();
 FILLCELL_X32 FILLER_40_434 ();
 FILLCELL_X4 FILLER_40_466 ();
 FILLCELL_X1 FILLER_40_470 ();
 FILLCELL_X8 FILLER_40_495 ();
 FILLCELL_X2 FILLER_40_503 ();
 FILLCELL_X16 FILLER_41_1 ();
 FILLCELL_X2 FILLER_41_17 ();
 FILLCELL_X8 FILLER_41_96 ();
 FILLCELL_X1 FILLER_41_104 ();
 FILLCELL_X4 FILLER_41_116 ();
 FILLCELL_X2 FILLER_41_120 ();
 FILLCELL_X8 FILLER_41_139 ();
 FILLCELL_X1 FILLER_41_147 ();
 FILLCELL_X4 FILLER_41_154 ();
 FILLCELL_X4 FILLER_41_163 ();
 FILLCELL_X1 FILLER_41_167 ();
 FILLCELL_X2 FILLER_41_180 ();
 FILLCELL_X2 FILLER_41_189 ();
 FILLCELL_X4 FILLER_41_210 ();
 FILLCELL_X1 FILLER_41_214 ();
 FILLCELL_X1 FILLER_41_222 ();
 FILLCELL_X1 FILLER_41_246 ();
 FILLCELL_X2 FILLER_41_271 ();
 FILLCELL_X1 FILLER_41_273 ();
 FILLCELL_X2 FILLER_41_277 ();
 FILLCELL_X8 FILLER_41_282 ();
 FILLCELL_X4 FILLER_41_290 ();
 FILLCELL_X8 FILLER_41_312 ();
 FILLCELL_X1 FILLER_41_320 ();
 FILLCELL_X4 FILLER_41_328 ();
 FILLCELL_X2 FILLER_41_332 ();
 FILLCELL_X8 FILLER_41_337 ();
 FILLCELL_X2 FILLER_41_345 ();
 FILLCELL_X8 FILLER_41_350 ();
 FILLCELL_X4 FILLER_41_382 ();
 FILLCELL_X8 FILLER_41_403 ();
 FILLCELL_X16 FILLER_41_418 ();
 FILLCELL_X1 FILLER_41_434 ();
 FILLCELL_X8 FILLER_41_464 ();
 FILLCELL_X4 FILLER_41_472 ();
 FILLCELL_X1 FILLER_41_476 ();
 FILLCELL_X8 FILLER_41_495 ();
 FILLCELL_X2 FILLER_41_503 ();
 FILLCELL_X4 FILLER_42_1 ();
 FILLCELL_X2 FILLER_42_5 ();
 FILLCELL_X1 FILLER_42_7 ();
 FILLCELL_X8 FILLER_42_28 ();
 FILLCELL_X4 FILLER_42_36 ();
 FILLCELL_X2 FILLER_42_40 ();
 FILLCELL_X16 FILLER_42_59 ();
 FILLCELL_X8 FILLER_42_75 ();
 FILLCELL_X1 FILLER_42_83 ();
 FILLCELL_X8 FILLER_42_101 ();
 FILLCELL_X4 FILLER_42_112 ();
 FILLCELL_X1 FILLER_42_116 ();
 FILLCELL_X16 FILLER_42_124 ();
 FILLCELL_X4 FILLER_42_140 ();
 FILLCELL_X1 FILLER_42_144 ();
 FILLCELL_X32 FILLER_42_162 ();
 FILLCELL_X4 FILLER_42_194 ();
 FILLCELL_X8 FILLER_42_222 ();
 FILLCELL_X2 FILLER_42_230 ();
 FILLCELL_X1 FILLER_42_232 ();
 FILLCELL_X1 FILLER_42_245 ();
 FILLCELL_X1 FILLER_42_257 ();
 FILLCELL_X4 FILLER_42_265 ();
 FILLCELL_X1 FILLER_42_276 ();
 FILLCELL_X1 FILLER_42_284 ();
 FILLCELL_X16 FILLER_42_292 ();
 FILLCELL_X8 FILLER_42_308 ();
 FILLCELL_X1 FILLER_42_316 ();
 FILLCELL_X2 FILLER_42_341 ();
 FILLCELL_X4 FILLER_42_389 ();
 FILLCELL_X2 FILLER_42_393 ();
 FILLCELL_X4 FILLER_42_403 ();
 FILLCELL_X1 FILLER_42_407 ();
 FILLCELL_X2 FILLER_42_473 ();
 FILLCELL_X1 FILLER_42_484 ();
 FILLCELL_X2 FILLER_42_502 ();
 FILLCELL_X1 FILLER_42_504 ();
 FILLCELL_X8 FILLER_43_1 ();
 FILLCELL_X4 FILLER_43_9 ();
 FILLCELL_X2 FILLER_43_13 ();
 FILLCELL_X2 FILLER_43_29 ();
 FILLCELL_X1 FILLER_43_38 ();
 FILLCELL_X2 FILLER_43_43 ();
 FILLCELL_X1 FILLER_43_45 ();
 FILLCELL_X4 FILLER_43_60 ();
 FILLCELL_X1 FILLER_43_64 ();
 FILLCELL_X2 FILLER_43_72 ();
 FILLCELL_X1 FILLER_43_74 ();
 FILLCELL_X2 FILLER_43_112 ();
 FILLCELL_X16 FILLER_43_121 ();
 FILLCELL_X8 FILLER_43_137 ();
 FILLCELL_X2 FILLER_43_145 ();
 FILLCELL_X16 FILLER_43_166 ();
 FILLCELL_X1 FILLER_43_182 ();
 FILLCELL_X4 FILLER_43_190 ();
 FILLCELL_X2 FILLER_43_194 ();
 FILLCELL_X1 FILLER_43_196 ();
 FILLCELL_X4 FILLER_43_204 ();
 FILLCELL_X1 FILLER_43_208 ();
 FILLCELL_X4 FILLER_43_216 ();
 FILLCELL_X2 FILLER_43_227 ();
 FILLCELL_X1 FILLER_43_253 ();
 FILLCELL_X4 FILLER_43_274 ();
 FILLCELL_X1 FILLER_43_278 ();
 FILLCELL_X4 FILLER_43_282 ();
 FILLCELL_X1 FILLER_43_286 ();
 FILLCELL_X8 FILLER_43_304 ();
 FILLCELL_X2 FILLER_43_312 ();
 FILLCELL_X2 FILLER_43_353 ();
 FILLCELL_X4 FILLER_43_372 ();
 FILLCELL_X2 FILLER_43_376 ();
 FILLCELL_X1 FILLER_43_378 ();
 FILLCELL_X1 FILLER_43_393 ();
 FILLCELL_X4 FILLER_43_397 ();
 FILLCELL_X2 FILLER_43_401 ();
 FILLCELL_X4 FILLER_43_417 ();
 FILLCELL_X2 FILLER_43_421 ();
 FILLCELL_X1 FILLER_43_450 ();
 FILLCELL_X2 FILLER_43_481 ();
 FILLCELL_X1 FILLER_43_483 ();
 FILLCELL_X8 FILLER_43_489 ();
 FILLCELL_X1 FILLER_43_504 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X2 FILLER_44_9 ();
 FILLCELL_X2 FILLER_44_18 ();
 FILLCELL_X8 FILLER_44_37 ();
 FILLCELL_X4 FILLER_44_45 ();
 FILLCELL_X1 FILLER_44_49 ();
 FILLCELL_X8 FILLER_44_70 ();
 FILLCELL_X2 FILLER_44_78 ();
 FILLCELL_X2 FILLER_44_87 ();
 FILLCELL_X1 FILLER_44_89 ();
 FILLCELL_X2 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_123 ();
 FILLCELL_X2 FILLER_44_155 ();
 FILLCELL_X2 FILLER_44_166 ();
 FILLCELL_X32 FILLER_44_171 ();
 FILLCELL_X4 FILLER_44_203 ();
 FILLCELL_X1 FILLER_44_207 ();
 FILLCELL_X8 FILLER_44_225 ();
 FILLCELL_X8 FILLER_44_257 ();
 FILLCELL_X4 FILLER_44_265 ();
 FILLCELL_X1 FILLER_44_279 ();
 FILLCELL_X2 FILLER_44_290 ();
 FILLCELL_X1 FILLER_44_292 ();
 FILLCELL_X8 FILLER_44_310 ();
 FILLCELL_X2 FILLER_44_318 ();
 FILLCELL_X2 FILLER_44_351 ();
 FILLCELL_X16 FILLER_44_356 ();
 FILLCELL_X2 FILLER_44_372 ();
 FILLCELL_X8 FILLER_44_398 ();
 FILLCELL_X2 FILLER_44_406 ();
 FILLCELL_X8 FILLER_44_415 ();
 FILLCELL_X2 FILLER_44_423 ();
 FILLCELL_X1 FILLER_44_425 ();
 FILLCELL_X8 FILLER_44_450 ();
 FILLCELL_X4 FILLER_44_458 ();
 FILLCELL_X2 FILLER_44_462 ();
 FILLCELL_X4 FILLER_44_473 ();
 FILLCELL_X8 FILLER_44_483 ();
 FILLCELL_X2 FILLER_44_491 ();
 FILLCELL_X4 FILLER_44_497 ();
 FILLCELL_X1 FILLER_44_501 ();
 FILLCELL_X2 FILLER_45_1 ();
 FILLCELL_X1 FILLER_45_27 ();
 FILLCELL_X8 FILLER_45_38 ();
 FILLCELL_X2 FILLER_45_46 ();
 FILLCELL_X1 FILLER_45_48 ();
 FILLCELL_X1 FILLER_45_59 ();
 FILLCELL_X8 FILLER_45_74 ();
 FILLCELL_X4 FILLER_45_82 ();
 FILLCELL_X2 FILLER_45_86 ();
 FILLCELL_X1 FILLER_45_88 ();
 FILLCELL_X4 FILLER_45_106 ();
 FILLCELL_X1 FILLER_45_110 ();
 FILLCELL_X8 FILLER_45_145 ();
 FILLCELL_X1 FILLER_45_153 ();
 FILLCELL_X8 FILLER_45_171 ();
 FILLCELL_X8 FILLER_45_213 ();
 FILLCELL_X2 FILLER_45_221 ();
 FILLCELL_X16 FILLER_45_226 ();
 FILLCELL_X4 FILLER_45_242 ();
 FILLCELL_X8 FILLER_45_253 ();
 FILLCELL_X4 FILLER_45_261 ();
 FILLCELL_X1 FILLER_45_299 ();
 FILLCELL_X2 FILLER_45_307 ();
 FILLCELL_X1 FILLER_45_309 ();
 FILLCELL_X8 FILLER_45_334 ();
 FILLCELL_X4 FILLER_45_342 ();
 FILLCELL_X4 FILLER_45_353 ();
 FILLCELL_X8 FILLER_45_364 ();
 FILLCELL_X2 FILLER_45_372 ();
 FILLCELL_X8 FILLER_45_379 ();
 FILLCELL_X1 FILLER_45_387 ();
 FILLCELL_X16 FILLER_45_427 ();
 FILLCELL_X2 FILLER_45_443 ();
 FILLCELL_X1 FILLER_45_445 ();
 FILLCELL_X8 FILLER_45_449 ();
 FILLCELL_X2 FILLER_45_457 ();
 FILLCELL_X2 FILLER_45_462 ();
 FILLCELL_X16 FILLER_45_470 ();
 FILLCELL_X2 FILLER_45_486 ();
 FILLCELL_X1 FILLER_45_488 ();
 FILLCELL_X2 FILLER_45_495 ();
 FILLCELL_X4 FILLER_45_500 ();
 FILLCELL_X1 FILLER_45_504 ();
 FILLCELL_X4 FILLER_46_1 ();
 FILLCELL_X2 FILLER_46_5 ();
 FILLCELL_X1 FILLER_46_7 ();
 FILLCELL_X1 FILLER_46_30 ();
 FILLCELL_X4 FILLER_46_85 ();
 FILLCELL_X2 FILLER_46_96 ();
 FILLCELL_X1 FILLER_46_98 ();
 FILLCELL_X2 FILLER_46_128 ();
 FILLCELL_X1 FILLER_46_137 ();
 FILLCELL_X2 FILLER_46_145 ();
 FILLCELL_X1 FILLER_46_147 ();
 FILLCELL_X8 FILLER_46_173 ();
 FILLCELL_X4 FILLER_46_181 ();
 FILLCELL_X8 FILLER_46_206 ();
 FILLCELL_X2 FILLER_46_214 ();
 FILLCELL_X4 FILLER_46_233 ();
 FILLCELL_X1 FILLER_46_244 ();
 FILLCELL_X1 FILLER_46_269 ();
 FILLCELL_X4 FILLER_46_275 ();
 FILLCELL_X1 FILLER_46_279 ();
 FILLCELL_X2 FILLER_46_286 ();
 FILLCELL_X1 FILLER_46_288 ();
 FILLCELL_X8 FILLER_46_296 ();
 FILLCELL_X4 FILLER_46_304 ();
 FILLCELL_X1 FILLER_46_308 ();
 FILLCELL_X8 FILLER_46_333 ();
 FILLCELL_X8 FILLER_46_358 ();
 FILLCELL_X1 FILLER_46_366 ();
 FILLCELL_X4 FILLER_46_374 ();
 FILLCELL_X1 FILLER_46_378 ();
 FILLCELL_X2 FILLER_46_394 ();
 FILLCELL_X1 FILLER_46_396 ();
 FILLCELL_X4 FILLER_46_419 ();
 FILLCELL_X2 FILLER_46_423 ();
 FILLCELL_X2 FILLER_46_442 ();
 FILLCELL_X2 FILLER_46_451 ();
 FILLCELL_X1 FILLER_46_453 ();
 FILLCELL_X2 FILLER_46_481 ();
 FILLCELL_X8 FILLER_46_492 ();
 FILLCELL_X4 FILLER_46_500 ();
 FILLCELL_X1 FILLER_46_504 ();
 FILLCELL_X16 FILLER_47_1 ();
 FILLCELL_X8 FILLER_47_17 ();
 FILLCELL_X4 FILLER_47_25 ();
 FILLCELL_X2 FILLER_47_29 ();
 FILLCELL_X1 FILLER_47_31 ();
 FILLCELL_X1 FILLER_47_49 ();
 FILLCELL_X2 FILLER_47_57 ();
 FILLCELL_X1 FILLER_47_59 ();
 FILLCELL_X16 FILLER_47_67 ();
 FILLCELL_X8 FILLER_47_83 ();
 FILLCELL_X4 FILLER_47_91 ();
 FILLCELL_X2 FILLER_47_95 ();
 FILLCELL_X1 FILLER_47_97 ();
 FILLCELL_X4 FILLER_47_108 ();
 FILLCELL_X2 FILLER_47_112 ();
 FILLCELL_X1 FILLER_47_114 ();
 FILLCELL_X2 FILLER_47_128 ();
 FILLCELL_X8 FILLER_47_154 ();
 FILLCELL_X4 FILLER_47_162 ();
 FILLCELL_X2 FILLER_47_166 ();
 FILLCELL_X16 FILLER_47_175 ();
 FILLCELL_X8 FILLER_47_191 ();
 FILLCELL_X2 FILLER_47_199 ();
 FILLCELL_X1 FILLER_47_201 ();
 FILLCELL_X2 FILLER_47_205 ();
 FILLCELL_X4 FILLER_47_243 ();
 FILLCELL_X4 FILLER_47_271 ();
 FILLCELL_X4 FILLER_47_284 ();
 FILLCELL_X8 FILLER_47_305 ();
 FILLCELL_X2 FILLER_47_313 ();
 FILLCELL_X1 FILLER_47_315 ();
 FILLCELL_X4 FILLER_47_337 ();
 FILLCELL_X1 FILLER_47_341 ();
 FILLCELL_X1 FILLER_47_351 ();
 FILLCELL_X2 FILLER_47_358 ();
 FILLCELL_X8 FILLER_47_363 ();
 FILLCELL_X1 FILLER_47_371 ();
 FILLCELL_X2 FILLER_47_379 ();
 FILLCELL_X1 FILLER_47_381 ();
 FILLCELL_X4 FILLER_47_399 ();
 FILLCELL_X2 FILLER_47_409 ();
 FILLCELL_X1 FILLER_47_414 ();
 FILLCELL_X8 FILLER_47_418 ();
 FILLCELL_X1 FILLER_47_426 ();
 FILLCELL_X4 FILLER_47_434 ();
 FILLCELL_X2 FILLER_47_445 ();
 FILLCELL_X1 FILLER_47_447 ();
 FILLCELL_X2 FILLER_47_475 ();
 FILLCELL_X2 FILLER_47_480 ();
 FILLCELL_X1 FILLER_47_482 ();
 FILLCELL_X4 FILLER_47_500 ();
 FILLCELL_X1 FILLER_47_504 ();
 FILLCELL_X2 FILLER_48_1 ();
 FILLCELL_X1 FILLER_48_3 ();
 FILLCELL_X4 FILLER_48_28 ();
 FILLCELL_X2 FILLER_48_32 ();
 FILLCELL_X2 FILLER_48_48 ();
 FILLCELL_X8 FILLER_48_53 ();
 FILLCELL_X4 FILLER_48_61 ();
 FILLCELL_X2 FILLER_48_65 ();
 FILLCELL_X1 FILLER_48_67 ();
 FILLCELL_X2 FILLER_48_76 ();
 FILLCELL_X4 FILLER_48_85 ();
 FILLCELL_X16 FILLER_48_106 ();
 FILLCELL_X4 FILLER_48_122 ();
 FILLCELL_X2 FILLER_48_126 ();
 FILLCELL_X1 FILLER_48_128 ();
 FILLCELL_X16 FILLER_48_153 ();
 FILLCELL_X1 FILLER_48_169 ();
 FILLCELL_X4 FILLER_48_187 ();
 FILLCELL_X8 FILLER_48_264 ();
 FILLCELL_X4 FILLER_48_272 ();
 FILLCELL_X2 FILLER_48_276 ();
 FILLCELL_X1 FILLER_48_278 ();
 FILLCELL_X32 FILLER_48_299 ();
 FILLCELL_X2 FILLER_48_338 ();
 FILLCELL_X2 FILLER_48_347 ();
 FILLCELL_X1 FILLER_48_366 ();
 FILLCELL_X1 FILLER_48_391 ();
 FILLCELL_X2 FILLER_48_398 ();
 FILLCELL_X4 FILLER_48_410 ();
 FILLCELL_X1 FILLER_48_414 ();
 FILLCELL_X1 FILLER_48_423 ();
 FILLCELL_X8 FILLER_48_458 ();
 FILLCELL_X1 FILLER_48_466 ();
 FILLCELL_X16 FILLER_48_484 ();
 FILLCELL_X4 FILLER_48_500 ();
 FILLCELL_X1 FILLER_48_504 ();
 FILLCELL_X4 FILLER_49_1 ();
 FILLCELL_X2 FILLER_49_5 ();
 FILLCELL_X16 FILLER_49_38 ();
 FILLCELL_X8 FILLER_49_57 ();
 FILLCELL_X2 FILLER_49_65 ();
 FILLCELL_X1 FILLER_49_67 ();
 FILLCELL_X2 FILLER_49_85 ();
 FILLCELL_X1 FILLER_49_87 ();
 FILLCELL_X16 FILLER_49_136 ();
 FILLCELL_X1 FILLER_49_152 ();
 FILLCELL_X1 FILLER_49_162 ();
 FILLCELL_X4 FILLER_49_176 ();
 FILLCELL_X1 FILLER_49_180 ();
 FILLCELL_X8 FILLER_49_188 ();
 FILLCELL_X4 FILLER_49_196 ();
 FILLCELL_X8 FILLER_49_214 ();
 FILLCELL_X4 FILLER_49_222 ();
 FILLCELL_X1 FILLER_49_226 ();
 FILLCELL_X8 FILLER_49_232 ();
 FILLCELL_X2 FILLER_49_240 ();
 FILLCELL_X1 FILLER_49_242 ();
 FILLCELL_X2 FILLER_49_263 ();
 FILLCELL_X8 FILLER_49_294 ();
 FILLCELL_X4 FILLER_49_302 ();
 FILLCELL_X2 FILLER_49_306 ();
 FILLCELL_X1 FILLER_49_308 ();
 FILLCELL_X2 FILLER_49_333 ();
 FILLCELL_X4 FILLER_49_359 ();
 FILLCELL_X1 FILLER_49_363 ();
 FILLCELL_X16 FILLER_49_371 ();
 FILLCELL_X8 FILLER_49_394 ();
 FILLCELL_X1 FILLER_49_402 ();
 FILLCELL_X4 FILLER_49_406 ();
 FILLCELL_X2 FILLER_49_410 ();
 FILLCELL_X1 FILLER_49_412 ();
 FILLCELL_X2 FILLER_49_437 ();
 FILLCELL_X2 FILLER_49_446 ();
 FILLCELL_X32 FILLER_49_452 ();
 FILLCELL_X16 FILLER_49_484 ();
 FILLCELL_X4 FILLER_49_500 ();
 FILLCELL_X1 FILLER_49_504 ();
 FILLCELL_X1 FILLER_50_1 ();
 FILLCELL_X16 FILLER_50_5 ();
 FILLCELL_X8 FILLER_50_21 ();
 FILLCELL_X4 FILLER_50_29 ();
 FILLCELL_X4 FILLER_50_57 ();
 FILLCELL_X2 FILLER_50_78 ();
 FILLCELL_X4 FILLER_50_87 ();
 FILLCELL_X1 FILLER_50_91 ();
 FILLCELL_X16 FILLER_50_109 ();
 FILLCELL_X1 FILLER_50_125 ();
 FILLCELL_X8 FILLER_50_133 ();
 FILLCELL_X4 FILLER_50_141 ();
 FILLCELL_X1 FILLER_50_145 ();
 FILLCELL_X2 FILLER_50_163 ();
 FILLCELL_X1 FILLER_50_165 ();
 FILLCELL_X2 FILLER_50_185 ();
 FILLCELL_X1 FILLER_50_187 ();
 FILLCELL_X1 FILLER_50_191 ();
 FILLCELL_X1 FILLER_50_209 ();
 FILLCELL_X1 FILLER_50_213 ();
 FILLCELL_X16 FILLER_50_221 ();
 FILLCELL_X1 FILLER_50_237 ();
 FILLCELL_X4 FILLER_50_243 ();
 FILLCELL_X16 FILLER_50_291 ();
 FILLCELL_X1 FILLER_50_338 ();
 FILLCELL_X1 FILLER_50_342 ();
 FILLCELL_X2 FILLER_50_353 ();
 FILLCELL_X8 FILLER_50_362 ();
 FILLCELL_X4 FILLER_50_370 ();
 FILLCELL_X1 FILLER_50_374 ();
 FILLCELL_X4 FILLER_50_399 ();
 FILLCELL_X1 FILLER_50_410 ();
 FILLCELL_X2 FILLER_50_425 ();
 FILLCELL_X4 FILLER_50_434 ();
 FILLCELL_X2 FILLER_50_438 ();
 FILLCELL_X16 FILLER_50_466 ();
 FILLCELL_X4 FILLER_50_482 ();
 FILLCELL_X2 FILLER_50_486 ();
 FILLCELL_X1 FILLER_50_488 ();
 FILLCELL_X8 FILLER_50_497 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X4 FILLER_51_33 ();
 FILLCELL_X1 FILLER_51_37 ();
 FILLCELL_X8 FILLER_51_65 ();
 FILLCELL_X4 FILLER_51_73 ();
 FILLCELL_X1 FILLER_51_77 ();
 FILLCELL_X8 FILLER_51_85 ();
 FILLCELL_X4 FILLER_51_93 ();
 FILLCELL_X1 FILLER_51_97 ();
 FILLCELL_X2 FILLER_51_105 ();
 FILLCELL_X16 FILLER_51_110 ();
 FILLCELL_X4 FILLER_51_126 ();
 FILLCELL_X2 FILLER_51_130 ();
 FILLCELL_X8 FILLER_51_135 ();
 FILLCELL_X2 FILLER_51_143 ();
 FILLCELL_X1 FILLER_51_145 ();
 FILLCELL_X4 FILLER_51_161 ();
 FILLCELL_X2 FILLER_51_168 ();
 FILLCELL_X1 FILLER_51_170 ();
 FILLCELL_X16 FILLER_51_176 ();
 FILLCELL_X8 FILLER_51_192 ();
 FILLCELL_X8 FILLER_51_224 ();
 FILLCELL_X2 FILLER_51_232 ();
 FILLCELL_X1 FILLER_51_234 ();
 FILLCELL_X16 FILLER_51_252 ();
 FILLCELL_X8 FILLER_51_268 ();
 FILLCELL_X16 FILLER_51_293 ();
 FILLCELL_X4 FILLER_51_309 ();
 FILLCELL_X2 FILLER_51_313 ();
 FILLCELL_X1 FILLER_51_315 ();
 FILLCELL_X4 FILLER_51_323 ();
 FILLCELL_X2 FILLER_51_327 ();
 FILLCELL_X2 FILLER_51_353 ();
 FILLCELL_X2 FILLER_51_372 ();
 FILLCELL_X4 FILLER_51_398 ();
 FILLCELL_X2 FILLER_51_402 ();
 FILLCELL_X8 FILLER_51_438 ();
 FILLCELL_X2 FILLER_51_446 ();
 FILLCELL_X1 FILLER_51_448 ();
 FILLCELL_X16 FILLER_51_481 ();
 FILLCELL_X8 FILLER_51_497 ();
 FILLCELL_X8 FILLER_52_1 ();
 FILLCELL_X4 FILLER_52_16 ();
 FILLCELL_X1 FILLER_52_20 ();
 FILLCELL_X16 FILLER_52_28 ();
 FILLCELL_X2 FILLER_52_44 ();
 FILLCELL_X8 FILLER_52_63 ();
 FILLCELL_X2 FILLER_52_71 ();
 FILLCELL_X1 FILLER_52_73 ();
 FILLCELL_X4 FILLER_52_81 ();
 FILLCELL_X1 FILLER_52_85 ();
 FILLCELL_X1 FILLER_52_93 ();
 FILLCELL_X4 FILLER_52_126 ();
 FILLCELL_X2 FILLER_52_130 ();
 FILLCELL_X8 FILLER_52_135 ();
 FILLCELL_X2 FILLER_52_143 ();
 FILLCELL_X4 FILLER_52_154 ();
 FILLCELL_X4 FILLER_52_194 ();
 FILLCELL_X2 FILLER_52_198 ();
 FILLCELL_X4 FILLER_52_230 ();
 FILLCELL_X1 FILLER_52_234 ();
 FILLCELL_X4 FILLER_52_238 ();
 FILLCELL_X1 FILLER_52_242 ();
 FILLCELL_X2 FILLER_52_257 ();
 FILLCELL_X1 FILLER_52_259 ();
 FILLCELL_X2 FILLER_52_284 ();
 FILLCELL_X1 FILLER_52_292 ();
 FILLCELL_X2 FILLER_52_303 ();
 FILLCELL_X1 FILLER_52_305 ();
 FILLCELL_X8 FILLER_52_311 ();
 FILLCELL_X16 FILLER_52_324 ();
 FILLCELL_X2 FILLER_52_340 ();
 FILLCELL_X16 FILLER_52_347 ();
 FILLCELL_X8 FILLER_52_368 ();
 FILLCELL_X4 FILLER_52_376 ();
 FILLCELL_X1 FILLER_52_380 ();
 FILLCELL_X2 FILLER_52_444 ();
 FILLCELL_X16 FILLER_52_460 ();
 FILLCELL_X8 FILLER_52_476 ();
 FILLCELL_X2 FILLER_52_484 ();
 FILLCELL_X2 FILLER_52_503 ();
 FILLCELL_X4 FILLER_53_1 ();
 FILLCELL_X1 FILLER_53_5 ();
 FILLCELL_X4 FILLER_53_30 ();
 FILLCELL_X8 FILLER_53_41 ();
 FILLCELL_X4 FILLER_53_49 ();
 FILLCELL_X8 FILLER_53_57 ();
 FILLCELL_X2 FILLER_53_65 ();
 FILLCELL_X1 FILLER_53_67 ();
 FILLCELL_X4 FILLER_53_109 ();
 FILLCELL_X1 FILLER_53_120 ();
 FILLCELL_X2 FILLER_53_128 ();
 FILLCELL_X1 FILLER_53_130 ();
 FILLCELL_X2 FILLER_53_138 ();
 FILLCELL_X1 FILLER_53_155 ();
 FILLCELL_X2 FILLER_53_180 ();
 FILLCELL_X2 FILLER_53_200 ();
 FILLCELL_X1 FILLER_53_202 ();
 FILLCELL_X16 FILLER_53_225 ();
 FILLCELL_X4 FILLER_53_241 ();
 FILLCELL_X1 FILLER_53_245 ();
 FILLCELL_X2 FILLER_53_259 ();
 FILLCELL_X1 FILLER_53_261 ();
 FILLCELL_X2 FILLER_53_268 ();
 FILLCELL_X1 FILLER_53_279 ();
 FILLCELL_X1 FILLER_53_292 ();
 FILLCELL_X16 FILLER_53_317 ();
 FILLCELL_X1 FILLER_53_333 ();
 FILLCELL_X8 FILLER_53_341 ();
 FILLCELL_X4 FILLER_53_349 ();
 FILLCELL_X2 FILLER_53_353 ();
 FILLCELL_X16 FILLER_53_376 ();
 FILLCELL_X8 FILLER_53_392 ();
 FILLCELL_X4 FILLER_53_400 ();
 FILLCELL_X2 FILLER_53_404 ();
 FILLCELL_X1 FILLER_53_406 ();
 FILLCELL_X16 FILLER_53_431 ();
 FILLCELL_X8 FILLER_53_447 ();
 FILLCELL_X4 FILLER_53_455 ();
 FILLCELL_X16 FILLER_53_463 ();
 FILLCELL_X8 FILLER_53_479 ();
 FILLCELL_X2 FILLER_53_487 ();
 FILLCELL_X4 FILLER_53_493 ();
 FILLCELL_X1 FILLER_53_497 ();
 FILLCELL_X1 FILLER_53_501 ();
 FILLCELL_X8 FILLER_54_1 ();
 FILLCELL_X2 FILLER_54_9 ();
 FILLCELL_X1 FILLER_54_11 ();
 FILLCELL_X2 FILLER_54_53 ();
 FILLCELL_X1 FILLER_54_55 ();
 FILLCELL_X1 FILLER_54_63 ();
 FILLCELL_X1 FILLER_54_104 ();
 FILLCELL_X2 FILLER_54_133 ();
 FILLCELL_X8 FILLER_54_138 ();
 FILLCELL_X1 FILLER_54_146 ();
 FILLCELL_X1 FILLER_54_179 ();
 FILLCELL_X1 FILLER_54_192 ();
 FILLCELL_X2 FILLER_54_203 ();
 FILLCELL_X2 FILLER_54_229 ();
 FILLCELL_X1 FILLER_54_231 ();
 FILLCELL_X2 FILLER_54_257 ();
 FILLCELL_X2 FILLER_54_281 ();
 FILLCELL_X1 FILLER_54_292 ();
 FILLCELL_X32 FILLER_54_304 ();
 FILLCELL_X4 FILLER_54_340 ();
 FILLCELL_X1 FILLER_54_344 ();
 FILLCELL_X8 FILLER_54_349 ();
 FILLCELL_X4 FILLER_54_357 ();
 FILLCELL_X32 FILLER_54_378 ();
 FILLCELL_X4 FILLER_54_410 ();
 FILLCELL_X4 FILLER_54_428 ();
 FILLCELL_X2 FILLER_54_432 ();
 FILLCELL_X1 FILLER_54_434 ();
 FILLCELL_X1 FILLER_54_442 ();
 FILLCELL_X2 FILLER_54_454 ();
 FILLCELL_X1 FILLER_54_456 ();
 FILLCELL_X2 FILLER_54_500 ();
 FILLCELL_X1 FILLER_54_504 ();
 FILLCELL_X16 FILLER_55_1 ();
 FILLCELL_X8 FILLER_55_17 ();
 FILLCELL_X4 FILLER_55_25 ();
 FILLCELL_X2 FILLER_55_51 ();
 FILLCELL_X1 FILLER_55_53 ();
 FILLCELL_X4 FILLER_55_71 ();
 FILLCELL_X2 FILLER_55_75 ();
 FILLCELL_X1 FILLER_55_77 ();
 FILLCELL_X8 FILLER_55_85 ();
 FILLCELL_X2 FILLER_55_93 ();
 FILLCELL_X32 FILLER_55_98 ();
 FILLCELL_X16 FILLER_55_130 ();
 FILLCELL_X4 FILLER_55_146 ();
 FILLCELL_X2 FILLER_55_150 ();
 FILLCELL_X1 FILLER_55_168 ();
 FILLCELL_X16 FILLER_55_175 ();
 FILLCELL_X4 FILLER_55_191 ();
 FILLCELL_X2 FILLER_55_195 ();
 FILLCELL_X1 FILLER_55_197 ();
 FILLCELL_X8 FILLER_55_218 ();
 FILLCELL_X4 FILLER_55_226 ();
 FILLCELL_X1 FILLER_55_230 ();
 FILLCELL_X4 FILLER_55_238 ();
 FILLCELL_X16 FILLER_55_266 ();
 FILLCELL_X1 FILLER_55_282 ();
 FILLCELL_X32 FILLER_55_290 ();
 FILLCELL_X4 FILLER_55_322 ();
 FILLCELL_X1 FILLER_55_326 ();
 FILLCELL_X4 FILLER_55_337 ();
 FILLCELL_X4 FILLER_55_345 ();
 FILLCELL_X1 FILLER_55_349 ();
 FILLCELL_X4 FILLER_55_354 ();
 FILLCELL_X4 FILLER_55_375 ();
 FILLCELL_X1 FILLER_55_379 ();
 FILLCELL_X16 FILLER_55_384 ();
 FILLCELL_X8 FILLER_55_400 ();
 FILLCELL_X2 FILLER_55_408 ();
 FILLCELL_X2 FILLER_55_415 ();
 FILLCELL_X1 FILLER_55_466 ();
 FILLCELL_X2 FILLER_55_471 ();
 FILLCELL_X1 FILLER_55_473 ();
 FILLCELL_X2 FILLER_56_1 ();
 FILLCELL_X1 FILLER_56_3 ();
 FILLCELL_X16 FILLER_56_21 ();
 FILLCELL_X8 FILLER_56_37 ();
 FILLCELL_X2 FILLER_56_45 ();
 FILLCELL_X16 FILLER_56_54 ();
 FILLCELL_X4 FILLER_56_70 ();
 FILLCELL_X2 FILLER_56_88 ();
 FILLCELL_X1 FILLER_56_90 ();
 FILLCELL_X4 FILLER_56_98 ();
 FILLCELL_X2 FILLER_56_102 ();
 FILLCELL_X4 FILLER_56_111 ();
 FILLCELL_X2 FILLER_56_115 ();
 FILLCELL_X4 FILLER_56_124 ();
 FILLCELL_X4 FILLER_56_135 ();
 FILLCELL_X2 FILLER_56_139 ();
 FILLCELL_X1 FILLER_56_141 ();
 FILLCELL_X4 FILLER_56_156 ();
 FILLCELL_X8 FILLER_56_167 ();
 FILLCELL_X1 FILLER_56_182 ();
 FILLCELL_X4 FILLER_56_200 ();
 FILLCELL_X2 FILLER_56_204 ();
 FILLCELL_X1 FILLER_56_206 ();
 FILLCELL_X4 FILLER_56_221 ();
 FILLCELL_X2 FILLER_56_225 ();
 FILLCELL_X2 FILLER_56_244 ();
 FILLCELL_X1 FILLER_56_246 ();
 FILLCELL_X8 FILLER_56_254 ();
 FILLCELL_X2 FILLER_56_262 ();
 FILLCELL_X2 FILLER_56_271 ();
 FILLCELL_X4 FILLER_56_278 ();
 FILLCELL_X2 FILLER_56_282 ();
 FILLCELL_X1 FILLER_56_284 ();
 FILLCELL_X2 FILLER_56_292 ();
 FILLCELL_X1 FILLER_56_369 ();
 FILLCELL_X2 FILLER_56_385 ();
 FILLCELL_X2 FILLER_56_394 ();
 FILLCELL_X8 FILLER_56_403 ();
 FILLCELL_X2 FILLER_56_422 ();
 FILLCELL_X4 FILLER_56_446 ();
 FILLCELL_X2 FILLER_56_458 ();
 FILLCELL_X2 FILLER_56_496 ();
 FILLCELL_X1 FILLER_56_498 ();
 FILLCELL_X4 FILLER_57_1 ();
 FILLCELL_X4 FILLER_57_29 ();
 FILLCELL_X4 FILLER_57_40 ();
 FILLCELL_X1 FILLER_57_44 ();
 FILLCELL_X4 FILLER_57_52 ();
 FILLCELL_X2 FILLER_57_56 ();
 FILLCELL_X1 FILLER_57_58 ();
 FILLCELL_X2 FILLER_57_69 ();
 FILLCELL_X2 FILLER_57_88 ();
 FILLCELL_X1 FILLER_57_90 ();
 FILLCELL_X2 FILLER_57_108 ();
 FILLCELL_X1 FILLER_57_110 ();
 FILLCELL_X2 FILLER_57_128 ();
 FILLCELL_X1 FILLER_57_130 ();
 FILLCELL_X8 FILLER_57_148 ();
 FILLCELL_X4 FILLER_57_156 ();
 FILLCELL_X8 FILLER_57_177 ();
 FILLCELL_X2 FILLER_57_185 ();
 FILLCELL_X1 FILLER_57_187 ();
 FILLCELL_X4 FILLER_57_202 ();
 FILLCELL_X2 FILLER_57_206 ();
 FILLCELL_X16 FILLER_57_225 ();
 FILLCELL_X2 FILLER_57_241 ();
 FILLCELL_X4 FILLER_57_260 ();
 FILLCELL_X2 FILLER_57_264 ();
 FILLCELL_X1 FILLER_57_266 ();
 FILLCELL_X4 FILLER_57_291 ();
 FILLCELL_X2 FILLER_57_295 ();
 FILLCELL_X16 FILLER_57_304 ();
 FILLCELL_X4 FILLER_57_320 ();
 FILLCELL_X1 FILLER_57_333 ();
 FILLCELL_X2 FILLER_57_344 ();
 FILLCELL_X1 FILLER_57_346 ();
 FILLCELL_X2 FILLER_57_362 ();
 FILLCELL_X1 FILLER_57_388 ();
 FILLCELL_X16 FILLER_57_406 ();
 FILLCELL_X2 FILLER_57_422 ();
 FILLCELL_X1 FILLER_57_424 ();
 FILLCELL_X16 FILLER_57_437 ();
 FILLCELL_X4 FILLER_57_453 ();
 FILLCELL_X2 FILLER_57_457 ();
 FILLCELL_X1 FILLER_57_459 ();
 FILLCELL_X8 FILLER_57_465 ();
 FILLCELL_X2 FILLER_57_473 ();
 FILLCELL_X1 FILLER_57_485 ();
 FILLCELL_X8 FILLER_57_494 ();
 FILLCELL_X4 FILLER_58_1 ();
 FILLCELL_X1 FILLER_58_5 ();
 FILLCELL_X4 FILLER_58_20 ();
 FILLCELL_X2 FILLER_58_24 ();
 FILLCELL_X8 FILLER_58_50 ();
 FILLCELL_X2 FILLER_58_58 ();
 FILLCELL_X8 FILLER_58_77 ();
 FILLCELL_X4 FILLER_58_85 ();
 FILLCELL_X2 FILLER_58_89 ();
 FILLCELL_X1 FILLER_58_91 ();
 FILLCELL_X4 FILLER_58_109 ();
 FILLCELL_X8 FILLER_58_130 ();
 FILLCELL_X2 FILLER_58_138 ();
 FILLCELL_X8 FILLER_58_152 ();
 FILLCELL_X4 FILLER_58_160 ();
 FILLCELL_X1 FILLER_58_164 ();
 FILLCELL_X1 FILLER_58_172 ();
 FILLCELL_X4 FILLER_58_180 ();
 FILLCELL_X8 FILLER_58_201 ();
 FILLCELL_X2 FILLER_58_226 ();
 FILLCELL_X1 FILLER_58_228 ();
 FILLCELL_X8 FILLER_58_232 ();
 FILLCELL_X4 FILLER_58_240 ();
 FILLCELL_X2 FILLER_58_244 ();
 FILLCELL_X1 FILLER_58_246 ();
 FILLCELL_X8 FILLER_58_258 ();
 FILLCELL_X1 FILLER_58_276 ();
 FILLCELL_X16 FILLER_58_294 ();
 FILLCELL_X8 FILLER_58_310 ();
 FILLCELL_X2 FILLER_58_318 ();
 FILLCELL_X1 FILLER_58_320 ();
 FILLCELL_X8 FILLER_58_340 ();
 FILLCELL_X1 FILLER_58_348 ();
 FILLCELL_X2 FILLER_58_368 ();
 FILLCELL_X4 FILLER_58_377 ();
 FILLCELL_X2 FILLER_58_381 ();
 FILLCELL_X1 FILLER_58_383 ();
 FILLCELL_X8 FILLER_58_388 ();
 FILLCELL_X4 FILLER_58_396 ();
 FILLCELL_X1 FILLER_58_400 ();
 FILLCELL_X8 FILLER_58_417 ();
 FILLCELL_X4 FILLER_58_425 ();
 FILLCELL_X4 FILLER_58_446 ();
 FILLCELL_X4 FILLER_58_454 ();
 FILLCELL_X1 FILLER_58_458 ();
 FILLCELL_X1 FILLER_58_463 ();
 FILLCELL_X1 FILLER_58_468 ();
 FILLCELL_X4 FILLER_58_480 ();
 FILLCELL_X1 FILLER_58_484 ();
 FILLCELL_X2 FILLER_58_502 ();
 FILLCELL_X1 FILLER_58_504 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X2 FILLER_59_33 ();
 FILLCELL_X1 FILLER_59_35 ();
 FILLCELL_X32 FILLER_59_53 ();
 FILLCELL_X8 FILLER_59_85 ();
 FILLCELL_X4 FILLER_59_97 ();
 FILLCELL_X2 FILLER_59_101 ();
 FILLCELL_X1 FILLER_59_110 ();
 FILLCELL_X16 FILLER_59_118 ();
 FILLCELL_X4 FILLER_59_134 ();
 FILLCELL_X2 FILLER_59_138 ();
 FILLCELL_X1 FILLER_59_140 ();
 FILLCELL_X4 FILLER_59_162 ();
 FILLCELL_X1 FILLER_59_166 ();
 FILLCELL_X4 FILLER_59_184 ();
 FILLCELL_X2 FILLER_59_188 ();
 FILLCELL_X1 FILLER_59_190 ();
 FILLCELL_X8 FILLER_59_198 ();
 FILLCELL_X4 FILLER_59_206 ();
 FILLCELL_X4 FILLER_59_217 ();
 FILLCELL_X1 FILLER_59_221 ();
 FILLCELL_X4 FILLER_59_251 ();
 FILLCELL_X2 FILLER_59_255 ();
 FILLCELL_X2 FILLER_59_281 ();
 FILLCELL_X1 FILLER_59_283 ();
 FILLCELL_X2 FILLER_59_287 ();
 FILLCELL_X8 FILLER_59_303 ();
 FILLCELL_X4 FILLER_59_311 ();
 FILLCELL_X2 FILLER_59_315 ();
 FILLCELL_X1 FILLER_59_342 ();
 FILLCELL_X16 FILLER_59_350 ();
 FILLCELL_X8 FILLER_59_366 ();
 FILLCELL_X2 FILLER_59_374 ();
 FILLCELL_X8 FILLER_59_414 ();
 FILLCELL_X4 FILLER_59_422 ();
 FILLCELL_X2 FILLER_59_433 ();
 FILLCELL_X8 FILLER_59_441 ();
 FILLCELL_X1 FILLER_59_449 ();
 FILLCELL_X2 FILLER_59_455 ();
 FILLCELL_X2 FILLER_59_500 ();
 FILLCELL_X16 FILLER_60_1 ();
 FILLCELL_X2 FILLER_60_17 ();
 FILLCELL_X1 FILLER_60_19 ();
 FILLCELL_X8 FILLER_60_27 ();
 FILLCELL_X1 FILLER_60_35 ();
 FILLCELL_X4 FILLER_60_58 ();
 FILLCELL_X2 FILLER_60_62 ();
 FILLCELL_X1 FILLER_60_64 ();
 FILLCELL_X8 FILLER_60_69 ();
 FILLCELL_X8 FILLER_60_94 ();
 FILLCELL_X4 FILLER_60_102 ();
 FILLCELL_X8 FILLER_60_123 ();
 FILLCELL_X8 FILLER_60_138 ();
 FILLCELL_X2 FILLER_60_146 ();
 FILLCELL_X1 FILLER_60_148 ();
 FILLCELL_X32 FILLER_60_156 ();
 FILLCELL_X4 FILLER_60_188 ();
 FILLCELL_X2 FILLER_60_192 ();
 FILLCELL_X1 FILLER_60_194 ();
 FILLCELL_X16 FILLER_60_216 ();
 FILLCELL_X1 FILLER_60_232 ();
 FILLCELL_X2 FILLER_60_257 ();
 FILLCELL_X1 FILLER_60_290 ();
 FILLCELL_X4 FILLER_60_315 ();
 FILLCELL_X2 FILLER_60_319 ();
 FILLCELL_X1 FILLER_60_321 ();
 FILLCELL_X4 FILLER_60_327 ();
 FILLCELL_X2 FILLER_60_331 ();
 FILLCELL_X1 FILLER_60_333 ();
 FILLCELL_X2 FILLER_60_342 ();
 FILLCELL_X8 FILLER_60_355 ();
 FILLCELL_X8 FILLER_60_419 ();
 FILLCELL_X8 FILLER_60_432 ();
 FILLCELL_X4 FILLER_60_440 ();
 FILLCELL_X4 FILLER_60_446 ();
 FILLCELL_X4 FILLER_60_453 ();
 FILLCELL_X4 FILLER_60_487 ();
 FILLCELL_X2 FILLER_60_491 ();
 FILLCELL_X2 FILLER_60_496 ();
 FILLCELL_X1 FILLER_60_498 ();
 FILLCELL_X4 FILLER_61_1 ();
 FILLCELL_X1 FILLER_61_5 ();
 FILLCELL_X2 FILLER_61_40 ();
 FILLCELL_X1 FILLER_61_42 ();
 FILLCELL_X2 FILLER_61_50 ();
 FILLCELL_X1 FILLER_61_52 ();
 FILLCELL_X1 FILLER_61_60 ();
 FILLCELL_X2 FILLER_61_85 ();
 FILLCELL_X1 FILLER_61_87 ();
 FILLCELL_X2 FILLER_61_158 ();
 FILLCELL_X1 FILLER_61_160 ();
 FILLCELL_X8 FILLER_61_164 ();
 FILLCELL_X4 FILLER_61_172 ();
 FILLCELL_X2 FILLER_61_176 ();
 FILLCELL_X8 FILLER_61_195 ();
 FILLCELL_X2 FILLER_61_210 ();
 FILLCELL_X16 FILLER_61_219 ();
 FILLCELL_X8 FILLER_61_235 ();
 FILLCELL_X4 FILLER_61_243 ();
 FILLCELL_X2 FILLER_61_254 ();
 FILLCELL_X1 FILLER_61_256 ();
 FILLCELL_X16 FILLER_61_260 ();
 FILLCELL_X8 FILLER_61_276 ();
 FILLCELL_X4 FILLER_61_284 ();
 FILLCELL_X8 FILLER_61_312 ();
 FILLCELL_X2 FILLER_61_320 ();
 FILLCELL_X1 FILLER_61_322 ();
 FILLCELL_X4 FILLER_61_325 ();
 FILLCELL_X2 FILLER_61_338 ();
 FILLCELL_X2 FILLER_61_357 ();
 FILLCELL_X1 FILLER_61_359 ();
 FILLCELL_X8 FILLER_61_387 ();
 FILLCELL_X4 FILLER_61_395 ();
 FILLCELL_X16 FILLER_61_421 ();
 FILLCELL_X1 FILLER_61_437 ();
 FILLCELL_X4 FILLER_61_440 ();
 FILLCELL_X1 FILLER_61_444 ();
 FILLCELL_X2 FILLER_61_448 ();
 FILLCELL_X1 FILLER_61_450 ();
 FILLCELL_X4 FILLER_61_455 ();
 FILLCELL_X8 FILLER_61_487 ();
 FILLCELL_X4 FILLER_61_499 ();
 FILLCELL_X2 FILLER_61_503 ();
 FILLCELL_X16 FILLER_62_1 ();
 FILLCELL_X1 FILLER_62_31 ();
 FILLCELL_X1 FILLER_62_59 ();
 FILLCELL_X2 FILLER_62_63 ();
 FILLCELL_X1 FILLER_62_65 ();
 FILLCELL_X2 FILLER_62_73 ();
 FILLCELL_X8 FILLER_62_85 ();
 FILLCELL_X8 FILLER_62_110 ();
 FILLCELL_X4 FILLER_62_149 ();
 FILLCELL_X1 FILLER_62_163 ();
 FILLCELL_X2 FILLER_62_171 ();
 FILLCELL_X1 FILLER_62_173 ();
 FILLCELL_X2 FILLER_62_198 ();
 FILLCELL_X2 FILLER_62_224 ();
 FILLCELL_X4 FILLER_62_250 ();
 FILLCELL_X8 FILLER_62_278 ();
 FILLCELL_X2 FILLER_62_286 ();
 FILLCELL_X32 FILLER_62_291 ();
 FILLCELL_X4 FILLER_62_323 ();
 FILLCELL_X1 FILLER_62_327 ();
 FILLCELL_X8 FILLER_62_348 ();
 FILLCELL_X4 FILLER_62_376 ();
 FILLCELL_X16 FILLER_62_393 ();
 FILLCELL_X8 FILLER_62_409 ();
 FILLCELL_X4 FILLER_62_417 ();
 FILLCELL_X1 FILLER_62_421 ();
 FILLCELL_X2 FILLER_62_436 ();
 FILLCELL_X2 FILLER_62_443 ();
 FILLCELL_X2 FILLER_62_461 ();
 FILLCELL_X8 FILLER_62_467 ();
 FILLCELL_X4 FILLER_62_475 ();
 FILLCELL_X1 FILLER_62_479 ();
 FILLCELL_X8 FILLER_62_497 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X16 FILLER_63_33 ();
 FILLCELL_X1 FILLER_63_49 ();
 FILLCELL_X4 FILLER_63_53 ();
 FILLCELL_X16 FILLER_63_64 ();
 FILLCELL_X8 FILLER_63_80 ();
 FILLCELL_X2 FILLER_63_88 ();
 FILLCELL_X1 FILLER_63_90 ();
 FILLCELL_X2 FILLER_63_94 ();
 FILLCELL_X1 FILLER_63_103 ();
 FILLCELL_X32 FILLER_63_107 ();
 FILLCELL_X2 FILLER_63_139 ();
 FILLCELL_X1 FILLER_63_141 ();
 FILLCELL_X16 FILLER_63_159 ();
 FILLCELL_X4 FILLER_63_175 ();
 FILLCELL_X2 FILLER_63_179 ();
 FILLCELL_X4 FILLER_63_198 ();
 FILLCELL_X1 FILLER_63_205 ();
 FILLCELL_X4 FILLER_63_216 ();
 FILLCELL_X2 FILLER_63_220 ();
 FILLCELL_X8 FILLER_63_225 ();
 FILLCELL_X1 FILLER_63_233 ();
 FILLCELL_X2 FILLER_63_241 ();
 FILLCELL_X1 FILLER_63_243 ();
 FILLCELL_X1 FILLER_63_251 ();
 FILLCELL_X1 FILLER_63_289 ();
 FILLCELL_X2 FILLER_63_297 ();
 FILLCELL_X8 FILLER_63_306 ();
 FILLCELL_X2 FILLER_63_314 ();
 FILLCELL_X2 FILLER_63_350 ();
 FILLCELL_X4 FILLER_63_366 ();
 FILLCELL_X1 FILLER_63_370 ();
 FILLCELL_X4 FILLER_63_385 ();
 FILLCELL_X1 FILLER_63_389 ();
 FILLCELL_X4 FILLER_63_401 ();
 FILLCELL_X1 FILLER_63_405 ();
 FILLCELL_X4 FILLER_63_411 ();
 FILLCELL_X1 FILLER_63_454 ();
 FILLCELL_X2 FILLER_63_488 ();
 FILLCELL_X4 FILLER_63_499 ();
 FILLCELL_X2 FILLER_63_503 ();
 FILLCELL_X16 FILLER_64_1 ();
 FILLCELL_X4 FILLER_64_17 ();
 FILLCELL_X2 FILLER_64_45 ();
 FILLCELL_X1 FILLER_64_47 ();
 FILLCELL_X1 FILLER_64_55 ();
 FILLCELL_X1 FILLER_64_66 ();
 FILLCELL_X1 FILLER_64_72 ();
 FILLCELL_X4 FILLER_64_90 ();
 FILLCELL_X1 FILLER_64_94 ();
 FILLCELL_X4 FILLER_64_126 ();
 FILLCELL_X2 FILLER_64_130 ();
 FILLCELL_X2 FILLER_64_139 ();
 FILLCELL_X8 FILLER_64_148 ();
 FILLCELL_X2 FILLER_64_156 ();
 FILLCELL_X4 FILLER_64_161 ();
 FILLCELL_X2 FILLER_64_165 ();
 FILLCELL_X16 FILLER_64_170 ();
 FILLCELL_X8 FILLER_64_186 ();
 FILLCELL_X4 FILLER_64_194 ();
 FILLCELL_X2 FILLER_64_198 ();
 FILLCELL_X8 FILLER_64_222 ();
 FILLCELL_X4 FILLER_64_230 ();
 FILLCELL_X4 FILLER_64_251 ();
 FILLCELL_X1 FILLER_64_255 ();
 FILLCELL_X4 FILLER_64_269 ();
 FILLCELL_X2 FILLER_64_276 ();
 FILLCELL_X8 FILLER_64_317 ();
 FILLCELL_X2 FILLER_64_325 ();
 FILLCELL_X1 FILLER_64_327 ();
 FILLCELL_X1 FILLER_64_351 ();
 FILLCELL_X1 FILLER_64_376 ();
 FILLCELL_X1 FILLER_64_395 ();
 FILLCELL_X4 FILLER_64_409 ();
 FILLCELL_X2 FILLER_64_413 ();
 FILLCELL_X8 FILLER_64_420 ();
 FILLCELL_X4 FILLER_64_428 ();
 FILLCELL_X1 FILLER_64_432 ();
 FILLCELL_X2 FILLER_64_437 ();
 FILLCELL_X1 FILLER_64_439 ();
 FILLCELL_X1 FILLER_64_443 ();
 FILLCELL_X2 FILLER_64_452 ();
 FILLCELL_X32 FILLER_64_468 ();
 FILLCELL_X4 FILLER_64_500 ();
 FILLCELL_X1 FILLER_64_504 ();
 FILLCELL_X16 FILLER_65_1 ();
 FILLCELL_X4 FILLER_65_17 ();
 FILLCELL_X1 FILLER_65_21 ();
 FILLCELL_X4 FILLER_65_39 ();
 FILLCELL_X1 FILLER_65_43 ();
 FILLCELL_X8 FILLER_65_116 ();
 FILLCELL_X1 FILLER_65_124 ();
 FILLCELL_X4 FILLER_65_156 ();
 FILLCELL_X2 FILLER_65_160 ();
 FILLCELL_X8 FILLER_65_169 ();
 FILLCELL_X4 FILLER_65_177 ();
 FILLCELL_X4 FILLER_65_205 ();
 FILLCELL_X8 FILLER_65_223 ();
 FILLCELL_X2 FILLER_65_231 ();
 FILLCELL_X2 FILLER_65_257 ();
 FILLCELL_X4 FILLER_65_266 ();
 FILLCELL_X2 FILLER_65_270 ();
 FILLCELL_X1 FILLER_65_272 ();
 FILLCELL_X2 FILLER_65_280 ();
 FILLCELL_X1 FILLER_65_282 ();
 FILLCELL_X32 FILLER_65_290 ();
 FILLCELL_X16 FILLER_65_322 ();
 FILLCELL_X8 FILLER_65_341 ();
 FILLCELL_X2 FILLER_65_349 ();
 FILLCELL_X1 FILLER_65_351 ();
 FILLCELL_X4 FILLER_65_359 ();
 FILLCELL_X2 FILLER_65_386 ();
 FILLCELL_X8 FILLER_65_421 ();
 FILLCELL_X4 FILLER_65_429 ();
 FILLCELL_X2 FILLER_65_433 ();
 FILLCELL_X1 FILLER_65_435 ();
 FILLCELL_X1 FILLER_65_443 ();
 FILLCELL_X1 FILLER_65_463 ();
 FILLCELL_X16 FILLER_65_481 ();
 FILLCELL_X8 FILLER_65_497 ();
 FILLCELL_X16 FILLER_66_1 ();
 FILLCELL_X8 FILLER_66_17 ();
 FILLCELL_X2 FILLER_66_25 ();
 FILLCELL_X1 FILLER_66_27 ();
 FILLCELL_X2 FILLER_66_35 ();
 FILLCELL_X1 FILLER_66_37 ();
 FILLCELL_X4 FILLER_66_45 ();
 FILLCELL_X2 FILLER_66_49 ();
 FILLCELL_X1 FILLER_66_68 ();
 FILLCELL_X32 FILLER_66_86 ();
 FILLCELL_X8 FILLER_66_118 ();
 FILLCELL_X4 FILLER_66_143 ();
 FILLCELL_X1 FILLER_66_147 ();
 FILLCELL_X2 FILLER_66_165 ();
 FILLCELL_X4 FILLER_66_177 ();
 FILLCELL_X1 FILLER_66_181 ();
 FILLCELL_X2 FILLER_66_213 ();
 FILLCELL_X1 FILLER_66_215 ();
 FILLCELL_X16 FILLER_66_219 ();
 FILLCELL_X2 FILLER_66_235 ();
 FILLCELL_X16 FILLER_66_241 ();
 FILLCELL_X1 FILLER_66_257 ();
 FILLCELL_X4 FILLER_66_265 ();
 FILLCELL_X2 FILLER_66_269 ();
 FILLCELL_X1 FILLER_66_271 ();
 FILLCELL_X4 FILLER_66_296 ();
 FILLCELL_X1 FILLER_66_300 ();
 FILLCELL_X16 FILLER_66_308 ();
 FILLCELL_X8 FILLER_66_324 ();
 FILLCELL_X16 FILLER_66_343 ();
 FILLCELL_X2 FILLER_66_359 ();
 FILLCELL_X1 FILLER_66_361 ();
 FILLCELL_X4 FILLER_66_378 ();
 FILLCELL_X2 FILLER_66_403 ();
 FILLCELL_X2 FILLER_66_414 ();
 FILLCELL_X2 FILLER_66_433 ();
 FILLCELL_X2 FILLER_66_452 ();
 FILLCELL_X32 FILLER_66_471 ();
 FILLCELL_X2 FILLER_66_503 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X16 FILLER_67_33 ();
 FILLCELL_X8 FILLER_67_49 ();
 FILLCELL_X4 FILLER_67_57 ();
 FILLCELL_X2 FILLER_67_61 ();
 FILLCELL_X1 FILLER_67_63 ();
 FILLCELL_X4 FILLER_67_67 ();
 FILLCELL_X32 FILLER_67_74 ();
 FILLCELL_X32 FILLER_67_106 ();
 FILLCELL_X8 FILLER_67_138 ();
 FILLCELL_X4 FILLER_67_146 ();
 FILLCELL_X1 FILLER_67_167 ();
 FILLCELL_X2 FILLER_67_185 ();
 FILLCELL_X1 FILLER_67_187 ();
 FILLCELL_X2 FILLER_67_201 ();
 FILLCELL_X1 FILLER_67_203 ();
 FILLCELL_X16 FILLER_67_221 ();
 FILLCELL_X8 FILLER_67_237 ();
 FILLCELL_X4 FILLER_67_245 ();
 FILLCELL_X4 FILLER_67_269 ();
 FILLCELL_X2 FILLER_67_273 ();
 FILLCELL_X1 FILLER_67_275 ();
 FILLCELL_X4 FILLER_67_279 ();
 FILLCELL_X1 FILLER_67_283 ();
 FILLCELL_X4 FILLER_67_287 ();
 FILLCELL_X2 FILLER_67_291 ();
 FILLCELL_X1 FILLER_67_293 ();
 FILLCELL_X4 FILLER_67_297 ();
 FILLCELL_X2 FILLER_67_301 ();
 FILLCELL_X2 FILLER_67_306 ();
 FILLCELL_X1 FILLER_67_308 ();
 FILLCELL_X4 FILLER_67_326 ();
 FILLCELL_X2 FILLER_67_333 ();
 FILLCELL_X1 FILLER_67_335 ();
 FILLCELL_X2 FILLER_67_339 ();
 FILLCELL_X1 FILLER_67_341 ();
 FILLCELL_X4 FILLER_67_345 ();
 FILLCELL_X2 FILLER_67_349 ();
 FILLCELL_X16 FILLER_67_356 ();
 FILLCELL_X8 FILLER_67_372 ();
 FILLCELL_X4 FILLER_67_380 ();
 FILLCELL_X2 FILLER_67_384 ();
 FILLCELL_X1 FILLER_67_401 ();
 FILLCELL_X1 FILLER_67_411 ();
 FILLCELL_X1 FILLER_67_417 ();
 FILLCELL_X8 FILLER_67_421 ();
 FILLCELL_X2 FILLER_67_429 ();
 FILLCELL_X8 FILLER_67_443 ();
 FILLCELL_X4 FILLER_67_451 ();
 FILLCELL_X2 FILLER_67_455 ();
 FILLCELL_X8 FILLER_67_463 ();
 FILLCELL_X4 FILLER_67_471 ();
 FILLCELL_X16 FILLER_67_478 ();
 FILLCELL_X8 FILLER_67_494 ();
 FILLCELL_X2 FILLER_67_502 ();
 FILLCELL_X1 FILLER_67_504 ();
endmodule
